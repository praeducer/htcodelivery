14edfd8a3f876ab45ab7cd265ed015edc34cafd4|4|372|34.937113|-80.837892|6.978426046781553|82bdabfce564510321727cd9f4722b92937edf63|2015-01-26 12:18:00|0|149|34.977331|-81.027334|00041116005954|(FE)BABY BOTTLE POP|4111600595|REGISTER BARS|47|CANDY|7|G1 GROCERY|1|1.59|0.0|1
14edfd8a3f876ab45ab7cd265ed015edc34cafd4|4|372|34.937113|-80.837892|6.978426046781553|82bdabfce564510321727cd9f4722b92937edf63|2015-01-26 12:18:00|0|149|34.977331|-81.027334|00203184000006|PORK BOSTON BUTT|20318400000|PREMIUM PORK|641|PORK|137|MEAT|2|23.41|11.74|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|e6bc40257eebe28008628db0ec553ca85f0bfe3e|2014-11-25 21:40:00|0|412|35.195689|-80.826724|00075500200014|TEXAS PETE HOTTER SAUCE|7550020001|MEAT SAUCES|76|CONDIMENTS|11|G1 GROCERY|1|1.29|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|cd9d14ffce2b14a1ce3eaeab07c890dfdbc3c137|2015-01-20 21:26:00|0|208|35.17739|-80.80146|00071921008291|DIG FOR 1 TTRADITION CRUST PEP|7192100989|SUPER PREMIUM PIZZA|284|FROZEN PIZZA|892|FROZEN|5|3.89|0.39|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|54af6277b6e884516cac7dd136c4f79aee8fc1e1|2015-02-04 19:10:00|0|412|35.195689|-80.826724|00071921008291|DIG FOR 1 TTRADITION CRUST PEP|7192100989|SUPER PREMIUM PIZZA|284|FROZEN PIZZA|892|FROZEN|5|3.89|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|c4ff8d949fd316f5b0e5c91e000cd36f6a0c09bb|2015-03-09 20:53:00|0|208|35.17739|-80.80146|00071921008291|DIG FOR 1 TTRADITION CRUST PEP|7192100989|SUPER PREMIUM PIZZA|284|FROZEN PIZZA|892|FROZEN|5|3.89|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|8e4229c78ec829d8ec02149805b486210eae74e9|2014-10-24 22:04:00|0|412|35.195689|-80.826724|00839743001513|YELLOW TAIL PINK MOSCATO|83974300151|NFS POP OTHER RED|9944|POPULAR (4-$7.99)|885|WINE|13|6.99|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|e7f52abc948c3795b98e11781543ef2821f2ca6c|2014-12-09 07:38:00|0|412|35.195689|-80.826724|00012546006088|TRIDENT SPEARMINT BTL|1254631053|PEG GUM|45|CANDY|7|G1 GROCERY|1|3.79|0.79|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|d9efaacf811a649f3afbb5c811e895f2dea06c3c|2014-11-25 21:46:00|0|412|35.195689|-80.826724|00839743001513|YELLOW TAIL PINK MOSCATO|83974300151|NFS POP OTHER RED|9944|POPULAR (4-$7.99)|885|WINE|13|5.99|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|382a61ff099be65a68fc88387f6ad7dc3999d011|2014-12-31 20:17:00|0|208|35.17739|-80.80146|00010900000215|REYNOLDS FOIL HEAVY DUTY 50 FT|1090000015|NFS-ALUMINUM FOIL|440|WRAPPING MATERIALS & BAGS|76|G1 GROCERY|1|3.99|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|e7f52abc948c3795b98e11781543ef2821f2ca6c|2014-12-09 07:38:00|0|412|35.195689|-80.826724|00024000507918|FRUIT NAT. MANDARIN ORANG 7 OZ|2400050785|FRESH JARRED FRUIT|578|OTHER MERCHANDISE|136|PRODUCE|4|1.5|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|c4ff8d949fd316f5b0e5c91e000cd36f6a0c09bb|2015-03-09 20:53:00|0|208|35.17739|-80.80146|00884395063013|LUCKS BEAN PINTO 29|88439506301|CANNED BEANS|242|VEGETABLES-CAN/JAR|39|G1 GROCERY|1|1.89|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|2f48e4568445fe930d4e39e44fffed5b818bf165|2014-10-13 14:36:00|0|208|35.17739|-80.80146|00754441777716|GREAT FISH WHITING FILLETS|75444177771|FISH FILLETS/STEAKS PKGD|663|FISH FILLETS/STEAKS|154|SEAFOOD|12|7.99|3.02|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|7260067d4b9244a0976dcda47e5c5862f8a4fe8a|2014-12-16 19:31:00|0|208|35.17739|-80.80146|00202518000002|HT NAT 90% LEAN GROUND BEEF|20251800000|NATURAL/ORGANIC BEEF|642|BEEF|49|MEAT|2|15.26|1.91|2
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|b0ab7811d88bdb3a5b32e6e02aa548cd45a8b834|2015-02-15 19:59:00|0|208|35.17739|-80.80146|00202518000002|HT NAT 90% LEAN GROUND BEEF|20251800000|NATURAL/ORGANIC BEEF|642|BEEF|49|MEAT|2|15.42|1.93|2
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|b0ab7811d88bdb3a5b32e6e02aa548cd45a8b834|2015-02-15 19:59:00|0|208|35.17739|-80.80146|00204069000005|COO GREEN CABBAGE||FRESH CABBAGE|530|FRESH PRODUCE|64|PRODUCE|4|3.38|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|e7f52abc948c3795b98e11781543ef2821f2ca6c|2014-12-09 07:38:00|0|412|35.195689|-80.826724|00305730196208|ADVIL ALLERGY&CONGESTION|30573019620|DEX ADULT/CHILDREN|4236|COUGH/COLD/SINUS|1200|HBC|17|10.59|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|f3f4487d7a42fa7916ed1850fb488b8039e58000|2015-02-17 19:15:00|0|412|35.195689|-80.826724|00300410606862|ORAL B INDICATOR TWIN SOFT #17|30041060686|TOOTH BRUSH-PREMIUM|4056|ORAL HYGIENE|1080|HBC|17|3.99|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|22d82c6e6c3b9854c18b00be9494843075d4e732|2014-10-13 13:36:00|0|412|35.195689|-80.826724|00208222000000|WC FRESH FLOUNDER FILLET (US)|20822200000|FISH FILLETS WILD CGHT|660|FISH FILLETS/STEAKS|154|SEAFOOD|12|3.95|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|90ac52504f452962f05c883f38af11521164ac09|2014-10-12 20:35:00|0|208|35.17739|-80.80146|00208222000000|WC FRESH FLOUNDER FILLET (US)|20822200000|FISH FILLETS WILD CGHT|660|FISH FILLETS/STEAKS|154|SEAFOOD|12|8.36|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|5bf0726886e91d2b41dead6e8d3f8b0fb5193fb9|2014-11-13 20:37:00|0|412|35.195689|-80.826724|00611443340266|KITCHEN BASICS STOCK TURKEY|61144334026|BROTH|214|SOUP|33|G1 GROCERY|1|7.38|0.9|2
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|635e647747bf5a3bd9ccc6e7789808bc890e9b06|2015-03-05 18:06:00|0|171|35.141204|-80.739|00201657000003|HT GROUND BEEF CHUCK 80% LEAN|20165700000|GROUND BEEF|297|BEEF|49|MEAT|2|5.25|1.17|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|635e647747bf5a3bd9ccc6e7789808bc890e9b06|2015-03-05 18:06:00|0|171|35.141204|-80.739|00041570056219|ALMOND BREEZE VANILLA|4157005617|ALMOND MILK|1265|MILK|57|DAIRY|3|3.25|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|635e647747bf5a3bd9ccc6e7789808bc890e9b06|2015-03-05 18:06:00|0|171|35.141204|-80.739|00042456005055|PIROULINE TIN CHOC HAZELNUT|4245600505|SPECIALTY COOKIES|1250|COOKIES|12|G1 GROCERY|1|5.99|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|54af6277b6e884516cac7dd136c4f79aee8fc1e1|2015-02-04 19:10:00|0|412|35.195689|-80.826724|00046704033203|TGIF LOADED FRIES CHEESE&BACON|4670406840|FROZEN SNACKS|1277|FROZEN SANDWICH AND SNACKS|279|FROZEN|5|3.99|0.65|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|da05fbbbb8102dea9bf6df2357b1d429d528cdd0|2014-12-17 19:31:00|0|208|35.17739|-80.80146|00046704033203|TGIF LOADED FRIES CHEESE&BACON|4670406840|FROZEN SNACKS|1277|FROZEN SANDWICH AND SNACKS|279|FROZEN|5|3.99|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|cd9d14ffce2b14a1ce3eaeab07c890dfdbc3c137|2015-01-20 21:26:00|0|208|35.17739|-80.80146|00046704068403|TGIF CHEDDAR & BACON POT SKINS|4670406840|FROZEN SNACKS|1277|FROZEN SANDWICH AND SNACKS|279|FROZEN|5|3.99|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|22fc4c32545e2649ac02785990f483449c244a64|2015-01-26 15:17:00|0|412|35.195689|-80.826724|00046704033203|TGIF LOADED FRIES CHEESE&BACON|4670406840|FROZEN SNACKS|1277|FROZEN SANDWICH AND SNACKS|279|FROZEN|5|3.99|0.65|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|5ba4a64f78c48e35ccb7245774882f7f4fec5684|2015-02-03 21:31:00|0|208|35.17739|-80.80146|00048500021828|PP TROP RASPBRY LEMONADE 59 OZ|4850002180|OTHER FRUIT JUICES|338|JUICES & DRINKS-REFRIGERATED|56|DAIRY|3|3.29|1.65|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|efd67486fa9be6e654d850ed2616429a5920f071|2014-11-27 13:43:00|0|412|35.195689|-80.826724|00043000009536|COOL WHIP WHIPPED TOPPING|4300000953|TOPPINGS FROZEN|272|DESSERTS FROZEN|307|FROZEN|5|2.0|1.01|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|20d577dc350ad05ec1b9e414df7146444a49d550|2014-12-28 13:34:00|0|412|35.195689|-80.826724|00018200149917|BUD LIGHT LIME 6PK LNNR|1820014991|DOMESTIC SINGLES/SIX PACKS|457|DOMESTIC BEER|82|BEER|16|7.99|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|f2a60a1a5fa2c037ce76fd2b6b7ad942a65b19f7|2014-10-03 18:26:00|0|208|35.17739|-80.80146|00009800123018|ROCHER|980012301|REGISTER BARS|47|CANDY|7|G1 GROCERY|1|1.5|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|382a61ff099be65a68fc88387f6ad7dc3999d011|2014-12-31 20:17:00|0|208|35.17739|-80.80146|00030400771712|ANGEL SOFT SOFT/STRONG 9DR|3040077171|NFS-TOILET TISSUE|427|PAPER/PLASTIC PRODUCTS|72|G1 GROCERY|1|6.99|1.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|657db625e28d2eaa29f8d42ccc3e96930dc4060e|2015-01-28 18:58:00|0|412|35.195689|-80.826724|00020000001104|GG NIBLET CORN BUTTER SAUCE|2000000065|BOX VEG|1275|VEGETABLES-FROZEN|50|FROZEN|5|1.89|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|9f32c3bb2632bee6cadb7eec615a7e8fedd3824c|2014-09-12 23:36:00|0|208|35.17739|-80.80146|00054400002669|A1 MARINADE MIX - ORIGINAL|5440000266|SEASONING PACKETS|80|SPICES/SEASONINGS/EXTRACTS|34|G1 GROCERY|1|1.49|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|d612f02b2556769e3971cbc629697502db30356e|2014-11-11 23:00:00|0|412|35.195689|-80.826724|00072036955500|BULK  BAGELS||BULK (BAGELS)|1635|BAGELS|375|BAKERY|14|0.75|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|d5940d560163c31c68191569828de9c800623160|2015-01-15 19:32:00|0|412|35.195689|-80.826724|00072036952981|OLD FASHION FUDGE CAKE SLICE|7203695298|DESSERT CAKES|1654|CAKES|381|BAKERY|14|2.59|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|54af6277b6e884516cac7dd136c4f79aee8fc1e1|2015-02-04 19:10:00|0|412|35.195689|-80.826724|00072036952981|OLD FASHION FUDGE CAKE SLICE|7203695298|DESSERT CAKES|1654|CAKES|381|BAKERY|14|2.59|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|cd9d14ffce2b14a1ce3eaeab07c890dfdbc3c137|2015-01-20 21:26:00|0|208|35.17739|-80.80146|00072036952981|OLD FASHION FUDGE CAKE SLICE|7203695298|DESSERT CAKES|1654|CAKES|381|BAKERY|14|2.59|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|c4ba739daf7aa5a685bf65adc8ed4c946af70f28|2014-12-15 15:49:00|0|208|35.17739|-80.80146|00072036880734|HT BAKER POTATO 4 CT PKG|7203688073|FRESH POTATOES|523|FRESH PRODUCE|64|PRODUCE|4|3.69|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|635e647747bf5a3bd9ccc6e7789808bc890e9b06|2015-03-05 18:06:00|0|171|35.141204|-80.739|00041780001887|UTZ RED HOT CHIP|4178000011|POTATO CHIPS|201|SNACKS|31|G1 GROCERY|1|4.29|1.3|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|8e1c58c48a31042e63c5374ab2eb19612a5d163e|2014-09-19 18:19:00|0|160|35.152722|-80.825175|00041780001887|UTZ RED HOT CHIP|4178000011|POTATO CHIPS|201|SNACKS|31|G1 GROCERY|1|8.58|2.14|2
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|20d577dc350ad05ec1b9e414df7146444a49d550|2014-12-28 13:34:00|0|412|35.195689|-80.826724|00051000159045|CHUNKY MW CHILI ROADHOUSE|5100014880|RTS MICROWAVE|1499|SOUP|33|G1 GROCERY|1|2.79|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|5ba4a64f78c48e35ccb7245774882f7f4fec5684|2015-02-03 21:31:00|0|208|35.17739|-80.80146|00051500222416|PILLSBURY BEST FLOUR-UNBLEACHD|5150020441|REMAINING FLOUR|103|FLOUR|15|G1 GROCERY|1|2.69|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|d5940d560163c31c68191569828de9c800623160|2015-01-15 19:32:00|0|412|35.195689|-80.826724|00071279231006|F.E. BABY SPRING SALAD MIX|7127923100|PACKAGED SALADS|555|FRESH PRODUCE|64|PRODUCE|4|1.99|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|9fa9bf07f2e593bc3f6439d4e0d6a0e7f72e9f8b|2014-12-26 19:10:00|0|412|35.195689|-80.826724|00071279231006|F.E. BABY SPRING SALAD MIX|7127923100|PACKAGED SALADS|555|FRESH PRODUCE|64|PRODUCE|4|1.99|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|a44a58f116c753073356093820799cd37b1f1971|2014-10-04 21:34:00|0|412|35.195689|-80.826724|00204879000004|HT TEXAS CAVIAR||SERVICE BAR|566|FRESH PRODUCE|64|PRODUCE|4|1.22|0.07|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|e7f52abc948c3795b98e11781543ef2821f2ca6c|2014-12-09 07:38:00|0|412|35.195689|-80.826724|00204826000002|KIWI EXPLOSION||FRESH CUT FRUIT|562|FRESH PRODUCE|64|PRODUCE|4|7.44|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|7260067d4b9244a0976dcda47e5c5862f8a4fe8a|2014-12-16 19:31:00|0|208|35.17739|-80.80146|00208895000000|FR TILAPIA FILLET|20889500000|FISH FLTS/STK FARM RAISD|648|FISH FILLETS/STEAKS|154|SEAFOOD|12|10.58|2.45|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|d9efaacf811a649f3afbb5c811e895f2dea06c3c|2014-11-25 21:46:00|0|412|35.195689|-80.826724|00051000138095|CHUNKY GRILLED SIRLOIN|5100000524|RTS CANNED|1201|SOUP|33|G1 GROCERY|1|1.99|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|5ba4a64f78c48e35ccb7245774882f7f4fec5684|2015-02-03 21:31:00|0|208|35.17739|-80.80146|00071025015621|BUNNY B&S ROLL|7102501562|DINNER ROLLS|1039|MEAL ACCOMPANIMENT|166|COMMERCIAL BAKERY|7|2.59|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|e6bc40257eebe28008628db0ec553ca85f0bfe3e|2014-11-25 21:40:00|0|412|35.195689|-80.826724|00071025015621|BUNNY B&S ROLL|7102501562|DINNER ROLLS|1039|MEAL ACCOMPANIMENT|166|COMMERCIAL BAKERY|7|2.59|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|7260067d4b9244a0976dcda47e5c5862f8a4fe8a|2014-12-16 19:31:00|0|208|35.17739|-80.80146|00072036320223|HT VEGETABLE OIL|7203632016|SALAD & COOKING OIL|195|SHORTENING/OIL|30|G1 GROCERY|1|3.0|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|a44a58f116c753073356093820799cd37b1f1971|2014-10-04 21:34:00|0|412|35.195689|-80.826724|00072940100430|VINE RIPE PASTA SC MUSHROOM|7294010041|PASTA SC VALUE|1221|PASTA SAUCES|275|G1 GROCERY|1|0.97|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|a7eb3d5a4877b1d4e554118fa8c81927a9c71126|2015-01-12 17:35:00|0|208|35.17739|-80.80146|00077782029833|JOHNSONVILLE BEEF BRATWURST|7778202983|SMOKED SAUSAGE LINKS|488|DINNER SAUSAGE|104|CASE READY MEATS|19|3.99|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|635e647747bf5a3bd9ccc6e7789808bc890e9b06|2015-03-05 18:06:00|0|171|35.141204|-80.739|00208965000008|HT FRESH CHICKEN DRUMMETTES|20896500000|FRESH HT CHICKEN|977|POULTRY|201|MEAT|2|7.359999999999999|0.0|2
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|54af6277b6e884516cac7dd136c4f79aee8fc1e1|2015-02-04 19:10:00|0|412|35.195689|-80.826724|00204011000008|BANANAS, YELLOW||FRESH BANANAS|502|FRESH PRODUCE|64|PRODUCE|4|0.67|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|ae9ead32ee800b4131d4db3a4d9ab8e8ab8d5b8f|2015-01-20 20:25:00|0|208|35.17739|-80.80146|00078000152166|CD GINGER ALE 12 PACK|7800001180|REGULAR|55|CARBONATED BEVERAGES|8|BEVERAGE|23|6.79|1.79|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|d4f584e05ff3f88e10db1fb946f0a77d9a1efac1|2014-10-20 15:56:00|0|412|35.195689|-80.826724|00039400015901|BUSH BKD BEAN EZO HMSTY|3940001606|BAKED BEANS|243|VEGETABLES-CAN/JAR|39|G1 GROCERY|1|1.39|0.39|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|b0ab7811d88bdb3a5b32e6e02aa548cd45a8b834|2015-02-15 19:59:00|0|208|35.17739|-80.80146|00074336100055|HUNTER  WHOLE MILK|7433610005|FRESH MILK|342|MILK|57|DAIRY|3|2.59|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|a44a58f116c753073356093820799cd37b1f1971|2014-10-04 21:34:00|0|412|35.195689|-80.826724|00070897013315|FOSTERS LAGER 25.4OZ CAN|7089701331|IMPORT BEER|459|IMPORT BEER|83|BEER|16|1.99|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|a44a58f116c753073356093820799cd37b1f1971|2014-10-04 21:34:00|0|412|35.195689|-80.826724|00076808280098|BARILLA PASTA THIN SPAG|7680828008|WHSE PASTA CORE|149|PASTA|23|G1 GROCERY|1|1.69|0.69|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|748a867f4d79bc8f0e0118f4f21bd668469edec1|2015-02-19 23:13:00|0|208|35.17739|-80.80146|00041260331091|OW GOLD THUMB TACKS|4126033109|TACKS & PAPER CLIPS|6764|SCHOOL & OFFICE SUPPLY|1564|GM|18|1.99|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|9d93788654c8fe94e01a11696dd195b6bb599e59|2014-10-01 23:51:00|0|208|35.17739|-80.80146|00044700000953|OSCAR MAYER BEEF FRANKS|4470007502|BEEF WIENERS|484|WIENERS|101|CASE READY MEATS|19|4.99|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|d5940d560163c31c68191569828de9c800623160|2015-01-15 19:32:00|0|412|35.195689|-80.826724|00041335332176|KENS DRS RANCH|4133533217|SALAD DRESSINGS-LIQUID|184|SALAD DRESSING/MAYONNAISE|28|G1 GROCERY|1|2.29|1.29|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|9f32c3bb2632bee6cadb7eec615a7e8fedd3824c|2014-09-12 23:36:00|0|208|35.17739|-80.80146|00041196406979|PROG ARTISAN SM WH BEAN WT VEG|4119640699|RTS ASEPTIC|1437|SOUP|33|G1 GROCERY|1|3.49|0.99|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|5ba4a64f78c48e35ccb7245774882f7f4fec5684|2015-02-03 21:31:00|0|208|35.17739|-80.80146|00030000315514|QKR MEDLEY PEACH ALMOND|3000031551|HOT CEREAL|60|CEREAL|9|G1 GROCERY|1|1.99|0.49|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|d612f02b2556769e3971cbc629697502db30356e|2014-11-11 23:00:00|0|412|35.195689|-80.826724|00024000507932|FRUIT NAT. NSA GRAPEFRT 6.5 OZ|2400050785|FRESH JARRED FRUIT|578|OTHER MERCHANDISE|136|PRODUCE|4|1.5|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|1f085a1fa268e94c8b9feb336ecfe54908818d1b|2014-11-12 19:58:00|0|412|35.195689|-80.826724|00068274934711|NESTLE PURE LIFE .5L 24PK|6827493471|NON CARBONATED WATER|31|BOTTLED WATER|4|G1 GROCERY|1|4.99|1.2|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|f9dc859b6851ef458ace7508afbf4db14f0cbaea|2014-12-05 19:43:00|0|412|35.195689|-80.826724|00068274934711|NESTLE PURE LIFE .5L 24PK|6827493471|NON CARBONATED WATER|31|BOTTLED WATER|4|G1 GROCERY|1|4.99|2.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|a44a58f116c753073356093820799cd37b1f1971|2014-10-04 21:34:00|0|412|35.195689|-80.826724|00068274934711|NESTLE PURE LIFE .5L 24PK|6827493471|NON CARBONATED WATER|31|BOTTLED WATER|4|G1 GROCERY|1|4.99|1.2|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|22d82c6e6c3b9854c18b00be9494843075d4e732|2014-10-13 13:36:00|0|412|35.195689|-80.826724|00025000047664|MINUTE MAID BERRY PUNCH|2500004748|OTHER FRUIT JUICES|338|JUICES & DRINKS-REFRIGERATED|56|DAIRY|3|2.0|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|d4f584e05ff3f88e10db1fb946f0a77d9a1efac1|2014-10-20 15:56:00|0|412|35.195689|-80.826724|00025000047664|MINUTE MAID BERRY PUNCH|2500004748|OTHER FRUIT JUICES|338|JUICES & DRINKS-REFRIGERATED|56|DAIRY|3|2.0|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|e7f52abc948c3795b98e11781543ef2821f2ca6c|2014-12-09 07:38:00|0|412|35.195689|-80.826724|00312546627543|(JHK) HALLS DEF VIT C CITRUS|31254662920|COUGH DROP-ADULT|4207|COUGH/COLD/SINUS|1200|HBC|17|2.29|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|b0ab7811d88bdb3a5b32e6e02aa548cd45a8b834|2015-02-15 19:59:00|0|208|35.17739|-80.80146|00033383490335|GREEN BELL PEPPER 2CT PK|3338349033|FRESH PEPPERS|533|FRESH PRODUCE|64|PRODUCE|4|1.27|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|ae9ead32ee800b4131d4db3a4d9ab8e8ab8d5b8f|2015-01-20 20:25:00|0|208|35.17739|-80.80146|00031200330147|OS 100% CRANBERRY JUICE|3120033014|CRANBERRY JUICE/DRINKS-SHELF|130|JUICES/DRINKS-SHELF STABLE|20|G1 GROCERY|1|7.98|1.99|2
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|9fa9bf07f2e593bc3f6439d4e0d6a0e7f72e9f8b|2014-12-26 19:10:00|0|412|35.195689|-80.826724|00051000167767|CHUNKY HR OLD FASH VEG BEEF|5100000524|RTS CANNED|1201|SOUP|33|G1 GROCERY|1|1.99|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|efd67486fa9be6e654d850ed2616429a5920f071|2014-11-27 13:43:00|0|412|35.195689|-80.826724|00070640034024|B BUNNY PREM HOMEMADE VANILLA|7064003404|PREMIUM ICE CREAM|252|ICE CREAM|45|FROZEN|5|6.79|2.81|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|e7f52abc948c3795b98e11781543ef2821f2ca6c|2014-12-09 07:38:00|0|412|35.195689|-80.826724|00013100501346|I/OHT HDAY FACIAL TISSUE SHPR|1310050134|NFS-FACIAL TISSUE|424|PAPER/PLASTIC PRODUCTS|72|G1 GROCERY|1|1.79|0.29|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|382a61ff099be65a68fc88387f6ad7dc3999d011|2014-12-31 20:17:00|0|208|35.17739|-80.80146|00204619000004|COO TURNIP GREENS, BULK||FRESH GREENS|535|FRESH PRODUCE|64|PRODUCE|4|1.67|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|f9dc859b6851ef458ace7508afbf4db14f0cbaea|2014-12-05 19:43:00|0|412|35.195689|-80.826724|00017400100773|SUCCESS RICE 4 BIB WHITE|1740010077|RICE-PACKAGED & BULK|239|RICE GRAINS AND BEANS|38|G1 GROCERY|1|2.79|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|e7f52abc948c3795b98e11781543ef2821f2ca6c|2014-12-09 07:38:00|0|412|35.195689|-80.826724|00312546631540|HALLS TROP FRUIT-63154|31254662380|COUGH DROP-ADULT|4207|COUGH/COLD/SINUS|1200|HBC|17|1.89|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|0fba0254bbb79fea55fa049358a36c9f3a9b4b61|2015-03-08 10:31:00|0|412|35.195689|-80.826724|00022000008992|EXTRA SPEARMINT|2200000899|REGISTER GUM|48|CANDY|7|G1 GROCERY|1|1.19|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|635e647747bf5a3bd9ccc6e7789808bc890e9b06|2015-03-05 18:06:00|0|171|35.141204|-80.739|00203316000003|PORK LOIN CHOPS BONE-IN THIN|20331600000|PREMIUM PORK|641|PORK|137|MEAT|2|10.21|0.0|2
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|9d93788654c8fe94e01a11696dd195b6bb599e59|2014-10-01 23:51:00|0|208|35.17739|-80.80146|00204011000008|BANANAS, YELLOW||FRESH BANANAS|502|FRESH PRODUCE|64|PRODUCE|4|0.53|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|c4ff8d949fd316f5b0e5c91e000cd36f6a0c09bb|2015-03-09 20:53:00|0|208|35.17739|-80.80146|00204011000008|BANANAS, YELLOW||FRESH BANANAS|502|FRESH PRODUCE|64|PRODUCE|4|0.4|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|9f32c3bb2632bee6cadb7eec615a7e8fedd3824c|2014-09-12 23:36:00|0|208|35.17739|-80.80146|00204011000008|BANANAS, YELLOW||FRESH BANANAS|502|FRESH PRODUCE|64|PRODUCE|4|0.31|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|e6bc40257eebe28008628db0ec553ca85f0bfe3e|2014-11-25 21:40:00|0|412|35.195689|-80.826724|00072036632203|HT GRADE A    LARGE EGGS|7203663220|EGGS|330|EGGS FRESH|55|DAIRY|3|1.45|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|9d93788654c8fe94e01a11696dd195b6bb599e59|2014-10-01 23:51:00|0|208|35.17739|-80.80146|00072036632203|HT GRADE A    LARGE EGGS|7203663220|EGGS|330|EGGS FRESH|55|DAIRY|3|1.45|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|7260067d4b9244a0976dcda47e5c5862f8a4fe8a|2014-12-16 19:31:00|0|208|35.17739|-80.80146|00070459005277|NY SOFT GARLIC PULL APARTS|7045900555|FROZEN GARLIC TOAST AND BRD|1461|FROZEN DOUGH|40|FROZEN|5|3.89|1.39|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|635e647747bf5a3bd9ccc6e7789808bc890e9b06|2015-03-05 18:06:00|0|171|35.141204|-80.739|00021788916291|BISCOFF COOKIES CRISP EURO|2178891629|SPECIALTY COOKIES|1250|COOKIES|12|G1 GROCERY|1|4.59|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|e7f52abc948c3795b98e11781543ef2821f2ca6c|2014-12-09 07:38:00|0|412|35.195689|-80.826724|00073852029437|PURELL OCEAN KISS PUMP BOTTLE|7385202390|ANTISEPTIC/DISINFECTANT|4828|FIRST AID|1235|HBC|17|1.79|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|635e647747bf5a3bd9ccc6e7789808bc890e9b06|2015-03-05 18:06:00|0|171|35.141204|-80.739|00201655000005|HT PREMIUM GRND BEEF 80% LEAN|20165500000|GROUND BEEF|297|BEEF|49|MEAT|2|5.79|0.73|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|d0411e9005a60617680e7bb993c072192d3176a1|2015-03-05 18:09:00|0|171|35.141204|-80.739|00201939000004|ANGUS BEEF SHORT RIBS|20193900000|ANGUS BEEF|299|BEEF|49|MEAT|2|11.02|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|635e647747bf5a3bd9ccc6e7789808bc890e9b06|2015-03-05 18:06:00|0|171|35.141204|-80.739|00201939000004|ANGUS BEEF SHORT RIBS|20193900000|ANGUS BEEF|299|BEEF|49|MEAT|2|19.71|0.0|2
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|7260067d4b9244a0976dcda47e5c5862f8a4fe8a|2014-12-16 19:31:00|0|208|35.17739|-80.80146|00070640004591|BB PERSONALS NSA DBL STRWBERRY|7064000461|SUPER PREMIUM ICE CREAM|275|ICE CREAM|45|FROZEN|5|1.34|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|22d82c6e6c3b9854c18b00be9494843075d4e732|2014-10-13 13:36:00|0|412|35.195689|-80.826724|00073420000066|DAISY SOUR CREAM|7342000006|SOUR CREAM|322|CULTURES|53|DAIRY|3|1.79|0.59|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|c4ba739daf7aa5a685bf65adc8ed4c946af70f28|2014-12-15 15:49:00|0|208|35.17739|-80.80146|00073420000110|DAISY SOUR CREAM|7342000011|SOUR CREAM|322|CULTURES|53|DAIRY|3|2.39|0.0|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|90ac52504f452962f05c883f38af11521164ac09|2014-10-12 20:35:00|0|208|35.17739|-80.80146|00027000612866|WESSON VEGETABLE OIL|2700061286|SALAD & COOKING OIL|195|SHORTENING/OIL|30|G1 GROCERY|1|4.59|1.09|1
14f71b19b67ee23ca147d8c4eda0ddb6204896e1|4|166|35.323246|-80.945176|1.8545010906496384|635e647747bf5a3bd9ccc6e7789808bc890e9b06|2015-03-05 18:06:00|0|171|35.141204|-80.739|00077975080047|SOH SOURDOUGH NIBBLERS|7797508005|PRETZELS|202|SNACKS|31|G1 GROCERY|1|3.49|0.99|1
