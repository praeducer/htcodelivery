customer|tier|homeStore|homeStoreLat|homeStoreLon|distance|receipt|datetime|onlineFlag|store|storeLat|storeLon|upc|desc|mupc|subcat|subcat_num|cat|cat_num|dept|dept_num|sales|discount|quantity
bdddad32053f7f53031d5dbfdc0692a01837373f|3|66|35.059823|-80.816172|0.8398516561798964|dd4b97177ebb1ea7b6732cc585ac8d0992ae1f87|2014-09-11 21:04:00|0|11|35.053394|-80.848528|00000000008070|24PK RECYCLING FEE|807|REGULAR|55|CARBONATED BEVERAGES|8|BEVERAGE|23|2.0|0.0|1
388acdabfcf14371f3e3715b783d2dd86eaef343|2|11|35.053394|-80.848528|1.4875527788777978|3f4560138de0fe76ca4e4cfa53eaf893a8fee8b1|2014-11-18 20:07:00|0|11|35.053394|-80.848528|00000000008070|24PK RECYCLING FEE|807|REGULAR|55|CARBONATED BEVERAGES|8|BEVERAGE|23|2.0|0.0|1
244a61514bf4e7cc8b53b1e86f1386b15e63fd2a|3|182|34.95459|-80.758228|19.173942376492086|7b656442ba85ad1e5a63d921cef06c69e622d780|2015-03-02 15:24:00|0|372|34.937113|-80.837892|00000000958940|CHEESE DANISH|95894|PASTRY|1599|STARBUCKS|370|COFFEE SHOP|22|2.45|0.0|1
fdc67de3d4ee9077be1fee92c19423b221c1e46a|2|317|35.024464|-80.847383|2.4816496149061793|cfc050d7c08982c1a2093e103493ab7cfd7dfac6|2014-12-16 10:12:00|0|372|34.937113|-80.837892|00000000958940|CHEESE DANISH|95894|PASTRY|1599|STARBUCKS|370|COFFEE SHOP|22|2.45|0.0|1
7abefb9b3f88d0fec923b34aba3fd231d95ee115|1|30|35.096737|-80.78468|0.8942038473266252|cfd7fe8b6ca0bd4438f6c4e3e7bbfeaccc574ee3|2014-10-02 16:08:00|0|372|34.937113|-80.837892|00000000958940|CHEESE DANISH|95894|PASTRY|1599|STARBUCKS|370|COFFEE SHOP|22|2.45|0.0|1
84d2310ad7d1c591f226386bb55e02cd1ed1bc6e|1|82|35.03469|-80.97058|2.4880644398940994|e9ef23c87e7a69578bfbfea87fd164b004087c61|2015-01-30 08:12:00|0|82|35.03469|-80.97058|00000000958940|CHEESE DANISH|95894|PASTRY|1599|STARBUCKS|370|COFFEE SHOP|22|2.45|1.23|1
341201b209fb1701d238bbc58a68d05037ded471|1|471|35.442529|-80.762919|3.1871599718814276|2c023c9a1c3071dcbdded317a178bd4b0d8d4fe2|2014-09-18 16:43:00|0|268|35.500972|-80.860108|00000000959570|SLTD CRML MOCHA FRAP GRAN|95957|NFS BEVERAGE BLEND|1597|NFS STARBUCKS|369|COFFEE SHOP|22|4.75|0.0|1
defa10073f7ec3e18521dda2ebfe5d7ba677b849|2|99|35.585842|-80.875654|1.7507069169423124|d9ca616accc6c4a5df79e67e049fa359e435faa0|2014-09-21 16:39:00|0|274|35.603432|-80.895009|00000000959570|SLTD CRML MOCHA FRAP GRAN|95957|NFS BEVERAGE BLEND|1597|NFS STARBUCKS|369|COFFEE SHOP|22|4.75|0.0|1
d7984a943579faa1f7871ed6e99575bcf1ac4ea2|2|157|35.124987|-80.709466|1.7907478604233464|56b5b36a538aa407a0dc757bc1779b5b33e163d8|2014-12-05 16:52:00|0|157|35.124987|-80.709466|00000000959570|SLTD CRML MOCHA FRAP GRAN|95957|NFS BEVERAGE BLEND|1597|NFS STARBUCKS|369|COFFEE SHOP|22|4.75|1.75|1
8d7d623dbf256d6792b6c34cd3c6df26c5fe2cec|2|157|35.124987|-80.709466|0.8515396021260951|78c97285ff7c1487b961147f9ba2a74c84a73870|2014-09-20 15:21:00|0|157|35.124987|-80.709466|00000000959570|SLTD CRML MOCHA FRAP GRAN|95957|NFS BEVERAGE BLEND|1597|NFS STARBUCKS|369|COFFEE SHOP|22|9.5|4.75|2
2fc86b6946aebfcd4ac59eec0e3921028e312a66|4|372|34.937113|-80.837892|20.379030753940455|9e967287f86e46ca8ead44b90865c31f0bdf4439|2014-10-19 15:09:00|0|372|34.937113|-80.837892|00000000959570|SLTD CRML MOCHA FRAP GRAN|95957|NFS BEVERAGE BLEND|1597|NFS STARBUCKS|369|COFFEE SHOP|22|4.75|0.0|1
559affaa6d1aefcb82c87f1256a975c09ec225cd|1|208|35.17739|-80.80146|2.335460904688238|a3ef61c4d6f2a72b58d5995b048a3f4058e2686e|2014-09-27 11:44:00|0|157|35.124987|-80.709466|00000000968840|CAFFE MOCHA GRANDE|96884|NFS BEVERAGE ESPRESSO|1589|NFS STARBUCKS|369|COFFEE SHOP|22|4.15|0.0|1
43c4e7d038650842db46e8c165e398a00e69f705|1|268|35.500972|-80.860108|4.368003822551078|75112a56364d4992d08569330d122d996c38c2f5|2014-11-17 06:51:00|0|268|35.500972|-80.860108|00000000968840|CAFFE MOCHA GRANDE|96884|NFS BEVERAGE ESPRESSO|1589|NFS STARBUCKS|369|COFFEE SHOP|22|4.15|0.0|1
b73a7f4e37273d5f5263cf9b421b37176e06b2a3|4|372|34.937113|-80.837892|21.404787733890718|1f9efcb09be135369a3c47daeaa9f9e04ce229a4|2014-11-22 10:40:00|0|475|35.061685|-80.994596|00000000968840|CAFFE MOCHA GRANDE|96884|NFS BEVERAGE ESPRESSO|1589|NFS STARBUCKS|369|COFFEE SHOP|22|4.15|0.0|1
43c4e7d038650842db46e8c165e398a00e69f705|1|268|35.500972|-80.860108|4.368003822551078|f0f072e82e91273e33b7604c551d962eac1d9679|2015-03-03 07:46:00|0|268|35.500972|-80.860108|00000000968840|CAFFE MOCHA GRANDE|96884|NFS BEVERAGE ESPRESSO|1589|NFS STARBUCKS|369|COFFEE SHOP|22|4.15|0.0|1
acd4bb36b708150dc2ab5cf1a58c677c762493ac|2|372|34.937113|-80.837892|1.2604840754487858|ffbaad30a17ec3e628c98f5fa6e8e05bf03f84d9|2014-12-14 11:32:00|0|372|34.937113|-80.837892|00000000968840|CAFFE MOCHA GRANDE|96884|NFS BEVERAGE ESPRESSO|1589|NFS STARBUCKS|369|COFFEE SHOP|22|4.15|0.0|1
ff1fb0d7a37f0afa26313d15a969442febb8196e|3|209|35.40953|-80.86175|1.206911972128497|eda8c4f089bc9906d8a4cf6fa654fe329085e665|2015-01-10 10:21:00|0|317|35.024464|-80.847383|00000000968840|CAFFE MOCHA GRANDE|96884|NFS BEVERAGE ESPRESSO|1589|NFS STARBUCKS|369|COFFEE SHOP|22|4.15|0.0|1
a9ccb5cfbd8f457a1d9282fdc7c21e0ef9fca622|4|4|35.106477|-80.806073|1.8606360681570644|86602249822946f5c8cb0b597e3fe4d634c95174|2015-01-21 13:06:00|0|372|34.937113|-80.837892|00000000968840|CAFFE MOCHA GRANDE|96884|NFS BEVERAGE ESPRESSO|1589|NFS STARBUCKS|369|COFFEE SHOP|22|4.15|0.0|1
6d1d2cb2cc186dd69ecb186d7aa72a3ac928f990|2|11|35.053394|-80.848528|0.1963563005113332|fb5bd376bebd03845c0635ceab65dd4798b98f40|2014-12-17 08:01:00|0|11|35.053394|-80.848528|00000000968840|CAFFE MOCHA GRANDE|96884|NFS BEVERAGE ESPRESSO|1589|NFS STARBUCKS|369|COFFEE SHOP|22|4.15|0.0|1
dacfdb33b1b94a2fa4414bb4c6446e8798041985|4|372|34.937113|-80.837892|14.940093292018869|03592cd8bc5427696c0c6aafaf993e369d069f20|2014-11-28 11:52:00|0|372|34.937113|-80.837892|00000000968840|CAFFE MOCHA GRANDE|96884|NFS BEVERAGE ESPRESSO|1589|NFS STARBUCKS|369|COFFEE SHOP|22|4.15|0.0|1
d3beed2865aae7921602f2091642da20adeeaf91|1|372|34.937113|-80.837892|0.8949185913142746|b631576e18a5af3a288e2c263fcbb7e779753aad|2015-02-10 14:36:00|0|372|34.937113|-80.837892|00000000968840|CAFFE MOCHA GRANDE|96884|NFS BEVERAGE ESPRESSO|1589|NFS STARBUCKS|369|COFFEE SHOP|22|4.15|0.0|1
b7e1959d2ca6e6b555705aa52fe92d50678b324a|4|274|35.603432|-80.895009|2.0639959800117906|2be1ac835c44c433b83e3a3bedbe83debb8ff5ac|2014-12-03 13:43:00|0|372|34.937113|-80.837892|00000000968840|CAFFE MOCHA GRANDE|96884|NFS BEVERAGE ESPRESSO|1589|NFS STARBUCKS|369|COFFEE SHOP|22|4.15|0.0|1
f7f76beca3f43fd3d06fd6a9d93cb3f39922edbc|1|27|35.037115|-80.8062|0.9424819307990322|b3c60047404cc53643fc533e5e1310861da0a11e|2014-12-13 14:06:00|0|11|35.053394|-80.848528|00000000968840|CAFFE MOCHA GRANDE|96884|NFS BEVERAGE ESPRESSO|1589|NFS STARBUCKS|369|COFFEE SHOP|22|8.3|0.0|2
e6f999a809e5b909ec20ce6f12c989ae63711a38|3|274|35.603432|-80.895009|3.1256013346120737|8acbaedf847f2e75bb2384ab3b187950412c6e05|2014-12-07 15:32:00|0|99|35.585842|-80.875654|00000000970270|VAN BEAN CREME FRAPP GRANDE|97027|NFS BEVERAGE BLEND|1597|NFS STARBUCKS|369|COFFEE SHOP|22|3.75|0.75|1
f2ed46f510e8828137c0f19e29512fbb7bf04fb2|3|99|35.585842|-80.875654|0.4945535443015718|315f38d259be8edeb040e86c60eac73d066d403e|2014-12-07 17:30:00|0|99|35.585842|-80.875654|00000000970270|VAN BEAN CREME FRAPP GRANDE|97027|NFS BEVERAGE BLEND|1597|NFS STARBUCKS|369|COFFEE SHOP|22|3.75|0.75|1
b76e7a1d7578ae3c4386136f595330bccf10c913|4|82|35.03469|-80.97058|6.040628599986319|25237fa90ec9bd3d1673383180c6d3d0b58348c5|2014-09-20 08:09:00|0|372|34.937113|-80.837892|00000000970270|VAN BEAN CREME FRAPP GRANDE|97027|NFS BEVERAGE BLEND|1597|NFS STARBUCKS|369|COFFEE SHOP|22|3.75|0.0|1
752b22ddbe76c42a2060a336efcd5462c3d24567|2|475|35.061685|-80.994596|0.5906819874356365|611269f01fe099d12306e0c9bce08560dee649d6|2014-12-01 10:56:00|0|372|34.937113|-80.837892|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
bfcbbed802139ac7669186d20877dd39482cb698|2|317|35.024464|-80.847383|2.5660420149431684|dd85821bcc59c8416056a69f3edc6befed45f6c4|2015-02-11 12:32:00|0|372|34.937113|-80.837892|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
860719f80abfd06486d232b8a90d277c8bb718da|1|317|35.024464|-80.847383|1.3246660865772504|4df21fd266fe59ac2cce9d4ba667a773857178fe|2014-10-16 14:46:00|0|372|34.937113|-80.837892|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
bfcbbed802139ac7669186d20877dd39482cb698|2|317|35.024464|-80.847383|2.5660420149431684|6471e36a9b0d1225e5e31a9e9c75ee4fafe1b847|2014-11-26 13:11:00|0|372|34.937113|-80.837892|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
81716d206ac9e2fd11f4990c9cc9a400913a8da1|2|372|34.937113|-80.837892|1.5946244690539713|3c78c1ec576716f126b69e3f76895299daa44311|2014-12-30 11:38:00|0|372|34.937113|-80.837892|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
4b763d22f21a9368d026ffce30541832b3d1d92a|4|30|35.096737|-80.78468|1.4696861862856192|8452edf40bdba2f78c971593108f11c57eec0ee3|2014-10-31 06:58:00|0|30|35.096737|-80.78468|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
fcc5d58e9957d711f521538a51cd8e539172b551|2|274|35.603432|-80.895009|0.4783380715738666|b316d2db5fa29f23170f9177c6f942f594f8f239|2015-03-03 14:22:00|0|268|35.500972|-80.860108|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
a3f4cb9e93abd3649c447f33b58f674ae0bf6a11|1|343|35.024332|-80.760919|1.3528897159292559|99378dec980b9d029df1de089c3dafa784490207|2015-01-07 17:19:00|0|343|35.024332|-80.760919|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
02f632f97e6ee0e343457799ff8d03e0c10efc57|3|60|35.006282|-80.562829|1.9508129485108234|16be678b2aed1bcebf29d1929731ed40b0cc94a5|2015-02-17 17:37:00|0|372|34.937113|-80.837892|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
bc2094ce69319750fe453163626c34f5f02ac440|1|317|35.024464|-80.847383|1.9351309237958876|13209104164c837754dc13ee1b0895df2a480bd2|2014-09-16 10:05:00|0|372|34.937113|-80.837892|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
e1b64d50bff78b58d231ac88e6d5a1f63571b2fe|1|182|34.95459|-80.758228|1.6523096976949503|c0b109b112c3e4906af55066340c029698849c65|2015-01-02 10:31:00|0|372|34.937113|-80.837892|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
ac97c9807f4e8ecfd8f521ec71942b189b872c95|4|46|35.28326|-80.66939|2.324395142558342|01075d93ccacff7565ae7ea7d25d293efd12a3e9|2015-02-15 12:34:00|0|157|35.124987|-80.709466|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
47be97d09e0003fbdc415c4bbbb20d3b1600e0cf|1|182|34.95459|-80.758228|2.7365265536039165|6aed5830473b60d2c081ad62fbfc7fa0895184d0|2015-02-16 14:26:00|0|372|34.937113|-80.837892|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
83ef7b48cfb4429025d2c7d9c24bc4b582f21ede|1|401|35.219587|-80.810056|0.674664642588163|77e83977695797905cbae373072f0426faf8e214|2015-01-03 12:06:00|0|401|35.219587|-80.810056|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
07b57d1183af18d93e71704ee187dff4c4860163|3|343|35.024332|-80.760919|1.623728066623682|453c5595d4fa9d79922bb58f30d862f60a16d203|2014-10-23 08:44:00|0|30|35.096737|-80.78468|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
fcc5d58e9957d711f521538a51cd8e539172b551|2|274|35.603432|-80.895009|0.4783380715738666|5bccd11cf82bc01f392acb017dee064d54a8a9b1|2014-10-07 13:33:00|0|268|35.500972|-80.860108|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
17fe33c60414bc1e1fc5eb342c1d9bc156262cf2|4|372|34.937113|-80.837892|15.014266051001554|374557575e792454415e94d407c31dab5ec47fff|2014-11-23 12:53:00|0|372|34.937113|-80.837892|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
af28a45ea9671b5d0a7dc5621443254b6107e505|1|182|34.95459|-80.758228|2.042017111701055|c09afc34d8057e86a8485a0b778c83dd8619d3db|2014-12-04 13:28:00|0|182|34.95459|-80.758228|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
b3f910f1762a90ccc704ed67d5558a0a0053ce17|1|182|34.95459|-80.758228|1.1405793117023135|b83012bb3d7004b432c5f6fd8ce80f09b702c1c3|2015-02-13 10:58:00|0|372|34.937113|-80.837892|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
e152fc2a3d1585d571a3531cf3108082295f0b31|4|30|35.096737|-80.78468|1.3618085366161023|be8f687cee60cd6f7aafa00e99261b27652bb3b7|2014-11-28 10:50:00|0|30|35.096737|-80.78468|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
ab2e0e98191b8e0155bb5afdcc911a1b9c4e2323|3|249|35.000049|-80.699686|1.9093686323325485|442358e5d3d0931872977237a35ed09cd35e0b0a|2014-10-09 09:53:00|0|182|34.95459|-80.758228|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
980185e36467e4c83cbc62b1c25ed702b6ffe667|2|372|34.937113|-80.837892|2.901017493607364|860777f692d2e4d559da9d0da1d4cc534ab73330|2014-10-04 08:38:00|0|372|34.937113|-80.837892|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
fcc5d58e9957d711f521538a51cd8e539172b551|2|274|35.603432|-80.895009|0.4783380715738666|5c18cb922ae8eb4e37c05c61cd7314c175313321|2014-12-17 08:17:00|0|268|35.500972|-80.860108|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
af5041fd5b8afb72759adfccd8c05c691fcab801|1|88|35.103409|-80.992182|2.202236641591022|240334af670831c1ed86f702fd259013a078cd51|2014-11-24 11:05:00|0|372|34.937113|-80.837892|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
bc08fefa4c8ec2cfb689abecbb76d0b0385ab12d|4|372|34.937113|-80.837892|14.384850774435352|fe085aac9a76e6c372ad441d4886bb431f038554|2014-11-18 15:31:00|0|372|34.937113|-80.837892|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|1.2|0.0|2
3e2be403d13acb3d49978546757a7ff908a48183|1|317|35.024464|-80.847383|2.110031931888723|9ca368414c5d9f866da83fa4541e11947e5bc2ef|2015-02-19 10:31:00|0|372|34.937113|-80.837892|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
6d6e6e417c49cf3c26edd0ad4df3c3227f670bf2|1|258|35.297134|-80.737839|1.0331409894584636|5e7eade70f7e8494b1df29d42e3b2605ddecbb0b|2014-12-20 09:32:00|0|258|35.297134|-80.737839|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
b65268f411a4740ecc39ed218be759e498a2e643|2|372|34.937113|-80.837892|4.209072079623996|c42d8acac949f495352d815022514da04db2ae87|2014-12-15 12:05:00|0|11|35.053394|-80.848528|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
5574863a022c4a0e8707b9004a5888e179c899c2|2|372|34.937113|-80.837892|1.524222570844152|434dc3477cf08f3191ac004b284ed2af9c791b66|2014-11-16 13:06:00|0|372|34.937113|-80.837892|00000000970630|ADD SOY|97063|NFS OTHER|1596|NFS STARBUCKS|369|COFFEE SHOP|22|0.6|0.0|1
8c4537928c38b0a42936ae1338f368eb6da6b75b|3|474|35.172688|-80.661096|0.3426118985698578|fecb17e3509565b2ea50197241bcb95605e7ac9e|2015-02-13 08:17:00|0|474|35.172688|-80.661096|00000000971620|TEVANA SPICE CHAI TEA LATTE G|97162|NFS BEVERAGE TEA|1582|NFS STARBUCKS|369|COFFEE SHOP|22|4.25|0.0|1
eeb4393b468b3138577519d2d1297e9cec4fe93b|1|45|35.066546|-80.771677|0.8065745752514656|1d296a8dfc6bbd13e30b6d4d0b87c216d3e2dc88|2015-01-26 16:07:00|0|45|35.066546|-80.771677|00000000971620|TEVANA SPICE CHAI TEA LATTE G|97162|NFS BEVERAGE TEA|1582|NFS STARBUCKS|369|COFFEE SHOP|22|4.25|0.0|1
68437280b0298718c0f0cd146b0ececadc12bae9|2|88|35.103409|-80.992182|3.590689780168165|44ef71df50d562157476483cb12e35f37790a194|2015-01-20 09:04:00|0|372|34.937113|-80.837892|00000000958680|PUMPKIN CREAM CHEESE MUFFINS|95868|PASTRY|1599|STARBUCKS|370|COFFEE SHOP|22|2.45|0.0|1
cd82b0089e475d7674fa91422e3b28311d1bde88|4|372|34.937113|-80.837892|4.253008124100085|20640865fb2f978c903e37c2a65630bb384786cb|2014-10-01 19:02:00|0|372|34.937113|-80.837892|00000000958680|PUMPKIN CREAM CHEESE MUFFINS|95868|PASTRY|1599|STARBUCKS|370|COFFEE SHOP|22|2.45|0.0|1
c76b21dfd0f2c66352dad9d8e62bafc37863b4b3|1|39|35.140781|-80.62331|1.5698730232053706|e0e0761a313939b7a216c3ac0e025571bc5509f4|2014-12-22 12:36:00|0|474|35.172688|-80.661096|00000000959120|PEPPERMNT WHITE CHOC. MOCHA 20|95912|NFS BEVERAGE BLEND|1597|NFS STARBUCKS|369|COFFEE SHOP|22|4.95|0.0|1
9d44568dded8166890c910aecbc70fbb51f36326|2|372|34.937113|-80.837892|5.458647515346652|959e3590cbc276706dcabbc7a4a2b61de2f31755|2015-01-03 08:13:00|0|372|34.937113|-80.837892|00000000969020|ICED WHITE CHOCO MOCHA VENTI|96902|NFS BEVERAGE ESPRESSO|1589|NFS STARBUCKS|369|COFFEE SHOP|22|4.95|0.0|1
b94422871341ac721517e7759e09991de07e4b1d|1|412|35.195689|-80.826724|0.7397863830403285|82e2503b451bf3051332692595122dfb86ce0ea8|2014-11-02 12:34:00|0|160|35.152722|-80.825175|00000772061209|BLAZE FIREFLY FLASHLIGHT|77206120|ALL OTHER TOYS|6450|TOYS|1556|GM|18|9.99|0.0|1
1c8e94670c63d78b3085b11946fa7fee1f84430f|4|121|35.444064|-80.995484|6.517504633353735|64908c459d229d46e467291c1222f60b343177d9|2014-12-22 17:03:00|0|121|35.444064|-80.995484|00000828259307|LADIES KNIT ROCHED GLOVES|82825930|WINTER GLOVES|7221|SEASONAL MERCHANDISE|1600|GM|18|4.99|1.0|1
38f556ebac7b94edea9804feacf92fa9ff1eb5b7|2|190|35.41832|-80.746334|1.13444600562727|8236e26ee710ce561042719a131a310ccded7f51|2015-01-04 08:26:00|0|190|35.41832|-80.746334|00000828259659|MENS KNIT WATCH CAP|82825968|WINTER GLOVES|7221|SEASONAL MERCHANDISE|1600|GM|18|2.99|0.5|1
61c2fea030ac6a1c5bb9ba2f3110567d40563bd5|1|220|35.341927|-80.764523|0.6471599659326277|32d0faabeae6bbf466113289a35ddb7cdb62807c|2014-11-18 07:38:00|0|220|35.341927|-80.764523|00000828259659|MENS KNIT WATCH CAP|82825968|WINTER GLOVES|7221|SEASONAL MERCHANDISE|1600|GM|18|2.99|0.5|1
d19aad74f8fda24ab6c6fd0f220837e38eee30d7|4|208|35.17739|-80.80146|0.9157543917344729|ac0a53a64dd75116253d64cebfb94524fef267d9|2014-11-28 16:48:00|0|167|35.318911|-80.780702|00000828259659|MENS KNIT WATCH CAP|82825968|WINTER GLOVES|7221|SEASONAL MERCHANDISE|1600|GM|18|2.99|0.5|1
9429970f38c1bfb83194d19c473ef1387f3106df|1|30|35.096737|-80.78468|1.2832971912169124|6b1a17d3026d94880130a39ccf6a8a5d0cb5900e|2014-11-16 19:21:00|0|147|35.082768|-80.732725|00000828259758|BOYS INSULATED FLEECE GLOVES|82825975|WINTER GLOVES|7221|SEASONAL MERCHANDISE|1600|GM|18|9.99|1.0|1
de971c00b3f018d18e7aeee56b8ef5ac93cc1993|1|218|35.175855|-80.85013|0.11804675656019406|00b18c8286ece38aa8f7d1fc9d01154298671fca|2015-01-12 15:21:00|0|11|35.053394|-80.848528|00000828259758|BOYS INSULATED FLEECE GLOVES|82825975|WINTER GLOVES|7221|SEASONAL MERCHANDISE|1600|GM|18|9.99|1.0|1
7ab9d203f0b0531f3b5228127bfc91b9d45d324f|1|66|35.059823|-80.816172|2.1670607516204012|6093ebd2ebbc31417951aefb0f852eeecb262f6e|2014-12-20 16:05:00|0|66|35.059823|-80.816172|00008005930025|SWEET POTATO GNOCCHI|800593001|FILLED PASTA|1886|PASTA|440|DELI|6|4.99|0.0|1
fddfe1385dac6e096e26faa4f56d5c63d89ffc47|2|182|34.95459|-80.758228|2.127999222498568|ed773588406b2e3704bc2d5d3b3c98bcb079214e|2014-09-15 15:45:00|0|182|34.95459|-80.758228|00008005930025|SWEET POTATO GNOCCHI|800593001|FILLED PASTA|1886|PASTA|440|DELI|6|4.99|0.0|1
e03e606b1eb253afdbb1fe46d977c6bfd60a9767|1|372|34.937113|-80.837892|3.1453311155349493|fc66f2fc604772943f77f347e528fcccddb82576|2015-01-18 15:03:00|0|27|35.037115|-80.8062|00008005930025|SWEET POTATO GNOCCHI|800593001|FILLED PASTA|1886|PASTA|440|DELI|6|4.99|0.0|1
ba50d6c4bc6c61810fb50285d50af750096deca3|4|122|35.372142|-80.782849|1.5954790766407045|0164cfae280db133a0930e83b5a60207cccaa9b8|2015-02-26 14:34:00|0|122|35.372142|-80.782849|00008005930025|SWEET POTATO GNOCCHI|800593001|FILLED PASTA|1886|PASTA|440|DELI|6|4.99|0.0|1
bf5a342f30c239e16d60c7fdb42e16e2c30e5563|2|82|35.03469|-80.97058|1.4450551659569657|117fe52e945cf6f794f99c20da945ae825017823|2014-10-27 22:47:00|0|82|35.03469|-80.97058|00008005930025|SWEET POTATO GNOCCHI|800593001|FILLED PASTA|1886|PASTA|440|DELI|6|4.99|0.0|1
7598ceb39d25cf64a7775ffc6c9dc4e33359eed8|3|121|35.444064|-80.995484|1.5775944655946195|dfa706808de66938c5a8759b933346adba4b90e3|2015-02-21 17:52:00|0|121|35.444064|-80.995484|00008005930025|SWEET POTATO GNOCCHI|800593001|FILLED PASTA|1886|PASTA|440|DELI|6|4.99|0.0|1
4029e8c40dc895dfafa43d70281e40130c04eab8|2|258|35.297134|-80.737839|0.1681928618912016|405ddc65fe7d3f44a961b4f0aeb75b1879bd06d0|2014-12-04 17:59:00|0|258|35.297134|-80.737839|00008005930025|SWEET POTATO GNOCCHI|800593001|FILLED PASTA|1886|PASTA|440|DELI|6|4.99|0.0|1
93d1e04e16abf71e0f3243fc07463ba928641cf9|4|66|35.059823|-80.816172|1.020415676089764|6431c968c66fdaa0200bfcdd65ee445eb2427b84|2014-12-28 10:43:00|0|66|35.059823|-80.816172|00008100003884|CG CLN SENS SKIN LMU CRM NAT-L|810000388|BRAND-COVER GIRL|3016|COSMETICS|1000|HBC|17|8.79|0.0|1
e07bc0e075e5d474ce3fd580d11db0ee00429565|2|475|35.061685|-80.994596|1.3834652594867658|24a298de1f1bc6fd686b6f9533bc00ca474d25e8|2014-09-12 16:19:00|0|475|35.061685|-80.994596|00008421383511|MINNIE MOUSE BEANIE CLIP|842138330|J HOOK LAMI PROGRAM|6821|J-HOOK|1580|GM|18|4.99|1.0|1
e203ac836840782441ae80837012cce35b5e360e|1|272|35.4437|-80.8955|0.6095109917973324|530348e37c8d17cbc563134db0db60a17e4e7cd6|2015-02-22 12:15:00|0|272|35.4437|-80.8955|00008421411429|I/OBLACK/WHITE RABBIT|842141142|EASTER PLUSH|7050|SEASONAL MERCHANDISE|1600|GM|18|9.99|1.0|1
79dc9328c12e01338bb0d725e4aa4c287d5f1357|3|208|35.17739|-80.80146|1.1109427890835786|83954ece349cc7777a6ba8bc50cf5bced92408ba|2014-11-09 13:12:00|0|208|35.17739|-80.80146|00009125003354|ANDERSON VALLEY BLOOD ORANGE|912500335|CRAFT BEER|458|DOMESTIC BEER|82|BEER|16|10.99|0.0|1
f019a5cc1f13d7413fbb83ff0142530399406b53|2|122|35.372142|-80.782849|0.4667695960651425|32b3bc1118ad81c9704bb6b338e0826aa019679c|2014-12-04 10:27:00|0|122|35.372142|-80.782849|00009281016137|PREVEN'BIG BOOK OF|928101613|MAGAZINES BI-MONTHLY|6788|MAGAZINES|1568|GM|18|10.99|0.0|1
504ab42c956393e7ab2ed8bd358fc9983c21f04a|1|171|35.141204|-80.739|0.49643500805130064|74dbdf713b3b94f2f8fba148949da97938a979a5|2014-12-04 09:06:00|0|157|35.124987|-80.709466|00009281016137|PREVEN'BIG BOOK OF|928101613|MAGAZINES BI-MONTHLY|6788|MAGAZINES|1568|GM|18|10.99|0.0|1
d37e0ac4d603a31edc5d849d402d39302b4d0225|4|182|34.95459|-80.758228|17.085606869705536|7762b060b35b1eeaf53508d9325c3d9b0a6926ae|2014-11-28 20:20:00|0|372|34.937113|-80.837892|00009281028765|TEATIME|928102876|MAGAZINES BI-MONTHLY|6788|MAGAZINES|1568|GM|18|5.99|0.0|1
0bc08d2ed59ac6bb882c1045bbb4a2d7ce7fc4b0|2|129|35.04711|-80.64817|0.8133730718143004|30b4ea3303d61941fc7100a08ee5555b64583da9|2015-01-27 16:38:00|0|129|35.04711|-80.64817|00009281502579|DEER & DEER HUNTIN|928150257|MAGAZINES BI-MONTHLY|6788|MAGAZINES|1568|GM|18|4.99|0.0|1
a1d1ca6476412bceaba4ac36d962a5bbfeab03bd|1|35|35.161696|-80.849471|0.9560219808819127|500829a5061780f0a9678426fe3f3556f342ebeb|2014-11-21 17:22:00|0|218|35.175855|-80.85013|00009300004084|MT OLV JALAPENO SLICES|930000405|PEPPERS|161|PICKLES/OLIVES/RELISHES|25|G1 GROCERY|1|4.49|1.5|1
08c8d8f993178631c524f7b4a410893e5efbb070|2|60|35.006282|-80.562829|15.967537984519032|566ea926b5c24de6088a3db9af952faf47d54d41|2015-02-07 09:47:00|0|60|35.006282|-80.562829|00009300004084|MT OLV JALAPENO SLICES|930000405|PEPPERS|161|PICKLES/OLIVES/RELISHES|25|G1 GROCERY|1|4.49|0.0|1
bb95169b2202a20a3184246788155382d40e9871|1|27|35.037115|-80.8062|0.37155304406119716|f7ea6086dfcf6fc24dd58ad70ed037fde267c8a7|2014-12-24 09:22:00|0|27|35.037115|-80.8062|00009300004084|MT OLV JALAPENO SLICES|930000405|PEPPERS|161|PICKLES/OLIVES/RELISHES|25|G1 GROCERY|1|4.49|0.0|1
ad887550379f3bd0410210e61b5ee732d63545dd|3|160|35.152722|-80.825175|1.181187507595615|5658c5ed31cb408ee76bb20a4d04929c4cd9cae0|2015-03-07 16:40:00|0|160|35.152722|-80.825175|00009300004084|MT OLV JALAPENO SLICES|930000405|PEPPERS|161|PICKLES/OLIVES/RELISHES|25|G1 GROCERY|1|4.49|0.5|1
86f768c3eb414602620b406a4d1574000c931d18|2|46|35.28326|-80.66939|2.2197899361091538|778e191a447c6957732a3d57cd9f2308ab27129e|2015-01-24 12:52:00|0|46|35.28326|-80.66939|00009300004084|MT OLV JALAPENO SLICES|930000405|PEPPERS|161|PICKLES/OLIVES/RELISHES|25|G1 GROCERY|1|4.49|0.0|1
79c737fb93d5bc96ed46ac428bf820ad646cfaf7|1|273|35.06858|-80.7007|1.0690335453483375|3e17dae9b83fe197f6d04bb2fc7477cf2bda0da3|2014-10-10 19:59:00|0|273|35.06858|-80.7007|00009300004084|MT OLV JALAPENO SLICES|930000405|PEPPERS|161|PICKLES/OLIVES/RELISHES|25|G1 GROCERY|1|4.49|0.0|1
642a4e46e1c4e3422b7c51fefec4dc7b7c09726d|1|343|35.024332|-80.760919|1.7616214294321515|92f06f37d328931253cecabcd4bd191c766a4df6|2014-11-11 18:09:00|0|40|35.052812|-80.770346|00009300004084|MT OLV JALAPENO SLICES|930000405|PEPPERS|161|PICKLES/OLIVES/RELISHES|25|G1 GROCERY|1|4.49|0.0|1
19349c088eb2cd43f2326ff2ce539dba6dd3ffc0|1|178|35.667941|-80.497332|6.095754995025354|cfbb1be4b16a665860ffc7c62ee9dfa8ecad13d3|2015-02-14 12:57:00|0|178|35.667941|-80.497332|00009300004084|MT OLV JALAPENO SLICES|930000405|PEPPERS|161|PICKLES/OLIVES/RELISHES|25|G1 GROCERY|1|4.49|0.0|1
87e6ac8869d8262cf130fd7635f428006b93dabe|1|182|34.95459|-80.758228|1.459051272210933|82df8d82c92e9dd6f9c551e63732de4d03fa2c2d|2015-02-16 20:10:00|0|182|34.95459|-80.758228|00009300004084|MT OLV JALAPENO SLICES|930000405|PEPPERS|161|PICKLES/OLIVES/RELISHES|25|G1 GROCERY|1|4.49|0.0|1
ced8f0c24693c24c02a5e87114c62cabf3862b9b|1|66|35.059823|-80.816172|0.8319029642140262|308b74f6bb73a8e982e96fb83a4432e058e33e3a|2015-02-21 16:10:00|0|66|35.059823|-80.816172|00009300004084|MT OLV JALAPENO SLICES|930000405|PEPPERS|161|PICKLES/OLIVES/RELISHES|25|G1 GROCERY|1|4.49|0.0|1
1c1cb70ff84ff398bf5b401708e83cb80d85f779|1|190|35.41832|-80.746334|1.1693425990296873|8ec4184348fa8938bf627bb3747e2cbf86f929a5|2014-10-05 17:14:00|0|190|35.41832|-80.746334|00009300004084|MT OLV JALAPENO SLICES|930000405|PEPPERS|161|PICKLES/OLIVES/RELISHES|25|G1 GROCERY|1|4.49|0.0|1
ebec0fcb0da111560db086b146ce4029291f8a12|3|166|35.323246|-80.945176|1.5799164780019128|b367ce0990c97493bd66ce13c36bb2d571918b61|2015-03-05 10:11:00|0|166|35.323246|-80.945176|00009300004084|MT OLV JALAPENO SLICES|930000405|PEPPERS|161|PICKLES/OLIVES/RELISHES|25|G1 GROCERY|1|4.49|0.5|1
06ac849b03629b6f1971b08f233095c883d3a07d|1|471|35.442529|-80.762919|3.1384540078386265|ecad9445b433448d8a20a9fb505beca65814d498|2014-11-30 17:47:00|0|61|35.204336|-80.844274|00009300004084|MT OLV JALAPENO SLICES|930000405|PEPPERS|161|PICKLES/OLIVES/RELISHES|25|G1 GROCERY|1|4.49|0.0|1
ed0e808f2d6d62d5ad153c62e4c8b8edac290634|1|160|35.152722|-80.825175|1.5263118921543266|eb50ae7789e391ffd42f9f0b2cd9492f0c205963|2015-02-07 13:14:00|0|160|35.152722|-80.825175|00009300004084|MT OLV JALAPENO SLICES|930000405|PEPPERS|161|PICKLES/OLIVES/RELISHES|25|G1 GROCERY|1|4.49|0.0|1
694c1d1e4cb9b3458d6e8fa64f10b4603268804a|2|401|35.219587|-80.810056|0.810296093403428|fb0d74ed73a9cc4a62bd809052c3da2d3843f422|2015-01-15 17:48:00|0|66|35.059823|-80.816172|00009300004084|MT OLV JALAPENO SLICES|930000405|PEPPERS|161|PICKLES/OLIVES/RELISHES|25|G1 GROCERY|1|4.49|0.0|1
b7fca67969aabe5f0d2f0eb2262840e205370814|1|209|35.40953|-80.86175|0.9644142548199185|d0912face65e2550bea3c1283ab3611aad9ca833|2015-01-23 13:32:00|0|272|35.4437|-80.8955|00009300004084|MT OLV JALAPENO SLICES|930000405|PEPPERS|161|PICKLES/OLIVES/RELISHES|25|G1 GROCERY|1|4.49|0.0|1
be79307384fbe74d1c28a1b76e2487bc7bd7198c|1|340|35.444615|-80.861571|1.8498571996604842|9f27cc25f0accb1a076cbd0087128d36430a4732|2015-01-06 12:45:00|0|340|35.444615|-80.861571|00009300004084|MT OLV JALAPENO SLICES|930000405|PEPPERS|161|PICKLES/OLIVES/RELISHES|25|G1 GROCERY|1|4.49|0.0|1
