homeStoreLat|receipt|sales|datetime|tier|mupc|homeStore|LatInt|onlineFlag|Cluster|subcat_num|storeLon|cat_num|storeLat|subcat|discount|dept_num|desc|customer|distance|upc|cat|dept|homeStoreLon|LonInt|store|quantity
35.318911|a92fd4fea4f3ae0c9d1666cb36d5c00208c984da|3.5|2015-02-14 14:50:00|4|20496000000|167|35.365524745616533|0|10|755|-80.945176|87|35.323246|NFS-BALLOONS|0.0|9|*BALLOONS|0bd7d2023e21f25e431ba35c792035d212585811|3.2208980459431045|00204960000005|FLORAL|FLORAL|-80.780702|80.780742074536306|166|1
35.318911|dd38b32a4384aa9d17e415a6a21290eeaf1773ee|10.78|2015-02-16 13:54:00|4|5100015318|167|35.365524637188123|0|32|137|-80.562829|20|35.006282|TOMATO & VEGETABLE JUICE|2.7|1|V8 VEG JUICE 6 PK|0bd7d2023e21f25e431ba35c792035d212585811|3.2208980459431045|00051000153180|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.780702|80.780831606766299|60|2
35.318911|4751d7b132f7126acde8732ae2d343ad7df4c056|10.78|2015-01-29 14:05:00|4|5100017100|167|35.365524637188123|0|32|137|-80.562829|20|35.006282|TOMATO & VEGETABLE JUICE|0.0|1|V8 LS VEG JUICE 6PK|0bd7d2023e21f25e431ba35c792035d212585811|3.2208980459431045|00051000171009|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.780702|80.780831606766299|60|2
35.140781|6627832dba0b2b874fab2b604fa9de3473efda04|2.69|2015-02-13 11:17:00|4|7203663217|39|35.172204825385748|0|37|330|-80.654118|55|35.123768|EGGS|0.69|3|HT GRADE A LARGE EGGS 18 CT|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|00072036632173|EGGS FRESH|DAIRY|-80.62331|80.623322194569553|473|1
35.140781|d7cce5cd02fa38b38359c31fdcb7d87e2188dc4a|8.49|2014-10-02 19:05:00|4|2301290136|39|35.172204825385748|0|37|1477|-80.654118|485|35.123768|SUSHI HYBRID|0.0|6|CRUNCHY ROLL SP|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|00023012901363|SUSHI|DELI|-80.62331|80.623322194569553|473|1
35.140781|0ad8bf5c44b5121e957520c4413a087cd8d07479|8.49|2014-10-11 16:43:00|4|2301290136|39|35.172204826560865|0|11|1477|-80.661096|485|35.172688|SUSHI HYBRID|0.0|6|CRUNCHY ROLL SP|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|00023012901363|SUSHI|DELI|-80.62331|80.623316182353093|474|1
35.140781|1db39fe244060d14edca4ddd6ea6262b1fa5aadf|2.69|2014-10-28 16:04:00|4|7203688023|39|0.6133223301722653|0|8|555|-80.62331|64|35.140781|PACKAGED SALADS|0.0|4|HT CURLY SPINACH,PKG|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|00072036880239|FRESH PRODUCE|PRODUCE|-80.62331|1.4071422133560694|39|1
35.140781|7a761e97f5d26de237b38d0a3cbe0b8bd7153ea9|5.99|2015-02-01 16:40:00|4|7756725423|39|35.172204826560865|0|11|252|-80.661096|45|35.172688|PREMIUM ICE CREAM|1.41|5|BREYERS CHOCOLATE I/C|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|00077567254207|ICE CREAM|FROZEN|-80.62331|80.623316182353093|474|1
35.140781|7f0620c5c7ae010668948eef23a9f6b6e7a1b0a9|6.98|2015-01-13 15:01:00|4||39|35.172204825385748|0|37|500|-80.654118|64|35.123768|FRESH APPLES|0.0|4|GOLD DEL APPLE, WA 56|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|00233285000001|FRESH PRODUCE|PRODUCE|-80.62331|80.623322194569553|473|1
35.140781|d71c322ebbd7a975815d7a703a6f212f422fbd10|3.99|2014-12-22 14:05:00|4|20405400000|39|35.172204826560865|0|11|504|-80.661096|64|35.172688|FRESH BERRIES|0.0|4|RED RASPBERRIES 6 OZ|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|00812049004419|FRESH PRODUCE|PRODUCE|-80.62331|80.623316182353093|474|1
35.140781|fb90fe3a32a33ed7075c88eb3859a7890d21454b|1.89|2014-09-15 20:03:00|4|1300079630|39|0.6133223301722653|0|8|69|-80.62331|26|35.140781|CANNED GRAVY|0.0|1|HEINZ GRAVY BROWN HOMESTYLE|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|00013000798006|PREPARED FOODS-DRY MIXES|G1 GROCERY|-80.62331|1.4071422133560694|39|1
35.140781|bcdde8440dcb26c7c148597894ed18889d76d649|2.69|2014-09-23 14:38:00|4|7203663996|39|35.172204826560865|0|11|342|-80.661096|57|35.172688|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|00072036631299|MILK|DAIRY|-80.62331|80.623316182353093|474|1
35.140781|cd96ef6d0c9f870999de2650839aeeea9d3c714b|2.29|2014-09-23 14:37:00|4|7203695175|39|35.172204826560865|0|11|1607|-80.661096|371|35.172688|FROZEN DOUGH (BREAD)|0.0|14|FRESH LRG FRENCH BREAD|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|00072036951755|BREAD|BAKERY|-80.62331|80.623316182353093|474|1
35.140781|cc5e8eac785379646c0ba80f3e811a985488f6dd|1.49|2014-11-10 16:02:00|4|7203688005|39|0.6133223301722653|0|8|555|-80.62331|64|35.140781|PACKAGED SALADS|0.0|4|HT GARDEN SALAD 16 OZ|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|00072036880055|FRESH PRODUCE|PRODUCE|-80.62331|1.4071422133560694|39|1
35.140781|2e5f997d6485145ad186aa8ad17acc472ce4654c|1.79|2015-02-10 14:26:00|4|7203671215|39|35.172204825385748|0|37|225|-80.654118|35|35.123768|SUGAR-GRANULATED|0.0|1|HT GRANULATED SUGAR|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|00072036712158|SUGAR/SUBSTITUTES|G1 GROCERY|-80.62331|80.623322194569553|473|1
35.03469|fd5c195e0ca73eba9d5d225bf13649737dd66216|6.78|2015-03-03 21:04:00|4|85631200220|82|0.6114706929155321|0|7|97|-80.97058|8|35.03469|ENERGY DRINKS|1.78|23|CORE POWER CHOCOLATE LIGHT|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|00856312002252|CARBONATED BEVERAGES|BEVERAGE|-80.97058|1.4132032182494703|82|2
35.03469|1ba2fbf22f2382740ec0b4d003a72d0e926af1a3|13.58|2014-10-03 16:24:00|4|1200080994|82|0.6114706929155321|0|7|54|-80.97058|8|35.03469|DIET|3.39|23|DT SIERRA MIST FRIDGEMATE|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|00012000810145|CARBONATED BEVERAGES|BEVERAGE|-80.97058|1.4132032182494703|82|2
35.03469|b86bb6f925f3511e8d7081c3ff1777a59ce015c3|6.49|2015-03-05 17:11:00|4|30997757708|82|0.6114706929155321|0|7|3005|-80.97058|1000|35.03469|BRAND-ALMAY|0.0|17|ALM LONGWEAR EMUR PADS 80CT|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|00309975924480|COSMETICS|HBC|-80.97058|1.4132032182494703|82|1
35.03469|1cb8cccc1c5c3f15201c9793a29e6f4da3ee104e|5.98|2014-09-11 19:08:00|4|7203688212|82|35.076192215652235|0|5|555|-80.994596|64|35.061685|PACKAGED SALADS|0.0|4|HT SPRING MIX|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|00072036882127|FRESH PRODUCE|PRODUCE|-80.97058|80.970588755830349|475|2
35.03469|f6c8eaa7e895369110d17e2217d613ed042b89aa|3.94|2015-02-11 16:54:00|4|7203629075|82|0.6114706929155321|0|7|1211|-80.97058|272|35.03469|HISP SALSA/DIPS|0.0|1|HT SALSA MEDIUM|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|00072036290755|HISPANIC PREP. FOODS|G1 GROCERY|-80.97058|1.4132032182494703|82|2
35.03469|63fcc53a9d3507682b2df22c51f9b4cb70d22069|1.99|2015-01-28 17:27:00|4|7127915102|82|0.6114706929155321|0|7|555|-80.97058|64|35.03469|PACKAGED SALADS|0.0|4|F.E. GREEN LEAF SHREDS|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|00071279151021|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|96f7f179b9cc578aa8bdc58b4e8978ccf1faa8a0|4.29|2014-10-10 10:20:00|4|4000031354|82|0.6114706929155321|0|7|727|-80.97058|7|35.03469|SEASONAL CANDY-SINGLE FAC|0.5|1|I/O(H14)M&M MC HALLOWEEN|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|00040000313540|CANDY|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|daab2cbec224e82c999fffcc5fcd79757df87e91|4.49|2015-02-18 17:22:00|4|4400002747|82|0.6114706929155321|0|7|91|-80.97058|13|35.03469|SPRAYED BUTTER CRACKERS|1.49|1|RITZ FRSH STACKS WHOLE WHEAT|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|00044000034832|CRACKERS|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|95dfa10894ef0c17effe983d2470565d02fc9be8|3.49|2014-11-12 16:33:00|4|4812127620|82|0.6114706929155321|0|7|1037|-80.97058|164|35.03469|ENGLISH MUFFINS|0.0|7|THOMAS LITE MULTIGRAIN EM PP|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|00048121276201|BREAKFAST|COMMERCIAL BAKERY|-80.97058|1.4132032182494703|82|1
35.03469|5221527095180cca124ccc31282e5208ea370594|5.7|2014-10-30 18:24:00|4|1800000401|82|0.6114706929155321|0|7|327|-80.97058|54|35.03469|DINNER ROLLS-REFRIGERATED|0.0|3|PILLSBURY CRESCENT ROLLS|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|00018000004010|DOUGH PRODUCTS|DAIRY|-80.97058|1.4132032182494703|82|2
35.03469|e94a547f0084a3c6ea0c5e3e6f98adf49ca31159|3.29|2015-01-06 17:00:00|4|7225091171|82|0.6114706929155321|0|7|1033|-80.97058|163|35.03469|HAMBURGER|0.0|7|NATOWN WHITEWHEAT HAMS|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|00072250911719|BUNS/ROLLS|COMMERCIAL BAKERY|-80.97058|1.4132032182494703|82|1
35.03469|ca1e9d5b0d50c6ee01ef543399f4099cb3ab746b|7.38|2015-01-12 16:47:00|4|7127925101|82|0.6114706929155321|0|7|555|-80.97058|64|35.03469|PACKAGED SALADS|0.0|4|F.E. SWEET BUTTER|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|00071279221038|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|2
35.03469|bb24a037ad67f3a4fdc8243f7ad251bb78a1c49e|11.07|2014-12-19 14:43:00|4|7127925101|82|0.6114706929155321|0|7|555|-80.97058|64|35.03469|PACKAGED SALADS|0.0|4|F.E. SWEET BUTTER|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|00071279221038|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|3
35.03469|dd287d77e524c1cdcaae0b4adf07d7f148a8494a|3.99|2014-12-29 20:08:00|4|2301290032|82|0.6114706929155321|0|7|1487|-80.97058|485|35.03469|SUSHI APPETIZERS|0.0|6|dumplings|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|00023012900328|SUSHI|DELI|-80.97058|1.4132032182494703|82|1
35.341927|d0cc4dbd03e9a3cfb10d9f70f56c2aa305d7cc31|4.69|2014-09-20 18:34:00|4|1600043779|220|35.383490730525274|0|6|1433|-80.605588|9|35.43259|GRANOLA|0.0|1|NV PROTEIN GRANOLA OATS HONEY|13f1ef39385226d7fb218594ad6647929f83128a|2.8719573987198292|00016000437791|CEREAL|G1 GROCERY|-80.764523|80.764607981189812|202|1
35.06858|f5272fd0f25ec2668eadc6d467d8b106c17ce827|6.79|2015-01-06 19:15:00|4|1200080994|273|0.612062184999033|0|9|55|-80.7007|8|35.06858|REGULAR|6.79|23|PEPSI FRIDGEMATE|1491831ee4d196c82983355845a5c9a99d794e89|1.1377023968546804|00012000809941|CARBONATED BEVERAGES|BEVERAGE|-80.7007|1.4084929236641879|273|1
35.06858|14f8817799cf0235ed39b882dd820f5dca0a8b4d|6.49|2014-10-28 11:38:00|4|1200080994|273|0.612062184999033|0|9|55|-80.7007|8|35.06858|REGULAR|6.49|23|PEPSI FRIDGEMATE|1491831ee4d196c82983355845a5c9a99d794e89|1.1377023968546804|00012000809941|CARBONATED BEVERAGES|BEVERAGE|-80.7007|1.4084929236641879|273|1
35.06858|7dece82219d67af550e4797d73bff578f273b9d0|9.99|2014-09-16 19:45:00|4|85877000246|273|0.612062184999033|0|9|458|-80.7007|82|35.06858|CRAFT BEER|0.0|16|OMB CHRISTMAS 12OZ 6PACK|1491831ee4d196c82983355845a5c9a99d794e89|1.1377023968546804|00858770002461|DOMESTIC BEER|BEER|-80.7007|1.4084929236641879|273|1
35.06858|a590e01007e2570a9888ec76fd2cda37bdec24cb|13.99|2014-09-19 19:51:00|4|86787200002|273|35.0850451503984|0|4|458|-80.699909|82|35.002628|CRAFT BEER|0.0|16|THE UNKNOWN VEHOPCIRAPTOR 22OZ|1491831ee4d196c82983355845a5c9a99d794e89|1.1377023968546804|00867872000022|DOMESTIC BEER|BEER|-80.7007|80.700713764055649|477|1
35.06858|5332ace6beabe16be86385eed3022df03b9b24fd|3.58|2014-10-25 10:00:00|4|4850001775|273|35.085045141086376|0|12|338|-80.661096|56|35.172688|OTHER FRUIT JUICES|1.58|3|TROPICANA RASP LEMONADE 12 OZ|1491831ee4d196c82983355845a5c9a99d794e89|1.1377023968546804|00048500021545|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.7007|80.700725442152319|474|2
35.059823|cfdbe030802581fb1a3d6077810473919a0dc7d2|5.35|2014-12-04 15:06:00|2|3700041759|66|35.068745252339973|0|0|388|-80.771677|66|35.066546|NFS-DISHWASH PWDR/LIQUID|1.06|1|CASCADE PAC CITRUS BRZ 15CT|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00037000806288|DETERGENTS|G1 GROCERY|-80.816172|80.816174955839742|45|1
35.059823|481f55220f0ba5e39c264bf8db8e4c43605236b0|4.49|2014-12-26 14:40:00|2|4000031532|66|35.068745252587782|0|0|727|-80.770346|7|35.052812|SEASONAL CANDY-SINGLE FAC|2.25|1|I/O(C14)M&M PLAIN CHRISTMAS|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00040000315322|CANDY|G1 GROCERY|-80.816172|80.816173461718321|40|1
35.059823|8c54796945a035791c43643a1534520bae7e43ec|2.99|2014-10-23 16:21:00|2|4145811704|66|35.068745252504428|0|0|265|-80.8062|307|35.037115|FROZEN PIES|0.0|5|EDWARDS CHOC SUNDAE SINGLES|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00041458117049|DESSERTS FROZEN|FROZEN|-80.816172|80.816174087217505|27|1
35.059823|3172d7bc90997eaefac7568b659971209539790e|5.79|2014-10-30 17:07:00|2|4440015600|66|35.068745252504428|0|0|293|-80.8062|48|35.037115|FROZEN SEAFOOD|2.79|5|GORTON'S 18CT FISHSTICKS|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00044400156509|FROZEN MEALS|FROZEN|-80.816172|80.816174087217505|27|1
35.059823|0b80da770f9605ed8bcaba64d0618cb515ca81c9|2.99|2014-09-25 16:23:00|2|4145811704|66|35.068745252504428|0|0|265|-80.8062|307|35.037115|FROZEN PIES|0.0|5|EDWARDS CHOC SUNDAE SINGLES|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00041458117049|DESSERTS FROZEN|FROZEN|-80.816172|80.816174087217505|27|1
35.059823|5b022333e709df5ca39f4208307e1e1bc5e71a2c|2.99|2014-11-13 16:03:00|2|4145811704|66|35.068745252504428|0|0|265|-80.8062|307|35.037115|FROZEN PIES|0.49|5|EDWARDS CHOC SUNDAE SINGLES|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00041458117049|DESSERTS FROZEN|FROZEN|-80.816172|80.816174087217505|27|1
35.059823|622f444a9157095cd052fc272cb33a731af69b2c|4.69|2014-12-26 14:40:00|2|4900002468|66|35.068745252587782|0|0|54|-80.770346|8|35.052812|DIET|1.19|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816173461718321|40|1
35.059823|935f9e083d5cf85225e0e8fc13a3e1b990826cfa|4.99|2015-02-12 16:14:00|2|4900002468|66|35.068745252504428|0|0|54|-80.8062|8|35.037115|DIET|1.0|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|1
35.059823|e5b074bf54ff7f3f28defe12fdc5dde9a0460968|4.99|2015-03-07 16:34:00|2|4900002468|66|35.068745252504428|0|0|54|-80.8062|8|35.037115|DIET|2.49|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|1
35.059823|25c629b14caf361cad0b70cd1b29ec64815d7d31|4.99|2015-01-15 15:57:00|2|4900002468|66|35.068745252504428|0|0|54|-80.8062|8|35.037115|DIET|2.5|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|1
35.059823|3f632921037688c2788a75fefd64838d3bb49e8a|4.99|2015-02-05 17:20:00|2|4900002468|66|35.068745252504428|0|0|54|-80.8062|8|35.037115|DIET|0.0|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|1
35.059823|f923ca73fd50afa8c12bdc1a681b2f156e73db1a|4.99|2015-01-01 15:04:00|2|4900002468|66|35.068745252339973|0|0|54|-80.771677|8|35.066546|DIET|1.0|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174955839742|45|1
35.059823|41c5da2906840bd780a72ec471e02f29fc7c40d3|4.69|2014-09-18 15:59:00|2|4900002468|66|35.068745252504428|0|0|54|-80.8062|8|35.037115|DIET|1.19|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|1
35.059823|e93870e45b839ecd6725983f1b980a0abdd8066c|4.69|2014-10-16 16:42:00|2|4900002468|66|0.6119093465164359|0|1|54|-80.816172|8|35.059823|DIET|0.0|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|1.4105082902580508|66|1
35.059823|53fc38435cfb362610cf3f291abac4f0be19a3be|4.69|2014-09-11 15:37:00|2|4900002468|66|35.068745252504428|0|0|54|-80.8062|8|35.037115|DIET|2.35|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|1
35.059823|487a33d65619150a87eb2f4b923ff928298cef22|4.69|2014-10-09 15:35:00|2|4900002468|66|35.068745252587782|0|0|54|-80.770346|8|35.052812|DIET|1.19|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816173461718321|40|1
35.059823|f9928f5d9957385f9899ad529196811e03268cd9|4.99|2015-02-25 12:00:00|2|4900002468|66|0.6119093465164359|0|1|54|-80.816172|8|35.059823|DIET|1.0|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|1.4105082902580508|66|1
35.059823|e916dab4a93fe339a082e901a05e722bfbe6a0cf|4.99|2015-02-19 16:10:00|2|4900002468|66|35.068745252504428|0|0|54|-80.8062|8|35.037115|DIET|2.5|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|1
35.059823|a13af3a3c3f8761e2630277d87b0a148fbccb8e5|4.69|2014-11-06 15:29:00|2|4900002468|66|35.068745252504428|0|0|54|-80.8062|8|35.037115|DIET|2.35|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|1
35.059823|c9c44524b63a6a286394cedd2ac5370d044a9f77|4.69|2014-12-18 15:59:00|2|4900002468|66|35.068745252504428|0|0|54|-80.8062|8|35.037115|DIET|1.19|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|1
35.059823|dc407dc526d87fc4c3ff6552da79a8ddf340a261|4.99|2015-01-08 15:52:00|2|4900002468|66|0.6119093465164359|0|1|54|-80.816172|8|35.059823|DIET|0.0|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|1.4105082902580508|66|1
35.059823|ac81691df00af01395105016df2815bf34a0e03a|9.38|2014-11-28 15:49:00|2|4900002468|66|35.068745252504428|0|0|54|-80.8062|8|35.037115|DIET|5.44|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|2
35.059823|cade03f00e3c2c06d93f53a2d8424f795d8251cb|4.69|2014-10-02 15:31:00|2|4900002468|66|35.068745252504428|0|0|54|-80.8062|8|35.037115|DIET|2.35|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|1
35.059823|45596165a660d6a528890874089ecafba6a53e99|4.69|2014-12-12 14:56:00|2|4900002468|66|35.068745252504428|0|0|54|-80.8062|8|35.037115|DIET|0.0|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|1
35.059823|801fb635b52c42649dd83315ae304ceb692a20fe|1.25|2015-01-22 16:16:00|2|4850001775|66|35.068745252504428|0|0|335|-80.8062|56|35.037115|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA PP ORIGINAL 12 OZ|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00048500017753|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.816172|80.816174087217505|27|1
35.059823|8e827d9d2d3b01e39276895351e0f7d21701bf8d|1.79|2014-10-25 16:34:00|2|4850001775|66|35.068745252339973|0|0|335|-80.771677|56|35.066546|ORANGE JUICE-REGRIGERATED|0.79|3|TROPICANA PP ORIGINAL 12 OZ|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00048500017753|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.816172|80.816174955839742|45|1
35.059823|917df65f81e48d99efd5338719fdd1661aa44db2|3.49|2014-12-11 16:14:00|2|7017715419|66|0.6119093465164359|0|1|233|-80.816172|37|35.059823|BLACK TEA|0.49|1|TWININGS DECAF EARL GREY|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00070177171674|TEA|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|866303475f5ca16c23095e253bc37def65f60809|4.23|2015-01-29 16:11:00|2||66|0.6119093465164359|0|1|529|-80.816172|64|35.059823|FRESH ASPARAGUS|2.12|4|GREEN  ASPARAGUS|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00204080000008|FRESH PRODUCE|PRODUCE|-80.816172|1.4105082902580508|66|1
35.059823|021dbee4854f83c9251e5f4db005786edb9941bc|8.98|2014-10-03 14:52:00|2|4164120104|66|35.068745252504428|0|0|899|-80.8062|205|35.037115|KOSHER FROZEN FOODS|0.0|5|GOLDEN PANCAKE POTATO|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00041641201036|FROZEN KOSHER|FROZEN|-80.816172|80.816174087217505|27|2
35.059823|87682e44f8d4e136b1786dc181a835fb84f2593e|12.35|2014-09-21 11:31:00|2|20598600000|66|35.068745252603684|0|0|1800|-80.760919|400|35.024332|FFM BEEF|0.0|6|HT ROAST  BEEF|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00205986000000|FFM MEAT|DELI|-80.816172|80.816173308875435|343|1
35.059823|86e9e285566b0d3191f696aa30c739a544da526c|1.77|2014-10-05 16:03:00|2|7203614049|66|35.068745252465455|0|0|104|-80.848528|16|35.053394|APPLESAUCE-CUPS|0.5|1|HT APPLESAUCE 6PK UNSWTND|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00072036140494|FRUIT-CAN/JAR|G1 GROCERY|-80.816172|80.816174322633771|11|1
35.059823|1de4a13ddefc7b0b0d03141d0f41948ddfd5f80e|3.99|2014-10-18 14:09:00|2|4000015140|66|35.068745252339973|0|0|46|-80.771677|7|35.066546|PKG CHOC|0.49|1|3 MUSKETEER FUN SIZE|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00040000151227|CANDY|G1 GROCERY|-80.816172|80.816174955839742|45|1
35.059823|790e64096132535ebf41d5620c82a93c562d7ee9|9.99|2014-09-13 14:29:00|2|4200044517|66|35.068745252339973|0|0|426|-80.771677|72|35.066546|NFS-PAPER TOWELS|3.0|1|BRAWNY 6 BIG ROLL PICK A SIZE|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00042000445177|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.816172|80.816174955839742|45|1
35.059823|b3d125ffa7fba9e294c372063ba80325d57c1cb2|4.49|2014-11-20 16:03:00|2|8265700312|66|35.068745252504428|0|0|31|-80.8062|4|35.037115|NON CARBONATED WATER|0.5|1|DEER PARK SPRG WATER .5 LTR|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00082657003122|BOTTLED WATER|G1 GROCERY|-80.816172|80.816174087217505|27|1
35.059823|3ef0637ae68418909a6b437732fa44389c0dd508|4.99|2015-01-24 16:35:00|2|8265750406|66|35.068745252339973|0|0|31|-80.771677|4|35.066546|NON CARBONATED WATER|1.49|1|(U)DEER PARK WATER 24PK .5LT|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00082657504063|BOTTLED WATER|G1 GROCERY|-80.816172|80.816174955839742|45|1
35.059823|7aab3718533712bf9522bb616f528effed1449f6|4.99|2015-02-15 15:19:00|2|8265750406|66|35.068745252339973|0|0|31|-80.771677|4|35.066546|NON CARBONATED WATER|0.5|1|(U)DEER PARK WATER 24PK .5LT|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00082657504063|BOTTLED WATER|G1 GROCERY|-80.816172|80.816174955839742|45|1
35.059823|6e5658a3ce89334d76e17e4791b7dfbf29079a77|2.89|2015-02-16 14:02:00|2|7203655029|66|0.6119093465164359|0|1|331|-80.816172|52|35.059823|NATURAL SLICED|1.22|3|HT RF PEPPER JACK SLICES|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00072036708694|CHEESE|DAIRY|-80.816172|1.4105082902580508|66|1
35.059823|549e7d818532d1e73b8ee1a6260ce500766289a7|2.19|2015-03-03 16:10:00|2|2880000001|66|0.6119093465164359|0|1|247|-80.816172|39|35.059823|VEGETABLES-FLANKER|0.0|1|HANOVER THREE BEAN SALAD|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00028800000013|VEGETABLES-CAN/JAR|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|e4402817c3ea7d62227503bf6120713ad3e30106|3.99|2014-12-24 16:21:00|2|88810911004|66|35.068745252339973|0|0|1046|-80.771677|173|35.066546|CAKES|2.0|7|HOSTESS CINN COFFEE CAKE|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00888109110048|SWEET BAKED GOODS|COMMERCIAL BAKERY|-80.816172|80.816174955839742|45|1
35.059823|dfdcd5a7d0f5fe83b0f037f0a9c0929f17e80636|4.99|2015-01-15 15:57:00|2|7099210227|66|35.068745252504428|0|0|6785|-80.8062|1568|35.037115|MAGAZINES WEEKLY|0.0|18|10227 PEOPLE|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00070992102273|MAGAZINES|GM|-80.816172|80.816174087217505|27|1
35.059823|d84c45cad2c021a1b19f3b50000d6cf3236ecff0|3.99|2015-02-12 16:11:00|2|4000042065|66|35.068745252504428|0|0|46|-80.8062|7|35.037115|PKG CHOC|1.99|1|I/O MM MILK CHOCOLATE BONUS|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00040000420651|CANDY|G1 GROCERY|-80.816172|80.816174087217505|27|1
35.059823|3042258cb06d2b5032a313ef80db5d508a48ba36|1.79|2014-10-21 14:47:00|2|2500000024|66|35.068745252504428|0|0|335|-80.8062|56|35.037115|ORANGE JUICE-REGRIGERATED|0.0|3|SIMPLY ORANGE JUICE PULP FREE|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00025000000249|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.816172|80.816174087217505|27|1
35.059823|701cf16ae1e93fe88a5be525e26ef64c4e7bdac3|2.79|2015-02-25 12:02:00|2|1130038110|66|0.6119093465164359|0|1|50|-80.816172|7|35.059823|PEG CANDY|0.0|1|BRACHS LEMON DROPS|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00011300384011|CANDY|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|7a5c1ae07f860411440819cd56b746420c75038f|2.79|2014-12-18 15:55:00|2|1130038110|66|35.068745252504428|0|0|50|-80.8062|7|35.037115|PEG CANDY|0.0|1|BRACHS LEMON DROPS|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00011300384011|CANDY|G1 GROCERY|-80.816172|80.816174087217505|27|1
35.059823|6da4ebebc76635a0baea9d47d5f2d9b407ff4bf1|2.79|2015-01-29 16:09:00|2|1130038110|66|0.6119093465164359|0|1|50|-80.816172|7|35.059823|PEG CANDY|0.0|1|BRACHS LEMON DROPS|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00011300384011|CANDY|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|92b638c2b775418722cce4a0016b197b1c2340a9|2.79|2015-01-01 15:05:00|2|1130038110|66|35.068745252339973|0|0|50|-80.771677|7|35.066546|PEG CANDY|0.0|1|BRACHS LEMON DROPS|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00011300384011|CANDY|G1 GROCERY|-80.816172|80.816174955839742|45|1
35.059823|059e1ac4ee3a32925e546231762fca8ec19e6d16|2.79|2015-01-08 15:53:00|2|1130038110|66|0.6119093465164359|0|1|50|-80.816172|7|35.059823|PEG CANDY|0.0|1|BRACHS LEMON DROPS|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00011300384011|CANDY|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|c85cdd0907d392574d365d1afab49d2f808624a2|2.79|2015-02-19 16:07:00|2|1130038110|66|35.068745252504428|0|0|50|-80.8062|7|35.037115|PEG CANDY|0.0|1|BRACHS LEMON DROPS|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00011300384011|CANDY|G1 GROCERY|-80.816172|80.816174087217505|27|1
35.059823|63025eaccedfdebca98d440d3802169a8d06cf5c|2.79|2015-03-07 16:29:00|2|1130038110|66|35.068745252504428|0|0|50|-80.8062|7|35.037115|PEG CANDY|0.0|1|BRACHS LEMON DROPS|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|00011300384011|CANDY|G1 GROCERY|-80.816172|80.816174087217505|27|1
