homeStoreLat|receipt|sales|datetime|z_CenLon|tier|mupc|homeStore|LatInt|onlineFlag|Cluster|subcat_num|storeLon|cat_num|storeLat|subcat|discount|dept_num|desc|customer|distance|z_CenLat|upc|cat|dept|homeStoreLon|LonInt|store|quantity
35.318911|a92fd4fea4f3ae0c9d1666cb36d5c00208c984da|3.5|2015-02-14 14:50:00|80.780380710856576|4|20496000000|167|35.365524745616533|0|48|755|-80.945176|87|35.323246|NFS-BALLOONS|0.0|9|*BALLOONS|0bd7d2023e21f25e431ba35c792035d212585811|3.2208980459431045|35.351085445956379|00204960000005|FLORAL|FLORAL|-80.780702|80.780742074536306|166|1
35.318911|dd38b32a4384aa9d17e415a6a21290eeaf1773ee|10.78|2015-02-16 13:54:00|80.780380710856576|4|5100015318|167|35.365524637188123|0|48|137|-80.562829|20|35.006282|TOMATO & VEGETABLE JUICE|2.7|1|V8 VEG JUICE 6 PK|0bd7d2023e21f25e431ba35c792035d212585811|3.2208980459431045|35.351085445956379|00051000153180|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.780702|80.780831606766299|60|2
35.318911|4751d7b132f7126acde8732ae2d343ad7df4c056|10.78|2015-01-29 14:05:00|80.780380710856576|4|5100017100|167|35.365524637188123|0|48|137|-80.562829|20|35.006282|TOMATO & VEGETABLE JUICE|0.0|1|V8 LS VEG JUICE 6PK|0bd7d2023e21f25e431ba35c792035d212585811|3.2208980459431045|35.351085445956379|00051000171009|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.780702|80.780831606766299|60|2
35.140781|6627832dba0b2b874fab2b604fa9de3473efda04|2.69|2015-02-13 11:17:00|80.632521683083056|4|7203663217|39|35.172204825385748|0|39|330|-80.654118|55|35.123768|EGGS|0.69|3|HT GRADE A LARGE EGGS 18 CT|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|35.177497916598789|00072036632173|EGGS FRESH|DAIRY|-80.62331|80.623322194569553|473|1
35.140781|d7cce5cd02fa38b38359c31fdcb7d87e2188dc4a|8.49|2014-10-02 19:05:00|80.632521683083056|4|2301290136|39|35.172204825385748|0|39|1477|-80.654118|485|35.123768|SUSHI HYBRID|0.0|6|CRUNCHY ROLL SP|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|35.177497916598789|00023012901363|SUSHI|DELI|-80.62331|80.623322194569553|473|1
35.140781|0ad8bf5c44b5121e957520c4413a087cd8d07479|8.49|2014-10-11 16:43:00|80.632521683083056|4|2301290136|39|35.172204826560865|0|39|1477|-80.661096|485|35.172688|SUSHI HYBRID|0.0|6|CRUNCHY ROLL SP|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|35.177497916598789|00023012901363|SUSHI|DELI|-80.62331|80.623316182353093|474|1
35.140781|1db39fe244060d14edca4ddd6ea6262b1fa5aadf|2.69|2014-10-28 16:04:00|1.4091206135396188|4|7203688023|39|0.6133223301722653|0|47|555|-80.62331|64|35.140781|PACKAGED SALADS|0.0|4|HT CURLY SPINACH,PKG|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|0.61242566243833529|00072036880239|FRESH PRODUCE|PRODUCE|-80.62331|1.4071422133560694|39|1
35.140781|7a761e97f5d26de237b38d0a3cbe0b8bd7153ea9|5.99|2015-02-01 16:40:00|80.632521683083056|4|7756725423|39|35.172204826560865|0|39|252|-80.661096|45|35.172688|PREMIUM ICE CREAM|1.41|5|BREYERS CHOCOLATE I/C|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|35.177497916598789|00077567254207|ICE CREAM|FROZEN|-80.62331|80.623316182353093|474|1
35.140781|7f0620c5c7ae010668948eef23a9f6b6e7a1b0a9|6.98|2015-01-13 15:01:00|80.632521683083056|4||39|35.172204825385748|0|39|500|-80.654118|64|35.123768|FRESH APPLES|0.0|4|GOLD DEL APPLE, WA 56|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|35.177497916598789|00233285000001|FRESH PRODUCE|PRODUCE|-80.62331|80.623322194569553|473|1
35.140781|d71c322ebbd7a975815d7a703a6f212f422fbd10|3.99|2014-12-22 14:05:00|80.632521683083056|4|20405400000|39|35.172204826560865|0|39|504|-80.661096|64|35.172688|FRESH BERRIES|0.0|4|RED RASPBERRIES 6 OZ|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|35.177497916598789|00812049004419|FRESH PRODUCE|PRODUCE|-80.62331|80.623316182353093|474|1
35.140781|fb90fe3a32a33ed7075c88eb3859a7890d21454b|1.89|2014-09-15 20:03:00|1.4091206135396188|4|1300079630|39|0.6133223301722653|0|47|69|-80.62331|26|35.140781|CANNED GRAVY|0.0|1|HEINZ GRAVY BROWN HOMESTYLE|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|0.61242566243833529|00013000798006|PREPARED FOODS-DRY MIXES|G1 GROCERY|-80.62331|1.4071422133560694|39|1
35.140781|bcdde8440dcb26c7c148597894ed18889d76d649|2.69|2014-09-23 14:38:00|80.632521683083056|4|7203663996|39|35.172204826560865|0|39|342|-80.661096|57|35.172688|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|35.177497916598789|00072036631299|MILK|DAIRY|-80.62331|80.623316182353093|474|1
35.140781|cd96ef6d0c9f870999de2650839aeeea9d3c714b|2.29|2014-09-23 14:37:00|80.632521683083056|4|7203695175|39|35.172204826560865|0|39|1607|-80.661096|371|35.172688|FROZEN DOUGH (BREAD)|0.0|14|FRESH LRG FRENCH BREAD|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|35.177497916598789|00072036951755|BREAD|BAKERY|-80.62331|80.623316182353093|474|1
35.140781|cc5e8eac785379646c0ba80f3e811a985488f6dd|1.49|2014-11-10 16:02:00|1.4091206135396188|4|7203688005|39|0.6133223301722653|0|47|555|-80.62331|64|35.140781|PACKAGED SALADS|0.0|4|HT GARDEN SALAD 16 OZ|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|0.61242566243833529|00072036880055|FRESH PRODUCE|PRODUCE|-80.62331|1.4071422133560694|39|1
35.140781|2e5f997d6485145ad186aa8ad17acc472ce4654c|1.79|2015-02-10 14:26:00|80.632521683083056|4|7203671215|39|35.172204825385748|0|39|225|-80.654118|35|35.123768|SUGAR-GRANULATED|0.0|1|HT GRANULATED SUGAR|0bf5dbf84014428eb44a49f7818f7ee9eb4e1869|2.1713105576209735|35.177497916598789|00072036712158|SUGAR/SUBSTITUTES|G1 GROCERY|-80.62331|80.623322194569553|473|1
35.03469|fd5c195e0ca73eba9d5d225bf13649737dd66216|6.78|2015-03-03 21:04:00|1.4132775322775095|4|85631200220|82|0.6114706929155321|0|58|97|-80.97058|8|35.03469|ENERGY DRINKS|1.78|23|CORE POWER CHOCOLATE LIGHT|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|0.61177642288969325|00856312002252|CARBONATED BEVERAGES|BEVERAGE|-80.97058|1.4132032182494703|82|2
35.03469|1ba2fbf22f2382740ec0b4d003a72d0e926af1a3|13.58|2014-10-03 16:24:00|1.4132775322775095|4|1200080994|82|0.6114706929155321|0|58|54|-80.97058|8|35.03469|DIET|3.39|23|DT SIERRA MIST FRIDGEMATE|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|0.61177642288969325|00012000810145|CARBONATED BEVERAGES|BEVERAGE|-80.97058|1.4132032182494703|82|2
35.03469|b86bb6f925f3511e8d7081c3ff1777a59ce015c3|6.49|2015-03-05 17:11:00|1.4132775322775095|4|30997757708|82|0.6114706929155321|0|58|3005|-80.97058|1000|35.03469|BRAND-ALMAY|0.0|17|ALM LONGWEAR EMUR PADS 80CT|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|0.61177642288969325|00309975924480|COSMETICS|HBC|-80.97058|1.4132032182494703|82|1
35.03469|1cb8cccc1c5c3f15201c9793a29e6f4da3ee104e|5.98|2014-09-11 19:08:00|80.970590786568081|4|7203688212|82|35.076192215652235|0|55|555|-80.994596|64|35.061685|PACKAGED SALADS|0.0|4|HT SPRING MIX|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|35.077427448337218|00072036882127|FRESH PRODUCE|PRODUCE|-80.97058|80.970588755830349|475|2
35.03469|f6c8eaa7e895369110d17e2217d613ed042b89aa|3.94|2015-02-11 16:54:00|1.4132775322775095|4|7203629075|82|0.6114706929155321|0|58|1211|-80.97058|272|35.03469|HISP SALSA/DIPS|0.0|1|HT SALSA MEDIUM|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|0.61177642288969325|00072036290755|HISPANIC PREP. FOODS|G1 GROCERY|-80.97058|1.4132032182494703|82|2
35.03469|63fcc53a9d3507682b2df22c51f9b4cb70d22069|1.99|2015-01-28 17:27:00|1.4132775322775095|4|7127915102|82|0.6114706929155321|0|58|555|-80.97058|64|35.03469|PACKAGED SALADS|0.0|4|F.E. GREEN LEAF SHREDS|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|0.61177642288969325|00071279151021|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|96f7f179b9cc578aa8bdc58b4e8978ccf1faa8a0|4.29|2014-10-10 10:20:00|1.4132775322775095|4|4000031354|82|0.6114706929155321|0|58|727|-80.97058|7|35.03469|SEASONAL CANDY-SINGLE FAC|0.5|1|I/O(H14)M&M MC HALLOWEEN|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|0.61177642288969325|00040000313540|CANDY|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|daab2cbec224e82c999fffcc5fcd79757df87e91|4.49|2015-02-18 17:22:00|1.4132775322775095|4|4400002747|82|0.6114706929155321|0|58|91|-80.97058|13|35.03469|SPRAYED BUTTER CRACKERS|1.49|1|RITZ FRSH STACKS WHOLE WHEAT|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|0.61177642288969325|00044000034832|CRACKERS|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|95dfa10894ef0c17effe983d2470565d02fc9be8|3.49|2014-11-12 16:33:00|1.4132775322775095|4|4812127620|82|0.6114706929155321|0|58|1037|-80.97058|164|35.03469|ENGLISH MUFFINS|0.0|7|THOMAS LITE MULTIGRAIN EM PP|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|0.61177642288969325|00048121276201|BREAKFAST|COMMERCIAL BAKERY|-80.97058|1.4132032182494703|82|1
35.03469|5221527095180cca124ccc31282e5208ea370594|5.7|2014-10-30 18:24:00|1.4132775322775095|4|1800000401|82|0.6114706929155321|0|58|327|-80.97058|54|35.03469|DINNER ROLLS-REFRIGERATED|0.0|3|PILLSBURY CRESCENT ROLLS|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|0.61177642288969325|00018000004010|DOUGH PRODUCTS|DAIRY|-80.97058|1.4132032182494703|82|2
35.03469|e94a547f0084a3c6ea0c5e3e6f98adf49ca31159|3.29|2015-01-06 17:00:00|1.4132775322775095|4|7225091171|82|0.6114706929155321|0|58|1033|-80.97058|163|35.03469|HAMBURGER|0.0|7|NATOWN WHITEWHEAT HAMS|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|0.61177642288969325|00072250911719|BUNS/ROLLS|COMMERCIAL BAKERY|-80.97058|1.4132032182494703|82|1
35.03469|ca1e9d5b0d50c6ee01ef543399f4099cb3ab746b|7.38|2015-01-12 16:47:00|1.4132775322775095|4|7127925101|82|0.6114706929155321|0|58|555|-80.97058|64|35.03469|PACKAGED SALADS|0.0|4|F.E. SWEET BUTTER|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|0.61177642288969325|00071279221038|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|2
35.03469|bb24a037ad67f3a4fdc8243f7ad251bb78a1c49e|11.07|2014-12-19 14:43:00|1.4132775322775095|4|7127925101|82|0.6114706929155321|0|58|555|-80.97058|64|35.03469|PACKAGED SALADS|0.0|4|F.E. SWEET BUTTER|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|0.61177642288969325|00071279221038|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|3
35.03469|dd287d77e524c1cdcaae0b4adf07d7f148a8494a|3.99|2014-12-29 20:08:00|1.4132775322775095|4|2301290032|82|0.6114706929155321|0|58|1487|-80.97058|485|35.03469|SUSHI APPETIZERS|0.0|6|dumplings|12f1e227f4b1ae744197fb1aeb73ee7dda981544|2.8677029200726714|0.61177642288969325|00023012900328|SUSHI|DELI|-80.97058|1.4132032182494703|82|1
35.341927|d0cc4dbd03e9a3cfb10d9f70f56c2aa305d7cc31|4.69|2014-09-20 18:34:00|80.779636304526477|4|1600043779|220|35.383490730525274|0|17|1433|-80.605588|9|35.43259|GRANOLA|0.0|1|NV PROTEIN GRANOLA OATS HONEY|13f1ef39385226d7fb218594ad6647929f83128a|2.8719573987198292|35.392509581117899|00016000437791|CEREAL|G1 GROCERY|-80.764523|80.764607981189812|202|1
35.06858|f5272fd0f25ec2668eadc6d467d8b106c17ce827|6.79|2015-01-06 19:15:00|1.4091206135396188|4|1200080994|273|0.612062184999033|0|47|55|-80.7007|8|35.06858|REGULAR|6.79|23|PEPSI FRIDGEMATE|1491831ee4d196c82983355845a5c9a99d794e89|1.1377023968546804|0.61242566243833529|00012000809941|CARBONATED BEVERAGES|BEVERAGE|-80.7007|1.4084929236641879|273|1
35.06858|14f8817799cf0235ed39b882dd820f5dca0a8b4d|6.49|2014-10-28 11:38:00|1.4091206135396188|4|1200080994|273|0.612062184999033|0|47|55|-80.7007|8|35.06858|REGULAR|6.49|23|PEPSI FRIDGEMATE|1491831ee4d196c82983355845a5c9a99d794e89|1.1377023968546804|0.61242566243833529|00012000809941|CARBONATED BEVERAGES|BEVERAGE|-80.7007|1.4084929236641879|273|1
35.06858|7dece82219d67af550e4797d73bff578f273b9d0|9.99|2014-09-16 19:45:00|1.4091206135396188|4|85877000246|273|0.612062184999033|0|47|458|-80.7007|82|35.06858|CRAFT BEER|0.0|16|OMB CHRISTMAS 12OZ 6PACK|1491831ee4d196c82983355845a5c9a99d794e89|1.1377023968546804|0.61242566243833529|00858770002461|DOMESTIC BEER|BEER|-80.7007|1.4084929236641879|273|1
35.06858|a590e01007e2570a9888ec76fd2cda37bdec24cb|13.99|2014-09-19 19:51:00|80.700712769248256|4|86787200002|273|35.0850451503984|0|42|458|-80.699909|82|35.002628|CRAFT BEER|0.0|16|THE UNKNOWN VEHOPCIRAPTOR 22OZ|1491831ee4d196c82983355845a5c9a99d794e89|1.1377023968546804|35.088667338853092|00867872000022|DOMESTIC BEER|BEER|-80.7007|80.700713764055649|477|1
35.06858|5332ace6beabe16be86385eed3022df03b9b24fd|3.58|2014-10-25 10:00:00|80.700712769248256|4|4850001775|273|35.085045141086376|0|42|338|-80.661096|56|35.172688|OTHER FRUIT JUICES|1.58|3|TROPICANA RASP LEMONADE 12 OZ|1491831ee4d196c82983355845a5c9a99d794e89|1.1377023968546804|35.088667338853092|00048500021545|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.7007|80.700725442152319|474|2
35.059823|cfdbe030802581fb1a3d6077810473919a0dc7d2|5.35|2014-12-04 15:06:00|80.816179662140996|2|3700041759|66|35.068745252339973|0|41|388|-80.771677|66|35.066546|NFS-DISHWASH PWDR/LIQUID|1.06|1|CASCADE PAC CITRUS BRZ 15CT|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00037000806288|DETERGENTS|G1 GROCERY|-80.816172|80.816174955839742|45|1
35.059823|481f55220f0ba5e39c264bf8db8e4c43605236b0|4.49|2014-12-26 14:40:00|80.816179662140996|2|4000031532|66|35.068745252587782|0|41|727|-80.770346|7|35.052812|SEASONAL CANDY-SINGLE FAC|2.25|1|I/O(C14)M&M PLAIN CHRISTMAS|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00040000315322|CANDY|G1 GROCERY|-80.816172|80.816173461718321|40|1
35.059823|8c54796945a035791c43643a1534520bae7e43ec|2.99|2014-10-23 16:21:00|80.816179662140996|2|4145811704|66|35.068745252504428|0|41|265|-80.8062|307|35.037115|FROZEN PIES|0.0|5|EDWARDS CHOC SUNDAE SINGLES|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00041458117049|DESSERTS FROZEN|FROZEN|-80.816172|80.816174087217505|27|1
35.059823|3172d7bc90997eaefac7568b659971209539790e|5.79|2014-10-30 17:07:00|80.816179662140996|2|4440015600|66|35.068745252504428|0|41|293|-80.8062|48|35.037115|FROZEN SEAFOOD|2.79|5|GORTON'S 18CT FISHSTICKS|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00044400156509|FROZEN MEALS|FROZEN|-80.816172|80.816174087217505|27|1
35.059823|0b80da770f9605ed8bcaba64d0618cb515ca81c9|2.99|2014-09-25 16:23:00|80.816179662140996|2|4145811704|66|35.068745252504428|0|41|265|-80.8062|307|35.037115|FROZEN PIES|0.0|5|EDWARDS CHOC SUNDAE SINGLES|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00041458117049|DESSERTS FROZEN|FROZEN|-80.816172|80.816174087217505|27|1
35.059823|5b022333e709df5ca39f4208307e1e1bc5e71a2c|2.99|2014-11-13 16:03:00|80.816179662140996|2|4145811704|66|35.068745252504428|0|41|265|-80.8062|307|35.037115|FROZEN PIES|0.49|5|EDWARDS CHOC SUNDAE SINGLES|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00041458117049|DESSERTS FROZEN|FROZEN|-80.816172|80.816174087217505|27|1
35.059823|622f444a9157095cd052fc272cb33a731af69b2c|4.69|2014-12-26 14:40:00|80.816179662140996|2|4900002468|66|35.068745252587782|0|41|54|-80.770346|8|35.052812|DIET|1.19|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816173461718321|40|1
35.059823|935f9e083d5cf85225e0e8fc13a3e1b990826cfa|4.99|2015-02-12 16:14:00|80.816179662140996|2|4900002468|66|35.068745252504428|0|41|54|-80.8062|8|35.037115|DIET|1.0|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|1
35.059823|e5b074bf54ff7f3f28defe12fdc5dde9a0460968|4.99|2015-03-07 16:34:00|80.816179662140996|2|4900002468|66|35.068745252504428|0|41|54|-80.8062|8|35.037115|DIET|2.49|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|1
35.059823|25c629b14caf361cad0b70cd1b29ec64815d7d31|4.99|2015-01-15 15:57:00|80.816179662140996|2|4900002468|66|35.068745252504428|0|41|54|-80.8062|8|35.037115|DIET|2.5|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|1
35.059823|3f632921037688c2788a75fefd64838d3bb49e8a|4.99|2015-02-05 17:20:00|80.816179662140996|2|4900002468|66|35.068745252504428|0|41|54|-80.8062|8|35.037115|DIET|0.0|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|1
35.059823|f923ca73fd50afa8c12bdc1a681b2f156e73db1a|4.99|2015-01-01 15:04:00|80.816179662140996|2|4900002468|66|35.068745252339973|0|41|54|-80.771677|8|35.066546|DIET|1.0|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174955839742|45|1
35.059823|41c5da2906840bd780a72ec471e02f29fc7c40d3|4.69|2014-09-18 15:59:00|80.816179662140996|2|4900002468|66|35.068745252504428|0|41|54|-80.8062|8|35.037115|DIET|1.19|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|1
35.059823|e93870e45b839ecd6725983f1b980a0abdd8066c|4.69|2014-10-16 16:42:00|1.4091206135396188|2|4900002468|66|0.6119093465164359|0|47|54|-80.816172|8|35.059823|DIET|0.0|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|0.61242566243833529|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|1.4105082902580508|66|1
35.059823|53fc38435cfb362610cf3f291abac4f0be19a3be|4.69|2014-09-11 15:37:00|80.816179662140996|2|4900002468|66|35.068745252504428|0|41|54|-80.8062|8|35.037115|DIET|2.35|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|1
35.059823|487a33d65619150a87eb2f4b923ff928298cef22|4.69|2014-10-09 15:35:00|80.816179662140996|2|4900002468|66|35.068745252587782|0|41|54|-80.770346|8|35.052812|DIET|1.19|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816173461718321|40|1
35.059823|f9928f5d9957385f9899ad529196811e03268cd9|4.99|2015-02-25 12:00:00|1.4091206135396188|2|4900002468|66|0.6119093465164359|0|47|54|-80.816172|8|35.059823|DIET|1.0|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|0.61242566243833529|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|1.4105082902580508|66|1
35.059823|e916dab4a93fe339a082e901a05e722bfbe6a0cf|4.99|2015-02-19 16:10:00|80.816179662140996|2|4900002468|66|35.068745252504428|0|41|54|-80.8062|8|35.037115|DIET|2.5|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|1
35.059823|a13af3a3c3f8761e2630277d87b0a148fbccb8e5|4.69|2014-11-06 15:29:00|80.816179662140996|2|4900002468|66|35.068745252504428|0|41|54|-80.8062|8|35.037115|DIET|2.35|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|1
35.059823|c9c44524b63a6a286394cedd2ac5370d044a9f77|4.69|2014-12-18 15:59:00|80.816179662140996|2|4900002468|66|35.068745252504428|0|41|54|-80.8062|8|35.037115|DIET|1.19|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|1
35.059823|dc407dc526d87fc4c3ff6552da79a8ddf340a261|4.99|2015-01-08 15:52:00|1.4091206135396188|2|4900002468|66|0.6119093465164359|0|47|54|-80.816172|8|35.059823|DIET|0.0|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|0.61242566243833529|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|1.4105082902580508|66|1
35.059823|ac81691df00af01395105016df2815bf34a0e03a|9.38|2014-11-28 15:49:00|80.816179662140996|2|4900002468|66|35.068745252504428|0|41|54|-80.8062|8|35.037115|DIET|5.44|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|2
35.059823|cade03f00e3c2c06d93f53a2d8424f795d8251cb|4.69|2014-10-02 15:31:00|80.816179662140996|2|4900002468|66|35.068745252504428|0|41|54|-80.8062|8|35.037115|DIET|2.35|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|1
35.059823|45596165a660d6a528890874089ecafba6a53e99|4.69|2014-12-12 14:56:00|80.816179662140996|2|4900002468|66|35.068745252504428|0|41|54|-80.8062|8|35.037115|DIET|0.0|23|DIET COKE .5 LITER/6 PK.|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.816172|80.816174087217505|27|1
35.059823|801fb635b52c42649dd83315ae304ceb692a20fe|1.25|2015-01-22 16:16:00|80.816179662140996|2|4850001775|66|35.068745252504428|0|41|335|-80.8062|56|35.037115|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA PP ORIGINAL 12 OZ|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00048500017753|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.816172|80.816174087217505|27|1
35.059823|8e827d9d2d3b01e39276895351e0f7d21701bf8d|1.79|2014-10-25 16:34:00|80.816179662140996|2|4850001775|66|35.068745252339973|0|41|335|-80.771677|56|35.066546|ORANGE JUICE-REGRIGERATED|0.79|3|TROPICANA PP ORIGINAL 12 OZ|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00048500017753|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.816172|80.816174955839742|45|1
35.059823|917df65f81e48d99efd5338719fdd1661aa44db2|3.49|2014-12-11 16:14:00|1.4091206135396188|2|7017715419|66|0.6119093465164359|0|47|233|-80.816172|37|35.059823|BLACK TEA|0.49|1|TWININGS DECAF EARL GREY|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|0.61242566243833529|00070177171674|TEA|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|866303475f5ca16c23095e253bc37def65f60809|4.23|2015-01-29 16:11:00|1.4091206135396188|2||66|0.6119093465164359|0|47|529|-80.816172|64|35.059823|FRESH ASPARAGUS|2.12|4|GREEN  ASPARAGUS|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|0.61242566243833529|00204080000008|FRESH PRODUCE|PRODUCE|-80.816172|1.4105082902580508|66|1
35.059823|021dbee4854f83c9251e5f4db005786edb9941bc|8.98|2014-10-03 14:52:00|80.816179662140996|2|4164120104|66|35.068745252504428|0|41|899|-80.8062|205|35.037115|KOSHER FROZEN FOODS|0.0|5|GOLDEN PANCAKE POTATO|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00041641201036|FROZEN KOSHER|FROZEN|-80.816172|80.816174087217505|27|2
35.059823|87682e44f8d4e136b1786dc181a835fb84f2593e|12.35|2014-09-21 11:31:00|80.816179662140996|2|20598600000|66|35.068745252603684|0|41|1800|-80.760919|400|35.024332|FFM BEEF|0.0|6|HT ROAST  BEEF|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00205986000000|FFM MEAT|DELI|-80.816172|80.816173308875435|343|1
35.059823|86e9e285566b0d3191f696aa30c739a544da526c|1.77|2014-10-05 16:03:00|80.816179662140996|2|7203614049|66|35.068745252465455|0|41|104|-80.848528|16|35.053394|APPLESAUCE-CUPS|0.5|1|HT APPLESAUCE 6PK UNSWTND|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00072036140494|FRUIT-CAN/JAR|G1 GROCERY|-80.816172|80.816174322633771|11|1
35.059823|1de4a13ddefc7b0b0d03141d0f41948ddfd5f80e|3.99|2014-10-18 14:09:00|80.816179662140996|2|4000015140|66|35.068745252339973|0|41|46|-80.771677|7|35.066546|PKG CHOC|0.49|1|3 MUSKETEER FUN SIZE|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00040000151227|CANDY|G1 GROCERY|-80.816172|80.816174955839742|45|1
35.059823|790e64096132535ebf41d5620c82a93c562d7ee9|9.99|2014-09-13 14:29:00|80.816179662140996|2|4200044517|66|35.068745252339973|0|41|426|-80.771677|72|35.066546|NFS-PAPER TOWELS|3.0|1|BRAWNY 6 BIG ROLL PICK A SIZE|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00042000445177|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.816172|80.816174955839742|45|1
35.059823|b3d125ffa7fba9e294c372063ba80325d57c1cb2|4.49|2014-11-20 16:03:00|80.816179662140996|2|8265700312|66|35.068745252504428|0|41|31|-80.8062|4|35.037115|NON CARBONATED WATER|0.5|1|DEER PARK SPRG WATER .5 LTR|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00082657003122|BOTTLED WATER|G1 GROCERY|-80.816172|80.816174087217505|27|1
35.059823|3ef0637ae68418909a6b437732fa44389c0dd508|4.99|2015-01-24 16:35:00|80.816179662140996|2|8265750406|66|35.068745252339973|0|41|31|-80.771677|4|35.066546|NON CARBONATED WATER|1.49|1|(U)DEER PARK WATER 24PK .5LT|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00082657504063|BOTTLED WATER|G1 GROCERY|-80.816172|80.816174955839742|45|1
35.059823|7aab3718533712bf9522bb616f528effed1449f6|4.99|2015-02-15 15:19:00|80.816179662140996|2|8265750406|66|35.068745252339973|0|41|31|-80.771677|4|35.066546|NON CARBONATED WATER|0.5|1|(U)DEER PARK WATER 24PK .5LT|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00082657504063|BOTTLED WATER|G1 GROCERY|-80.816172|80.816174955839742|45|1
35.059823|6e5658a3ce89334d76e17e4791b7dfbf29079a77|2.89|2015-02-16 14:02:00|1.4091206135396188|2|7203655029|66|0.6119093465164359|0|47|331|-80.816172|52|35.059823|NATURAL SLICED|1.22|3|HT RF PEPPER JACK SLICES|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|0.61242566243833529|00072036708694|CHEESE|DAIRY|-80.816172|1.4105082902580508|66|1
35.059823|549e7d818532d1e73b8ee1a6260ce500766289a7|2.19|2015-03-03 16:10:00|1.4091206135396188|2|2880000001|66|0.6119093465164359|0|47|247|-80.816172|39|35.059823|VEGETABLES-FLANKER|0.0|1|HANOVER THREE BEAN SALAD|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|0.61242566243833529|00028800000013|VEGETABLES-CAN/JAR|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|e4402817c3ea7d62227503bf6120713ad3e30106|3.99|2014-12-24 16:21:00|80.816179662140996|2|88810911004|66|35.068745252339973|0|41|1046|-80.771677|173|35.066546|CAKES|2.0|7|HOSTESS CINN COFFEE CAKE|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00888109110048|SWEET BAKED GOODS|COMMERCIAL BAKERY|-80.816172|80.816174955839742|45|1
35.059823|dfdcd5a7d0f5fe83b0f037f0a9c0929f17e80636|4.99|2015-01-15 15:57:00|80.816179662140996|2|7099210227|66|35.068745252504428|0|41|6785|-80.8062|1568|35.037115|MAGAZINES WEEKLY|0.0|18|10227 PEOPLE|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00070992102273|MAGAZINES|GM|-80.816172|80.816174087217505|27|1
35.059823|d84c45cad2c021a1b19f3b50000d6cf3236ecff0|3.99|2015-02-12 16:11:00|80.816179662140996|2|4000042065|66|35.068745252504428|0|41|46|-80.8062|7|35.037115|PKG CHOC|1.99|1|I/O MM MILK CHOCOLATE BONUS|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00040000420651|CANDY|G1 GROCERY|-80.816172|80.816174087217505|27|1
35.059823|3042258cb06d2b5032a313ef80db5d508a48ba36|1.79|2014-10-21 14:47:00|80.816179662140996|2|2500000024|66|35.068745252504428|0|41|335|-80.8062|56|35.037115|ORANGE JUICE-REGRIGERATED|0.0|3|SIMPLY ORANGE JUICE PULP FREE|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00025000000249|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.816172|80.816174087217505|27|1
35.059823|701cf16ae1e93fe88a5be525e26ef64c4e7bdac3|2.79|2015-02-25 12:02:00|1.4091206135396188|2|1130038110|66|0.6119093465164359|0|47|50|-80.816172|7|35.059823|PEG CANDY|0.0|1|BRACHS LEMON DROPS|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|0.61242566243833529|00011300384011|CANDY|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|7a5c1ae07f860411440819cd56b746420c75038f|2.79|2014-12-18 15:55:00|80.816179662140996|2|1130038110|66|35.068745252504428|0|41|50|-80.8062|7|35.037115|PEG CANDY|0.0|1|BRACHS LEMON DROPS|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00011300384011|CANDY|G1 GROCERY|-80.816172|80.816174087217505|27|1
35.059823|6da4ebebc76635a0baea9d47d5f2d9b407ff4bf1|2.79|2015-01-29 16:09:00|1.4091206135396188|2|1130038110|66|0.6119093465164359|0|47|50|-80.816172|7|35.059823|PEG CANDY|0.0|1|BRACHS LEMON DROPS|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|0.61242566243833529|00011300384011|CANDY|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|92b638c2b775418722cce4a0016b197b1c2340a9|2.79|2015-01-01 15:05:00|80.816179662140996|2|1130038110|66|35.068745252339973|0|41|50|-80.771677|7|35.066546|PEG CANDY|0.0|1|BRACHS LEMON DROPS|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00011300384011|CANDY|G1 GROCERY|-80.816172|80.816174955839742|45|1
35.059823|059e1ac4ee3a32925e546231762fca8ec19e6d16|2.79|2015-01-08 15:53:00|1.4091206135396188|2|1130038110|66|0.6119093465164359|0|47|50|-80.816172|7|35.059823|PEG CANDY|0.0|1|BRACHS LEMON DROPS|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|0.61242566243833529|00011300384011|CANDY|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|c85cdd0907d392574d365d1afab49d2f808624a2|2.79|2015-02-19 16:07:00|80.816179662140996|2|1130038110|66|35.068745252504428|0|41|50|-80.8062|7|35.037115|PEG CANDY|0.0|1|BRACHS LEMON DROPS|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00011300384011|CANDY|G1 GROCERY|-80.816172|80.816174087217505|27|1
35.059823|63025eaccedfdebca98d440d3802169a8d06cf5c|2.79|2015-03-07 16:29:00|80.816179662140996|2|1130038110|66|35.068745252504428|0|41|50|-80.8062|7|35.037115|PEG CANDY|0.0|1|BRACHS LEMON DROPS|211d1fa65abd67186b4f552be4497cc972dc61b8|0.6165061128897139|35.070508771677183|00011300384011|CANDY|G1 GROCERY|-80.816172|80.816174087217505|27|1
35.372142|f8c7a3cf653837a9e684d216e67683eaec98d27f|11.58|2014-09-17 18:46:00|1.4102725052409182|3|5833618000|122|0.617360341382972|0|1|254|-80.782849|892|35.372142|PREMIUM PIZZA|1.79|5|RISTORANTE MOZZARELLA PIZZA|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|0.61833652052202714|00058336180002|FROZEN PIZZA|FROZEN|-80.782849|1.4099266941914086|122|2
35.372142|b7d6fdf3df68139d81e9b580a9484254a22a75f7|6.3|2014-09-27 22:29:00|1.4102725052409182|3|7265500105|122|0.617360341382972|0|1|1278|-80.782849|48|35.372142|SINGLE SERVE NUTRITIONAL|2.3|5|HC CAFE STEAMERS CHK MARGARITA|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|0.61833652052202714|00072655001053|FROZEN MEALS|FROZEN|-80.782849|1.4099266941914086|122|2
35.372142|7fc52af9824b75ab640982644b6b37b9f1c423d6|3.79|2015-02-27 13:24:00|1.4102725052409182|3|3700034885|122|0.617360341382972|0|1|425|-80.782849|72|35.372142|NFS-PAPER NAPKINS|0.0|1|BOUNTY QUILTED NAPKINS 200CT|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|0.61833652052202714|00037000348856|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|d8ddcab280fb96fd40d2bbe888ec1db09e725795|5.97|2014-12-03 19:20:00|1.4102725052409182|3|81483201043|122|0.617360341382972|0|1|4207|-80.782849|1200|35.372142|COUGH DROP-ADULT|2.9699999999999998|17|LUDENS S/F WILD CHERRY BAG|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|0.61833652052202714|00814832010539|COUGH/COLD/SINUS|HBC|-80.782849|1.4099266941914086|122|3
35.372142|69c3032ecc15d0da3baf795a1eced70cc9b6e9d9|4.79|2014-12-31 19:28:00|1.4102725052409182|3|18685200031|122|0.617360341382972|0|1|275|-80.782849|45|35.372142|SUPER PREMIUM ICE CREAM|0.8|5|TALENTI CARIBB COCONUT GELATO|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|0.61833652052202714|00186852000327|ICE CREAM|FROZEN|-80.782849|1.4099266941914086|122|1
35.372142|f2c8f1725b28f4dd48b3289edf8d027f69cfd35d|8.17|2014-10-20 19:14:00|1.4102725052409182|3|20895700000|122|0.617360341382972|0|1|977|-80.782849|201|35.372142|FRESH HT CHICKEN|2.85|2|HT VALUE PK CHCKN LEG QUARTERS|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|0.61833652052202714|00208957000009|POULTRY|MEAT|-80.782849|1.4099266941914086|122|1
35.372142|ceb01845bda510804d64d632675c052028c0c2a9|4.59|2014-09-30 13:26:00|80.779636304526477|3|7535303362|122|35.376092266991911|0|17|6253|-80.709466|1550|35.124987|TAPES/DUCT TAPE|0.0|18|DUCK TAPE 1.88X15 YD NEON PINK|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|35.392509581117899|00075353033623|HARDWARE|GM|-80.782849|80.78285984128712|157|1
35.372142|f0fcf6c9e592419f2b83fa266e7312553c840944|3.99|2015-02-02 18:34:00|1.4102725052409182|3|7218069274|122|0.617360341382972|0|1|1277|-80.782849|279|35.372142|FROZEN SNACKS|0.99|5|PAGODA CRM CHEESE WONTONS|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|0.61833652052202714|00072180698568|FROZEN SANDWICH AND SNACKS|FROZEN|-80.782849|1.4099266941914086|122|1
35.372142|025ec6d673344734967a5e3ed3cc4f8148504174|3.99|2014-10-24 10:24:00|1.4102725052409182|3|89299200227|122|0.617360341382972|0|1|4237|-80.782849|1200|35.372142|MEDICATED LIP CARE|1.49|17|(FE) OS HNYSUCKLE HNYDEW  BALM|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|0.61833652052202714|00892992002298|COUGH/COLD/SINUS|HBC|-80.782849|1.4099266941914086|122|1
35.372142|3d1cf2b479bc623742709585228e4f0f7e2510ac|3.99|2014-10-31 18:30:00|1.4102725052409182|3|81793900034|122|0.617360341382972|0|1|722|-80.782849|73|35.372142|NFS-HAND SOAPS|2.02|1|METHOD HAND SOAP BOTAN GARDEN|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|0.61833652052202714|00817939011942|PERSONAL SOAP/BATH ADDITIVES|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|3aa7af96673a5f1908d821e606d11df31949b35e|12.97|2014-11-21 15:12:00|1.4102725052409182|3|7203697650|122|0.617360341382972|0|1|8433|-80.782849|1769|35.372142|ALKALINE AA|5.98|18|HT AA BATTERIES 24PK|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|0.61833652052202714|00072036976505|BATTERY & FLASHLIGHT|GM|-80.782849|1.4099266941914086|122|1
35.372142|dabdc88e97fe33ecfe291b489dfbe4b051d76e9b|28.24|2014-10-27 18:23:00|1.4102725052409182|3|20137100000|122|0.617360341382972|0|1|296|-80.782849|49|35.372142|RANCHER BEEF|5.19|2|VALUE PK T-BONE STEAKS|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|0.61833652052202714|00201371000006|BEEF|MEAT|-80.782849|1.4099266941914086|122|1
35.372142|33972375588e26156c005f6e9ecbbd208fecca9c|1.69|2014-10-28 13:17:00|80.779636304526477|3|4900000044|122|35.376092266991911|0|17|54|-80.709466|8|35.124987|DIET|0.0|23|CB COKE ZERO 20 OZ|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|35.392509581117899|00049000040869|CARBONATED BEVERAGES|BEVERAGE|-80.782849|80.78285984128712|157|1
35.372142|36d9119edfbc27667b3785b75ef5982c71cf957e|2.45|2014-11-26 15:09:00|1.4102725052409182|3|7203663217|122|0.617360341382972|0|1|330|-80.782849|55|35.372142|EGGS|0.0|3|HT GRADE A LARGE EGGS 18 CT|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|0.61833652052202714|00072036632173|EGGS FRESH|DAIRY|-80.782849|1.4099266941914086|122|1
35.372142|db2796e614f9a96f3dacc900f7ded23a9335c3b8|4.9|2014-09-26 16:57:00|80.779636304526477|3|7203663217|122|35.376092276777776|0|17|330|-80.764523|55|35.341927|EGGS|0.9|3|HT GRADE A LARGE EGGS 18 CT|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|35.392509581117899|00072036632173|EGGS FRESH|DAIRY|-80.782849|80.782850117093091|220|2
35.372142|ba7d44ab355e29a7747ae16fd66e63b77861b357|3.99|2014-10-04 14:50:00|1.4102725052409182|3|2500005542|122|0.617360341382972|0|1|335|-80.782849|56|35.372142|ORANGE JUICE-REGRIGERATED|0.99|3|SIMPLY ORANGE WITH MANGO|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|0.61833652052202714|00025000054372|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.782849|1.4099266941914086|122|1
35.372142|99c91b71a836dc5249a571511b502dff115b2be2|3.99|2015-01-15 18:50:00|1.4102725052409182|3|7247000221|122|0.617360341382972|0|1|1641|-80.782849|377|35.372142|PACKAGED DONUTS|0.0|14|K K 6 FUDGE ICED W/CREME    PP|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|0.61833652052202714|00072470002211|DONUTS|BAKERY|-80.782849|1.4099266941914086|122|1
35.372142|ec3e37676f4b51a35b79d42b972028d923c47228|4.55|2014-09-24 19:32:00|1.4102725052409182|3|7457000400|122|0.617360341382972|0|1|275|-80.782849|45|35.372142|SUPER PREMIUM ICE CREAM|1.21|5|H DAZS PINEAPPLE COCONUT|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|0.61833652052202714|00074570610075|ICE CREAM|FROZEN|-80.782849|1.4099266941914086|122|1
35.372142|34a95d1a51bc76f7d80f282a109dafa435ccbeaf|3.95|2014-09-19 21:08:00|1.4102725052409182|3|7457000400|122|0.617360341382972|0|1|275|-80.782849|45|35.372142|SUPER PREMIUM ICE CREAM|0.0|5|H DAZS PINEAPPLE COCONUT|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|0.61833652052202714|00074570610075|ICE CREAM|FROZEN|-80.782849|1.4099266941914086|122|1
35.372142|340d06464b1f83edfce3d8252252fab3045f1679|3.95|2014-09-15 18:52:00|1.4102725052409182|3|7457000400|122|0.617360341382972|0|1|275|-80.782849|45|35.372142|SUPER PREMIUM ICE CREAM|0.0|5|H DAZS PINEAPPLE COCONUT|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|0.61833652052202714|00074570610075|ICE CREAM|FROZEN|-80.782849|1.4099266941914086|122|1
35.372142|f0c3f4cf82577cdc8d376fa9c003dc8032ff9727|1.59|2014-12-17 18:47:00|1.4102725052409182|3|7203638020|122|0.617360341382972|0|1|226|-80.782849|35|35.372142|SUGAR-POWDERED|0.0|1|HT CONFECTIONERS SUGAR|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|0.61833652052202714|00072036380302|SUGAR/SUBSTITUTES|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|40ee555e5700df61ccf9ed5798010a01b5772f31|13.99|2014-10-29 12:27:00|80.779636304526477|3|3680007390|122|35.376092266991911|0|17|4234|-80.709466|1200|35.124987|PSE SOLID DOSE|4.2|17|(PP) PSE TC LORATADINE D-24|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|35.392509581117899|00036800073906|COUGH/COLD/SINUS|HBC|-80.782849|80.78285984128712|157|1
35.372142|4c25ff7371d07c6d19bde79eeb07035bb2ec643f|1.29|2014-10-18 15:32:00|80.779636304526477|3|2200000899|122|35.376092276058856|0|17|48|-80.746334|7|35.41832|REGISTER GUM|0.0|1|EXTRA SPEARMINT|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|35.392509581117899|00022000008992|CANDY|G1 GROCERY|-80.782849|80.782852129019801|190|1
35.372142|93fafbb1688b8e94796c6a7d9b05633ed40786df|2.49|2014-10-02 19:59:00|1.4102725052409182|3|3760401465|122|0.617360341382972|0|1|6821|-80.782849|1580|35.372142|J HOOK LAMI PROGRAM|0.0|18|FLEX STRAW 150CT-NEON|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|0.61833652052202714|00037604014652|J-HOOK|GM|-80.782849|1.4099266941914086|122|1
35.372142|34039ed9d78397bcf679e6016bcc8530fb39da2c|9.58|2014-09-22 19:25:00|1.4102725052409182|3|18685200031|122|0.617360341382972|0|1|275|-80.782849|45|35.372142|SUPER PREMIUM ICE CREAM|0.0|5|TALENTI CRML APPLE PIE GELATO|233c51d7f3a2b452a5e63422f55277987103f4a1|0.27295459302329644|0.61833652052202714|00186852000860|ICE CREAM|FROZEN|-80.782849|1.4099266941914086|122|2
35.17739|de0f5ae969045454dbbd54dc6979394f2043c772|1.59|2014-09-12 15:35:00|80.801203185414451|4|78616201000|208|35.193014467442438|0|24|31|-80.826724|4|35.195689|NON CARBONATED WATER|0.59|1|VIT WATER XXX 20 OZ|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00786162150004|BOTTLED WATER|G1 GROCERY|-80.80146|80.801461451627773|412|1
35.17739|15d9ed403b6f92de296693c17ace445e0574d3d0|1.49|2015-03-03 15:20:00|80.801203185414451|4|7618316363|208|35.193014467442438|0|24|99|-80.826724|32|35.195689|LIQUID TEA|0.49|1|SNAPPLE KIWI STRAWBERRY|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00076183163634|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.80146|80.801461451627773|412|1
35.17739|ef1e2c66b553f1ed538f664fa60ea232edbd12e2|2.98|2015-03-05 23:04:00|1.4094857484078087|4|7618316363|208|0.613961277758128|0|26|99|-80.80146|32|35.17739|LIQUID TEA|0.98|1|SNAPPLE KIWI STRAWBERRY|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|0.61471665291522548|00076183163634|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.80146|1.4102515174184975|208|2
35.17739|9c9949f8f80907b0874652a43c6d5bc74cfcce85|2.5|2014-10-05 18:56:00|80.801203185414451|4|78142100610|208|35.193014467442438|0|24|1601|-80.826724|371|35.195689|BRANDED BREAD|0.51|14|LA BREA WHEAT BAGUETTE|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00781421521182|BREAD|BAKERY|-80.80146|80.801461451627773|412|1
35.17739|6071c14972f0123448780ac08cedb80822a41718|3.49|2015-03-02 20:40:00|80.801203185414451|4|4850002115|208|35.193014467442438|0|24|338|-80.826724|56|35.195689|OTHER FRUIT JUICES|0.99|3|DOLE BLENDS-ORANGE PEACH MANGO|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00048500021125|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.80146|80.801461451627773|412|1
35.17739|f15a7e42fd27a45696df2eedb757033f43a0f223|8.58|2015-01-09 11:38:00|80.801203185414451|4|2840015636|208|35.193014467442438|0|24|204|-80.826724|31|35.195689|TORTILLA CHIPS|2.15|1|DORTIOS NACHO CHEESE|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00028400156363|SNACKS|G1 GROCERY|-80.80146|80.801461451627773|412|2
35.17739|7a0e6f51005a4bae65f600bb76751eac0bd0dd36|10.15|2014-12-29 11:14:00|1.4094857484078087|4|20895700000|208|0.613961277758128|0|26|977|-80.80146|201|35.17739|FRESH HT CHICKEN|3.54|2|HT VALUE PK CHCKN LEG QUARTERS|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|0.61471665291522548|00208957000009|POULTRY|MEAT|-80.80146|1.4102515174184975|208|1
35.17739|0266ba2a85cac531c77dcb757fb2f316adbc254f|2.68|2014-10-14 15:25:00|80.801203185414451|4|7203698078|208|35.193014467442438|0|24|242|-80.826724|39|35.195689|CANNED BEANS|0.68|1|HT BEANS KIDNEY LIGHT RED|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00072036411150|VEGETABLES-CAN/JAR|G1 GROCERY|-80.80146|80.801461451627773|412|4
35.17739|c4d9b80547b74e5d8834086007d799f35dc1d8a1|1.34|2014-10-02 10:31:00|80.801203185414451|4|7047045916|208|35.193014467442438|0|24|685|-80.826724|61|35.195689|GREEK|0.0|3|YOPLAIT GREEK BLEND STWBRY RAS|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00070470459158|YOGURT|DAIRY|-80.80146|80.801461451627773|412|1
35.17739|0eb12c5586c6a9c9c0c8642010d72c5831d03576|2.5|2014-10-07 15:12:00|80.801203185414451|4|7203695204|208|35.193014467442438|0|24|1603|-80.826724|371|35.195689|PRIVATE LABEL BREAD|0.51|14|BAND OF BAKERS BAGUETTE|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00072036952042|BREAD|BAKERY|-80.80146|80.801461451627773|412|1
35.17739|4048bcbd79e3eac27a984a47c60769c573e3d9f5|2.99|2014-12-11 15:16:00|80.801203185414451|4|7203698526|208|35.193014467442438|0|24|201|-80.826724|31|35.195689|POTATO CHIPS|0.49|1|HT TRADER KETTLE CHIP RED FAT|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00072036985262|SNACKS|G1 GROCERY|-80.80146|80.801461451627773|412|1
35.17739|ab72b387f2c9dd769bff8213a91f4f8ebe662f0a|2.47|2014-09-12 12:03:00|80.801203185414451|4||208|35.193014467442438|0|24|501|-80.826724|64|35.195689|FRESH PEARS|0.37|4|BARTLETT PEARS|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00204409000009|FRESH PRODUCE|PRODUCE|-80.80146|80.801461451627773|412|1
35.17739|b5c49e6731e168df1b32ebd3a8b1f5cd7e99d8df|1.0|2015-02-22 22:17:00|1.4094857484078087|4||208|0.613961277758128|0|26|512|-80.80146|64|35.17739|FRSH PROD FRSH FRUIT REM|0.0|4|MANGOS|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|0.61471665291522548|00204959000009|FRESH PRODUCE|PRODUCE|-80.80146|1.4102515174184975|208|1
35.17739|29b1e664d4e385f126f2e0b3f628957b9f0d5054|1.0|2015-02-01 20:05:00|1.4094857484078087|4||208|0.613961277758128|0|26|512|-80.80146|64|35.17739|FRSH PROD FRSH FRUIT REM|0.0|4|MANGOS|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|0.61471665291522548|00204959000009|FRESH PRODUCE|PRODUCE|-80.80146|1.4102515174184975|208|1
35.17739|34357680eb660569792d6aaa848eb66dfa12fd94|1.79|2014-10-10 13:59:00|80.801203185414451|4|7342000006|208|35.193014467442438|0|24|322|-80.826724|53|35.195689|SOUR CREAM|0.59|3|DAISY SOUR CREAM|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00073420000066|CULTURES|DAIRY|-80.80146|80.801461451627773|412|1
35.17739|cd96c522e358795f5a7a22b6a593848e41ce87b3|2.89|2014-10-26 20:53:00|1.4094857484078087|4|7618364374|208|0.613961277758128|0|26|99|-80.80146|32|35.17739|LIQUID TEA|0.9|1|SNAPPLE HALF & HALF|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|0.61471665291522548|00076183001035|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|36bf6e7c2dd00406071ff00f9e298ddfdac8b9c9|2.69|2014-11-13 10:31:00|80.801203185414451|4|3663202720|208|35.193014467442438|0|24|688|-80.826724|61|35.195689|LIGHT|0.0|3|DANNON FRUIT ON BOTTOM PEACH|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00036632018267|YOGURT|DAIRY|-80.80146|80.801461451627773|412|1
35.17739|6b86b098a4e4bc8a1e25ff7742aa97fe627af372|3.59|2014-10-03 14:01:00|80.801203185414451|4|7433610102|208|35.193014467442438|0|24|342|-80.826724|57|35.195689|FRESH MILK|0.0|3|HIGHLAND CREST WHOLE MILK|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00074336879203|MILK|DAIRY|-80.80146|80.801461451627773|412|1
35.17739|8bd103a2d38a80e11015ac17e1cdf117148c4ae4|2.99|2015-01-26 15:26:00|1.4094857484078087|4|7433610102|208|0.613961277758128|0|26|342|-80.80146|57|35.17739|FRESH MILK|0.0|3|HIGHLAND CREST WHOLE MILK|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|0.61471665291522548|00074336879203|MILK|DAIRY|-80.80146|1.4102515174184975|208|1
35.17739|dea553131e71cd42f9082e8a1d3ab295d64a0793|4.29|2015-02-02 16:22:00|1.4094857484078087|4|2840016014|208|0.613961277758128|0|26|201|-80.80146|31|35.17739|POTATO CHIPS|1.79|1|LAYS CLASSIC|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|0.61471665291522548|00028400160148|SNACKS|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|bc1fc9b380a8c55454d36f618771e7c1c8589944|2.99|2015-01-15 11:14:00|80.801203185414451|4|3120020007|208|35.193014467442438|0|24|130|-80.826724|20|35.195689|CRANBERRY JUICE/DRINKS-SHELF|0.0|1|OSPRAY CRANBERRY JUICE|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00031200200075|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.80146|80.801461451627773|412|1
35.17739|17c0a548d4a8e13d3d202d6e44c84e2fa87a63d5|1.67|2015-02-04 16:07:00|80.801203185414451|4|7203614011|208|35.193014467442438|0|24|110|-80.826724|16|35.195689|FRUIT-CORE|0.33|1|HT PEACHES HALVES HS 15|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00072036140104|FRUIT-CAN/JAR|G1 GROCERY|-80.80146|80.801461451627773|412|1
35.17739|3e38270de98aac1200bc49a3c43eb4c24248ed6e|1.17|2014-11-14 11:48:00|80.801203185414451|4|7203628044|208|35.193014467442438|0|24|161|-80.826724|25|35.195689|PEPPERS|0.0|1|HT JALAPENO SLICES|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00072036280442|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.80146|80.801461451627773|412|1
35.17739|389076976c6833bb68d593389477fc2dd05ed94c|2.99|2014-10-17 14:12:00|80.801203185414451|4|20443000000|208|35.193014467442438|0|24|510|-80.826724|64|35.195689|FRESH PINEAPPLE|0.0|4|GOLD PINEAPPLES|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00643126072003|FRESH PRODUCE|PRODUCE|-80.80146|80.801461451627773|412|1
35.17739|f6f565802265b52a1bb4652779310c72c6c184f2|5.35|2014-12-16 11:47:00|80.801203185414451|4|7203697668|208|35.193014467442438|0|24|317|-80.826724|52|35.195689|CHUNK AND BAR CHEESE|2.35|3|HT MOZZARELLA CHEESE|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00072036980472|CHEESE|DAIRY|-80.80146|80.801461451627773|412|1
35.17739|c5bbba4143d5d909b8d0f072a1ecba3a58c25e36|0.37|2014-12-22 18:53:00|1.4094857484078087|4|7203659035|208|0.613961277758128|0|26|688|-80.80146|61|35.17739|LIGHT|0.0|3|HT NONFAT PEACH YOGURT|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|0.61471665291522548|00072036570413|YOGURT|DAIRY|-80.80146|1.4102515174184975|208|1
35.17739|111bc9085b3fef9d1390555a7b6f27ff2ed97aed|0.74|2015-01-08 15:52:00|80.801203185414451|4|7203659035|208|35.193014467442438|0|24|688|-80.826724|61|35.195689|LIGHT|0.07|3|HT NONFAT PEACH YOGURT|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00072036570413|YOGURT|DAIRY|-80.80146|80.801461451627773|412|2
35.17739|b2b63463e4a0c505577341a7af8220e1b89da233|1.77|2015-02-26 22:13:00|1.4094857484078087|4|7203657031|208|0.613961277758128|0|26|322|-80.80146|53|35.17739|SOUR CREAM|0.0|3|HT SOUR CREAM|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|0.61471665291522548|00072036570314|CULTURES|DAIRY|-80.80146|1.4102515174184975|208|1
35.17739|d3251d9c36615a8ab97e1c57da0388efb8734da6|2.67|2014-09-21 20:08:00|1.4094857484078087|4|7047045916|208|0.613961277758128|0|26|685|-80.80146|61|35.17739|GREEK|0.67|3|YOPLAIT GREEK BLEND BLUEBERRY|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|0.61471665291522548|00070470459165|YOGURT|DAIRY|-80.80146|1.4102515174184975|208|2
35.17739|fead43e444382b4405e3748537f48c73c1e84657|2.29|2014-10-30 10:25:00|80.801203185414451|4|7203695175|208|35.193014467442438|0|24|1607|-80.826724|371|35.195689|FROZEN DOUGH (BREAD)|0.0|14|FRESH LRG FRENCH BREAD|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00072036951755|BREAD|BAKERY|-80.80146|80.801461451627773|412|1
35.17739|8e5c98a036dd0c434886d4f72a70633491e821cb|1.5|2015-02-19 15:12:00|80.801203185414451|4||208|35.193014467442438|0|24|1617|-80.826724|373|35.195689|ROLLS BULK|0.0|14|BULK ROLLS|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00072036955555|ROLLS|BAKERY|-80.80146|80.801461451627773|412|2
35.17739|5e88984f116dda6c1667ebb51594951a69cb2386|1.5|2015-03-05 15:14:00|80.801203185414451|4||208|35.193014467442438|0|24|1635|-80.826724|375|35.195689|BULK (BAGELS)|0.0|14|BULK  BAGELS|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00072036955500|BAGELS|BAKERY|-80.80146|80.801461451627773|412|2
35.17739|74599b03c4b0ce7b5871c7f1543a7709b8d67906|1.99|2015-02-28 16:07:00|80.801203185414451|4|7203695644|208|35.193014467442438|0|24|1647|-80.826724|379|35.195689|PACKAGED MUFFINS|0.0|14|2CT RAISIN BRAN MUFFINS|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00072036956446|MUFFINS|BAKERY|-80.80146|80.801461451627773|412|1
35.17739|08cdbb2d82d5e40d2924093ac33d17b99bcc3c86|1.29|2014-10-16 10:22:00|80.801203185414451|4|1657191030|208|35.193014467442438|0|24|30|-80.826724|4|35.195689|CARBONATED WATER|0.29|1|SPARKLING ICE PEACH NECTARINE|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00016571940348|BOTTLED WATER|G1 GROCERY|-80.80146|80.801461451627773|412|1
35.17739|326f1dd6b5b03ccc089de0c4058cc548308faa6d|1.29|2015-02-13 11:20:00|80.801203185414451|4|1657191030|208|35.193014467442438|0|24|30|-80.826724|4|35.195689|CARBONATED WATER|0.29|1|SPARKLING ICE PEACH NECTARINE|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00016571940348|BOTTLED WATER|G1 GROCERY|-80.80146|80.801461451627773|412|1
35.17739|472ec5bd4da4ff36eaeedcfe4743ca5293060afe|1.29|2015-02-24 15:29:00|80.801203185414451|4|1657191030|208|35.193014467442438|0|24|30|-80.826724|4|35.195689|CARBONATED WATER|0.29|1|SPARKLING ICE PEACH NECTARINE|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00016571940348|BOTTLED WATER|G1 GROCERY|-80.80146|80.801461451627773|412|1
35.17739|e8c0956609f99ecfa1a233098613166328b776c7|1.29|2014-11-22 15:44:00|80.801203185414451|4|1657191030|208|35.193014467442438|0|24|30|-80.826724|4|35.195689|CARBONATED WATER|0.29|1|SPARKLING ICE PEACH NECTARINE|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00016571940348|BOTTLED WATER|G1 GROCERY|-80.80146|80.801461451627773|412|1
35.17739|6e8b252dc5b78aa1a163881a710a3aad20136e03|2.58|2014-09-30 11:19:00|80.801203185414451|4|1657191030|208|35.193014467442438|0|24|30|-80.826724|4|35.195689|CARBONATED WATER|0.58|1|SPARKLING ICE PEACH NECTARINE|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00016571940348|BOTTLED WATER|G1 GROCERY|-80.80146|80.801461451627773|412|2
35.17739|67cb48e57cbfbf4f9d72b409106b5635d986b19a|0.74|2014-09-28 17:52:00|80.801203185414451|4|7203659035|208|35.193014467442438|0|24|688|-80.826724|61|35.195689|LIGHT|0.0|3|HT NONFAT PLAIN YOGURT|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00072036040299|YOGURT|DAIRY|-80.80146|80.801461451627773|412|2
35.17739|128e19ac2a58e885b1440220bf3956e917e250c1|4.99|2015-01-09 11:37:00|80.801203185414451|4|1111018700|208|35.193014467442438|0|24|1647|-80.826724|379|35.195689|PACKAGED MUFFINS|2.5|14|FFM 4 CT LEMON POPPY MUFFIN|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00011110187048|MUFFINS|BAKERY|-80.80146|80.801461451627773|412|1
35.17739|28420ec3dde5e810e810937221d949612028466f|2.59|2014-11-02 18:24:00|80.801203185414451|4|2100061223|208|35.193014467442438|0|24|316|-80.826724|52|35.195689|CREAM CHEESE|0.0|3|PHILLY CREAM CHEESE - BRICK|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00021000612239|CHEESE|DAIRY|-80.80146|80.801461451627773|412|1
35.17739|2877208d6f11c926ae106876419d56ab08aa70ff|1.33|2014-11-04 11:50:00|80.801203185414451|4||208|35.193014467442438|0|24|500|-80.826724|64|35.195689|FRESH APPLES|0.67|4|GOLD DEL APPLE, WA 72|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00204020000006|FRESH PRODUCE|PRODUCE|-80.80146|80.801461451627773|412|1
35.17739|5373f35402ec6b6cd04ad3e768172d751fc95f77|4.69|2015-03-02 20:39:00|80.801203185414451|4|7756712130|208|35.193014467442438|0|24|251|-80.826724|43|35.195689|NON-DAIRY NOVELTIES|0.0|5|POPSICLE RAINBOW|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00077567021533|FROZEN NOVELTIES|FROZEN|-80.80146|80.801461451627773|412|1
35.17739|d2cb707b8f8d1170be1c4daffc8c6dbd17693e2c|3.49|2014-12-05 14:55:00|80.801203185414451|4|664|208|35.193014467442438|0|24|1639|-80.826724|377|35.195689|BULK (DONUTS)|0.0|14|PICK 6  DONUTS|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00000000006640|DONUTS|BAKERY|-80.80146|80.801461451627773|412|1
35.17739|6ce655e50234cea792ecb298c20378f85834487b|3.49|2014-11-19 16:27:00|80.801203185414451|4|664|208|35.193014467442438|0|24|1639|-80.826724|377|35.195689|BULK (DONUTS)|0.0|14|PICK 6  DONUTS|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00000000006640|DONUTS|BAKERY|-80.80146|80.801461451627773|412|1
35.17739|99e4ee7752e3ac52990969deb61b5cbc4c9c1dd9|3.49|2014-09-18 17:05:00|80.801203185414451|4|664|208|35.193014467442438|0|24|1639|-80.826724|377|35.195689|BULK (DONUTS)|0.0|14|PICK 6  DONUTS|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00000000006640|DONUTS|BAKERY|-80.80146|80.801461451627773|412|1
35.17739|b8f5af8a3532466818051e0f9aad525513c781b5|3.49|2015-02-13 11:19:00|80.801203185414451|4|664|208|35.193014467442438|0|24|1639|-80.826724|377|35.195689|BULK (DONUTS)|0.0|14|PICK 6  DONUTS|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00000000006640|DONUTS|BAKERY|-80.80146|80.801461451627773|412|1
35.17739|1783fa2dbac2242b5db6aed4cb375f5dbd246264|3.49|2015-01-18 16:55:00|80.801203185414451|4|664|208|35.193014467442438|0|24|1639|-80.826724|377|35.195689|BULK (DONUTS)|0.0|14|PICK 6  DONUTS|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00000000006640|DONUTS|BAKERY|-80.80146|80.801461451627773|412|1
35.17739|9899c367154fbb3da4ded7c5fa993854a98db4f8|1.39|2014-10-03 14:00:00|80.801203185414451|4|7618316356|208|35.193014467442438|0|24|99|-80.826724|32|35.195689|LIQUID TEA|0.39|1|SNAPPLE PEACH TEA 16 OZ|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00076183163566|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.80146|80.801461451627773|412|1
35.17739|310a9c9cbe3df8a2c1449aa4f2507964b4e8fc1c|6.23|2014-09-12 12:04:00|80.801203185414451|4||208|35.193014467442438|0|24|500|-80.826724|64|35.195689|FRESH APPLES|0.0|4|GRANNY SMITH APPLES 72|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00204017000002|FRESH PRODUCE|PRODUCE|-80.80146|80.801461451627773|412|1
35.17739|990df473239838b1f3e2756b757b9f1b1514393b|4.27|2014-10-23 10:25:00|80.801203185414451|4||208|35.193014467442438|0|24|565|-80.826724|64|35.195689|REDUCED PRODUCE|0.0|4|PRODUCE REWRAP BY LB|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00204844000008|FRESH PRODUCE|PRODUCE|-80.80146|80.801461451627773|412|3
35.17739|75e9c714935e90c8bee3bb3000b099647e4678f2|2.75|2014-09-26 10:25:00|80.801203185414451|4||208|35.193014467442438|0|24|565|-80.826724|64|35.195689|REDUCED PRODUCE|0.0|4|PRODUCE REWRAP BY CT|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00204845000007|FRESH PRODUCE|PRODUCE|-80.80146|80.801461451627773|412|2
35.17739|7715f6e2cd4c6b3b66ec83bba53546abfe194129|2.0|2014-09-18 10:25:00|80.801203185414451|4|812|208|35.193014467442438|0|24|1639|-80.826724|377|35.195689|BULK (DONUTS)|0.0|14|NEW BULK DONUT CODE|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00000000008120|DONUTS|BAKERY|-80.80146|80.801461451627773|412|2
35.17739|5fc23bc7a041dfb898ffe876c85a076446db1bd7|4.0|2014-10-21 12:00:00|80.801203185414451|4|812|208|35.193014467442438|0|24|1639|-80.826724|377|35.195689|BULK (DONUTS)|0.0|14|NEW BULK DONUT CODE|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00000000008120|DONUTS|BAKERY|-80.80146|80.801461451627773|412|4
35.17739|5271663a5a0582305a144dd8893ca8b6943f4092|4.0|2014-09-11 10:28:00|80.801203185414451|4|812|208|35.193014467442438|0|24|1639|-80.826724|377|35.195689|BULK (DONUTS)|0.0|14|NEW BULK DONUT CODE|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00000000008120|DONUTS|BAKERY|-80.80146|80.801461451627773|412|4
35.17739|5f8f44b20a8be1f7147b6578b9b29f88f21684e1|15.88|2015-01-09 11:36:00|80.801203185414451|4|27085500000|208|35.193014467442438|0|24|973|-80.826724|201|35.195689|FRESH PERDUE CHICKEN|0.0|2|PERDUE OVEN STUFFER ROASTER|244c651d0c08ee39c810d3fccc38a04cad5b986a|1.079612971647154|35.194272495053255|00270855000009|POULTRY|MEAT|-80.80146|80.801461451627773|412|1
35.43259|52c1b134147faeb19d23d5e1c933a3fe3f8ed9af|13.99|2015-02-02 14:27:00|1.4057311447477159|4|7203695696|202|0.6184153580092175|0|52|1653|-80.605588|381|35.43259|CELEBRATION CAKES|0.0|14|1/8 SHEET DL MBL W/WHT BUTCRM|27423e3f281a66e2a181650a903e91a474a10224|0.8357089404423385|0.6209993146566879|00072036956965|CAKES|BAKERY|-80.605588|1.406832906106031|202|1
35.43259|5a8488134dca104fe9da95df479e67c0fe84781a|6.79|2014-11-30 18:39:00|1.4057311447477159|4|7800001180|202|0.6184153580092175|0|52|55|-80.605588|8|35.43259|REGULAR|1.4|23|CHEERWINE 12PK CANS|27423e3f281a66e2a181650a903e91a474a10224|0.8357089404423385|0.6209993146566879|00070925000102|CARBONATED BEVERAGES|BEVERAGE|-80.605588|1.406832906106031|202|1
35.43259|88206386295759ec6c23d10e6d6ec984a0309a34|5.99|2014-12-30 17:04:00|80.607132136635443|4|3746605490|202|35.444684614858581|0|9|727|-80.746334|7|35.41832|SEASONAL CANDY-SINGLE FAC|3.0|1|I/O(C14)LINDOR HOLIDAY MC BAG|27423e3f281a66e2a181650a903e91a474a10224|0.8357089404423385|35.47365851958088|00037466054902|CANDY|G1 GROCERY|-80.605588|80.605599735963409|190|1
35.43259|03886c6af2c5a9c3aa93009199ace22cbd5c9e02|8.99|2014-11-23 17:38:00|80.607132136635443|4|87126011085|202|35.444684594172351|0|9|740|-80.737839|87|35.297134|NFS-ROSE BQT|0.0|9|BUNCH- 10 CONSUMER ROSE|27423e3f281a66e2a181650a903e91a474a10224|0.8357089404423385|35.47365851958088|00871260110859|FLORAL|FLORAL|-80.605588|80.605617858894675|258|1
35.43259|911672b212c305c4bb904b39b0dbd9b2ab7aed80|5.0|2014-09-28 09:14:00|1.4057311447477159|4|2400016286|202|0.6184153580092175|0|52|245|-80.605588|39|35.43259|VEGETABLES-CORE|0.0|1|DEL MONTE GRN BEANS CUT|27423e3f281a66e2a181650a903e91a474a10224|0.8357089404423385|0.6209993146566879|00024000162865|VEGETABLES-CAN/JAR|G1 GROCERY|-80.605588|1.406832906106031|202|4
35.43259|c45c1d456a85f435a3a8b20559a2f1b61b485174|3.75|2015-02-18 19:57:00|1.4057311447477159|4|5250005005|202|0.6184153580092175|0|52|182|-80.605588|28|35.43259|MAYO|0.0|1|DUKES MAYONNAISE 32|27423e3f281a66e2a181650a903e91a474a10224|0.8357089404423385|0.6209993146566879|00052500050054|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.605588|1.406832906106031|202|1
35.43259|6fc5236cf2f94dded31367f550d04c28f05c28cf|9.99|2014-10-02 21:17:00|80.607132136635443|4|8500001667|202|35.444684598067283|0|9|9945|-80.66939|885|35.28326|NFS POP OTHER WHITE|0.0|13|CB-BAREFOOT MOSCATO 1.5L|27423e3f281a66e2a181650a903e91a474a10224|0.8357089404423385|35.47365851958088|00085000016671|POPULAR (4-$7.99)|WINE|-80.605588|80.605615379184812|46|1
35.43259|e1b61ae8286ab2fd555e063d8fcd55162170a22f|6.57|2015-01-18 12:18:00|1.4057311447477159|4|2400001830|202|0.6184153580092175|0|52|245|-80.605588|39|35.43259|VEGETABLES-CORE|0.0|1|DEL MONTE GRN BEANS CUT 28.|27423e3f281a66e2a181650a903e91a474a10224|0.8357089404423385|0.6209993146566879|00024000018308|VEGETABLES-CAN/JAR|G1 GROCERY|-80.605588|1.406832906106031|202|3
35.43259|72bf338a3b1fb4f6165680d68d39cf7fd8959988|4.99|2015-02-04 20:58:00|1.4057311447477159|4|1111018700|202|0.6184153580092175|0|52|1647|-80.605588|379|35.43259|PACKAGED MUFFINS|2.49|14|FFM 4 CT BLUEBERRY MUFFIN|27423e3f281a66e2a181650a903e91a474a10224|0.8357089404423385|0.6209993146566879|00011110187000|MUFFINS|BAKERY|-80.605588|1.406832906106031|202|1
35.43259|615022c8ebd409fd6f3cf485b9c5497d03c884a1|4.49|2014-11-27 13:18:00|1.4057311447477159|4|5210000263|202|0.6184153580092175|0|52|1245|-80.605588|34|35.43259|SINGLE SPICES|1.35|1|MC POULTRY SEASONING|27423e3f281a66e2a181650a903e91a474a10224|0.8357089404423385|0.6209993146566879|00052100002637|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.605588|1.406832906106031|202|1
35.43259|9201b88f48edc4af4bee00c4f34a89104f1d968f|14.99|2014-11-21 20:32:00|1.4057311447477159|4|3410057256|202|0.6184153580092175|0|52|455|-80.605588|82|35.43259|DOMESTIC PREMIUM 12PK&>|0.0|16|MILLER LITE 18PK 12OZ BTL|27423e3f281a66e2a181650a903e91a474a10224|0.8357089404423385|0.6209993146566879|00034100572563|DOMESTIC BEER|BEER|-80.605588|1.406832906106031|202|1
35.03469|76cbb4cc80c083bef8a5b8284e97adf8b1bba096|37.1|2014-11-01 10:55:00|1.4132775322775095|4|7203608135|82|0.6114706929155321|0|58|82|-80.97058|11|35.03469|VINEGAR|0.0|1|HT VINEGAR WHITE DISTILLED 128|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|0.61177642288969325|00072036081353|CONDIMENTS|G1 GROCERY|-80.97058|1.4132032182494703|82|14
35.03469|e3f8534c096824f277ad81911e42bdfd76211036|3.39|2015-01-17 09:47:00|80.970593795509558|4|7203646021|82|35.066747962327092|0|4|1463|-80.994596|42|35.061685|REGULAR FROZEN FRUIT|0.0|5|HT BERRY MEDLEY|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|35.073829668338668|00072036460622|FROZEN FRUIT|FROZEN|-80.97058|80.970586762569255|475|1
35.03469|56f71cd0b7986ebfd14ce3bef92f60664bd5d7b7|1.39|2014-10-27 19:47:00|1.4132775322775095|4|7203624015|82|0.6114706929155321|0|58|149|-80.97058|23|35.03469|WHSE PASTA CORE|0.42|1|HT PASTA SPAGHETTI 16|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|0.61177642288969325|00072036240156|PASTA|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|3b531c8d1d0a2a28857a2cdcf6e6da0fcf99d464|4.33|2015-02-01 13:15:00|80.970593795509558|4|20358700000|82|35.066747962327092|0|4|656|-80.994596|137|35.061685|STR MDE VALUE ADDED PORK|2.17|2|CAJUN & RICE STUFFED PORK CHOP|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|35.073829668338668|00203587000009|PORK|MEAT|-80.97058|80.970586762569255|475|1
35.03469|77585b3d39f195e0ef737ec0f980e449aaa595c8|3.05|2015-01-27 13:11:00|80.970593795509558|4|20165700000|82|35.066747953909534|0|4|297|-80.848528|49|35.053394|GROUND BEEF|0.34|2|HT GROUND BEEF CHUCK 80% LEAN|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|35.073829668338668|00201657000003|BEEF|MEAT|-80.97058|80.970609172601343|11|1
35.03469|0271191c1d2c109d9bae84de8a120e2edc911df5|3.73|2014-12-30 12:34:00|80.970593795509558|4|20165700000|82|35.066747953909534|0|4|297|-80.848528|49|35.053394|GROUND BEEF|0.83|2|HT GROUND BEEF CHUCK 80% LEAN|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|35.073829668338668|00201657000003|BEEF|MEAT|-80.97058|80.970609172601343|11|1
35.03469|bf9af20ca64d6c2d28ecec47c0121c2b5e4f1ec7|1.99|2014-09-17 17:43:00|80.970593795509558|4|3599530782|82|35.066747951169035|0|4|6412|-81.027334|1556|34.977331|CARS/TRUCKS/MOTORCYCLES|0.0|18|MATCHBOX BASIC CARS|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|35.073829668338668|00035995307827|TOYS|GM|-80.97058|80.970613365006798|149|1
35.03469|1501191fcfb185c62f09af5ca07b0bf1303e8c77|4.99|2014-11-24 18:49:00|1.4132775322775095|4|3800031834|82|0.6114706929155321|0|58|74|-80.97058|9|35.03469|RTE CEREAL ALL FAMILY|0.0|1|KELL MINI WHEATS BITE LG BOX|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|0.61177642288969325|00038000318344|CEREAL|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|ee5bfd8f853c899365bdbd224d83d33e9c04da6d|2.5|2014-12-23 18:08:00|80.970593795509558|4|78142100610|82|35.066747962327092|0|4|1601|-80.994596|371|35.061685|BRANDED BREAD|0.0|14|LA BREA WHEAT BAGUETTE|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|35.073829668338668|00781421521182|BREAD|BAKERY|-80.97058|80.970586762569255|475|1
35.03469|4e16e1b903deb891a94a365958645fb9a80cf1a9|19.98|2014-12-13 17:52:00|1.4132775322775095|4|7203695262|82|0.6114706929155321|0|58|1671|-80.97058|383|35.03469|CHEESE CAKE|0.0|14|HAZELNUT CHEESECAKE|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|0.61177642288969325|00072036953285|PASTRY CASE|BAKERY|-80.97058|1.4132032182494703|82|2
35.03469|268d2b66812b2763dc77aa907b7a6f15f880c93c|13.99|2014-12-31 12:25:00|80.970593795509558|4|7203688033|82|35.066747953909534|0|4|563|-80.848528|64|35.053394|FRESH VEGETABLE/FRUIT TRAYS|1.0|4|HT VEGETABLE TRAY, LARGE|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|35.073829668338668|00072036880338|FRESH PRODUCE|PRODUCE|-80.97058|80.970609172601343|11|1
35.03469|3ba76f5fc3deb04f3e25a457da3288a0fc16cdfc|8.85|2015-01-12 18:59:00|80.970593795509558|4|2370001409|82|35.066747962327092|0|4|291|-80.994596|48|35.061685|FROZEN POUTLRY|0.0|5|TYSON SOUTHERN CKN TENDERLOINS|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|35.073829668338668|00023700014856|FROZEN MEALS|FROZEN|-80.97058|80.970586762569255|475|1
35.03469|b241f9f917534766adc1c3228ce4c7703b3ff5d2|3.79|2015-01-16 07:45:00|80.970593795509558|4|7774529186|82|35.066747953909534|0|4|555|-80.848528|64|35.053394|PACKAGED SALADS|0.0|4|R.P. BISTRO SANTA FE SALAD|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|35.073829668338668|00077745291888|FRESH PRODUCE|PRODUCE|-80.97058|80.970609172601343|11|1
35.03469|a6c815c15446bb8162326080fa2b2c40e94ebe96|30.729999999999997|2015-01-07 20:06:00|1.4132775322775095|4|7120228515|82|0.6114706929155321|0|58|1463|-80.97058|42|35.03469|REGULAR FROZEN FRUIT|0.0|5|DOLE PINEAPPLE CHUNKS|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|0.61177642288969325|00071202285151|FROZEN FRUIT|FROZEN|-80.97058|1.4132032182494703|82|7
35.03469|09a9b8b6c7b92c2ba28054c5a0fb5e84084b414b|3.98|2015-02-02 12:47:00|80.970593795509558|4|7127923100|82|35.066747953909534|0|4|555|-80.848528|64|35.053394|PACKAGED SALADS|0.0|4|F.E. BABY SPRING SALAD MIX|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|35.073829668338668|00071279231006|FRESH PRODUCE|PRODUCE|-80.97058|80.970609172601343|11|2
35.03469|b5d7110adc68646ca23c663c25dfa2de3a8e168a|3.54|2014-12-23 18:07:00|80.970593795509558|4|7203698067|82|35.066747962327092|0|4|365|-80.994596|56|35.061685|REFRIGERATED TEAS|0.0|3|HARRIS TEETER SWEET TEA|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|35.073829668338668|00072036980670|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.97058|80.970586762569255|475|2
35.03469|02174f7049e5bdd34d70996b5b78b48a9c906427|6.49|2015-02-14 09:23:00|80.970593795509558|4|8139200005|82|35.066747962327092|0|4|9983|-80.994596|889|35.061685|NFS-SPARKLING|0.0|13|J. ROGET SPUMANTE|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|35.073829668338668|00081392000052|SPARKLING|WINE|-80.97058|80.970586762569255|475|1
35.03469|ca9bc7b71fd643abf7f8de0cdad11572cedc021d|0.94|2014-11-12 18:12:00|1.4132775322775095|4|7248600220|82|0.6114706929155321|0|58|11|-80.97058|2|35.03469|MUFFIN MIXES|0.0|1|JIFFY CORN MUFFIN MIX|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|0.61177642288969325|00072486002205|BAKING MIXES|G1 GROCERY|-80.97058|1.4132032182494703|82|2
35.03469|fcf2f5303a9b5e6c91d738aa3168eee22fdcf6fe|3.79|2014-11-29 11:18:00|80.970593795509558|4|2500005542|82|35.066747962327092|0|4|335|-80.994596|56|35.061685|ORANGE JUICE-REGRIGERATED|0.79|3|SIMPLY ORANGE ORIGINAL|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|35.073829668338668|00025000055423|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.97058|80.970586762569255|475|1
35.03469|a00a09a95f5d4a68e95726c7c31d3c62832e4eb9|3.29|2015-03-08 19:20:00|1.4132775322775095|4|5250005002|82|0.6114706929155321|0|58|182|-80.97058|28|35.03469|MAYO|0.0|1|DUKES MAYONNAISE 16|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|0.61177642288969325|00052500050023|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|6628ee287615d7f712f29bed5eeb15599352a41d|2.99|2014-09-10 18:07:00|1.4132775322775095|4|2880010314|82|0.6114706929155321|0|58|245|-80.97058|39|35.03469|VEGETABLES-CORE|0.0|1|HANOVER GREEN BEAN CUT 50|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|0.61177642288969325|00028800103141|VEGETABLES-CAN/JAR|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|d61ee2185604c6c5c0095414e6e2a09e3925a2a7|8.99|2014-12-31 17:17:00|1.4132775322775095|4|61278110230|82|0.6114706929155321|0|58|265|-80.97058|307|35.03469|FROZEN PIES|0.0|5|M CALLENDER LEM MERINGUE PIE|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|0.61177642288969325|00612781102301|DESSERTS FROZEN|FROZEN|-80.97058|1.4132032182494703|82|1
35.03469|8864be3b336f93f569432b93220e27c0361ff8b0|3.79|2014-12-19 07:55:00|80.970593795509558|4|1254631053|82|35.066747953909534|0|4|48|-80.848528|7|35.053394|REGISTER GUM|0.79|1|DENTYNE ICE SPEARMINT BTL|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|35.073829668338668|00012546310796|CANDY|G1 GROCERY|-80.97058|80.970609172601343|11|1
35.03469|5f52a153aab2e1e54b8286a8a66783b06dda8949|13.99|2014-11-17 17:08:00|1.4132775322775095|4|75452700201|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|NEW BELGIUM FOLLY VARIETY 12PK|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|0.61177642288969325|00754527002015|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|df65ad45ae64f0499fbbaeefe4754e82ec796964|4.59|2014-10-27 17:30:00|1.4132775322775095|4|7581002425|82|0.6114706929155321|0|58|79|-80.97058|273|35.03469|ASIAN SAUCES/SEASONINGS|0.6|1|SAN J ORG TAMARI LITE 50% LSD|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|0.61177642288969325|00075810024256|ASIAN PREP. FOODS|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|713b7ba71e96c07e55ebe44eae7aa9c016c34ff6|3.79|2014-12-19 12:35:00|80.970593795509558|4|7774529186|82|35.066747953909534|0|4|555|-80.848528|64|35.053394|PACKAGED SALADS|0.0|4|R.P. BISTRO MEDITERRANEAN|2e3a421afda9e30afcb803cd65fb1305f8126c1e|2.2151278126251195|35.073829668338668|00077745294988|FRESH PRODUCE|PRODUCE|-80.97058|80.970609172601343|11|1
34.95459|fdf6f226b3f220a40072132c39e66dc473addfa3|1.99|2014-12-03 18:12:00|1.4091206135396188|3|3900004504|182|0.6100726841846847|0|47|114|-80.758228|14|34.95459|PUMPKIN|0.0|1|LIBBY SOLID PACK PUMPKIN|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00039000045049|DESSERTS/GELS/SYRUPS|G1 GROCERY|-80.758228|1.4094969766762753|182|1
34.95459|30e46cab0deef2417f30ec6b8532e958496b6273|3.89|2014-09-23 16:44:00|1.4091206135396188|3|3800039125|182|0.6100726841846847|0|47|74|-80.758228|9|34.95459|RTE CEREAL ALL FAMILY|0.9|1|KELLOGG RICE KRISPIES 9|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00038000318443|CEREAL|G1 GROCERY|-80.758228|1.4094969766762753|182|1
34.95459|19b263eeb6fcfdfcf8bc8d56b09ce4f8df7a9968|2.69|2015-02-24 08:37:00|1.4091206135396188|3|4119640471|182|0.6100726841846847|0|47|1201|-80.758228|33|34.95459|RTS CANNED|0.69|1|PROG LIGHT BEEF POT ROAST|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00041196404814|SOUP|G1 GROCERY|-80.758228|1.4094969766762753|182|1
34.95459|b76b0fb635387ebddd5738e7cd172fa1452d759c|10.99|2014-10-25 14:33:00|1.4091206135396188|3|4740000126|182|0.6100726841846847|0|47|3917|-80.758228|1075|34.95459|DISPOSABLE RAZOE-MEN|3.0|17|(FE) GIL FUSION DISPOSBL RZR|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00047400001268|SHAVING NEEDS/MEN HAIR|HBC|-80.758228|1.4094969766762753|182|1
34.95459|379b830faac506b33a696bd2dbacc7f7e9a387a6|3.09|2015-01-07 18:46:00|1.4091206135396188|3|7225001854|182|0.6100726841846847|0|47|1034|-80.758228|163|34.95459|HOT DOG|0.0|7|NATOWN 8PK BUTTER HOTS|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00072250018548|BUNS/ROLLS|COMMERCIAL BAKERY|-80.758228|1.4094969766762753|182|1
34.95459|ced20af6a1a160e304f239fc735b87b579400e6d|1.37|2015-03-09 17:31:00|1.4091206135396188|3|7203690021|182|0.6100726841846847|0|47|1033|-80.758228|163|34.95459|HAMBURGER|0.0|7|H T HAMBURGER BUNS|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00072036900210|BUNS/ROLLS|COMMERCIAL BAKERY|-80.758228|1.4094969766762753|182|1
34.95459|6251fe3aef34fb09c9e799f8ab83f7d3c6223010|3.49|2014-12-17 15:34:00|1.4091206135396188|3|4069503007|182|0.6100726841846847|0|47|555|-80.758228|64|34.95459|PACKAGED SALADS|0.0|4|ROMIANE HEARTS|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00033383651620|FRESH PRODUCE|PRODUCE|-80.758228|1.4094969766762753|182|1
34.95459|e1bbd94324f305cf1a84687c1c7c30cc9b8a2974|5.49|2015-01-20 12:24:00|1.4091206135396188|3|2301290132|182|0.6100726841846847|0|47|1477|-80.758228|485|34.95459|SUSHI HYBRID|0.0|6|SPICY CALIFORNIA ROLL SP|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00023012901325|SUSHI|DELI|-80.758228|1.4094969766762753|182|1
34.95459|abb38d027ad743977e31b941d3abd47ad7d1c3bf|3.09|2015-02-15 13:59:00|1.4091206135396188|3|7225002313|182|0.6100726841846847|0|47|1033|-80.758228|163|34.95459|HAMBURGER|0.0|7|NATOWN 8PK BUTTER HAMS|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00072250023139|BUNS/ROLLS|COMMERCIAL BAKERY|-80.758228|1.4094969766762753|182|1
34.95459|87e08cb9ed0fca04fcb8e9dfc1a32eed450f4b2f|6.58|2014-10-01 17:54:00|1.4091206135396188|3|7225091171|182|0.6100726841846847|0|47|1033|-80.758228|163|34.95459|HAMBURGER|0.0|7|NATOWN WHITEWHEAT HAMS|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00072250911719|BUNS/ROLLS|COMMERCIAL BAKERY|-80.758228|1.4094969766762753|182|2
34.95459|07c6471d54a6336ce89e77db87a0191300b1644a|2.69|2015-03-05 18:44:00|1.4091206135396188|3|7225001739|182|0.6100726841846847|0|47|1025|-80.758228|162|34.95459|WHITE|0.0|7|NATOWN WHITEWHEAT RTOP BRD|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00072250017398|SLICED BREAD|COMMERCIAL BAKERY|-80.758228|1.4094969766762753|182|1
34.95459|f1bdb9414d61aff7dad57c0ab3869ff1c7779a5e|3.55|2014-11-08 19:54:00|1.4091206135396188|3|7433610102|182|0.6100726841846847|0|47|342|-80.758228|57|34.95459|FRESH MILK|0.0|3|HIGHLAND CREST 2% REDUCE FAT|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00074336101021|MILK|DAIRY|-80.758228|1.4094969766762753|182|1
34.95459|03ddc57ff2991a3ed24e08be82cef7fe374782d5|6.98|2014-12-24 12:41:00|1.4091206135396188|3|7203688136|182|0.6100726841846847|0|47|556|-80.758228|64|34.95459|PACKAGED VEGETABLES|1.0|4|HT CELERY & CARROTS AQUA PACK|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00072036881267|FRESH PRODUCE|PRODUCE|-80.758228|1.4094969766762753|182|2
34.95459|6bd090fb488a238fedf0c8d63c8dd8bd55244d6f|8.59|2014-12-22 20:15:00|1.4091206135396188|3|7050105370|182|0.6100726841846847|0|47|3237|-80.758228|1020|34.95459|ACNE PRODUCTS|1.72|17|(E)NEUT PINK GRPFRT ACNE SCRUB|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00070501053607|FACIAL CLEANSER & MOISTURIZER|HBC|-80.758228|1.4094969766762753|182|1
34.95459|186a25fbd3cc9977924070944e606b56c43f615c|1.69|2014-12-18 07:29:00|1.4091206135396188|3|1200000129|182|0.6100726841846847|0|47|55|-80.758228|8|34.95459|REGULAR|0.0|23|CB DR PEPPER 20 OZ NR SINGLE|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00078000082401|CARBONATED BEVERAGES|BEVERAGE|-80.758228|1.4094969766762753|182|1
34.95459|da52666f707e8f35a1a9d78ba8b9c4e8aa7a4e82|5.99|2014-11-20 06:44:00|1.4091206135396188|3|88552321821|182|0.6100726841846847|0|47|1403|-80.758228|389|34.95459|THAW AND SELL PIES|1.0|14|"8"" NO SGR ADD PUMPKIN PIE"|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00885523218213|PIES|BAKERY|-80.758228|1.4094969766762753|182|1
34.95459|64d99b0882767a41599b48f5a2f50f4221c0b28f|2.99|2014-11-14 16:03:00|1.4091206135396188|3|3800035900|182|0.6100726841846847|0|47|41|-80.758228|6|34.95459|BREAKFAST BARS|0.0|1|KLGS NUTRI GRN BAR APPLE CINN|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00038000356001|BREAKFAST FOODS|G1 GROCERY|-80.758228|1.4094969766762753|182|1
34.95459|735ecc4d018322c802295e3882d87876c7cc0628|35.99|2014-11-15 11:05:00|1.4091206135396188|3|20496600000|182|0.6100726841846847|0|47|1153|-80.758228|87|34.95459|NFS-FRESH CUT ARRANGE|0.0|9|*MIXED VASE ARRANGEMENTS|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00204966000009|FLORAL|FLORAL|-80.758228|1.4094969766762753|182|1
34.95459|79a9c3d32200ac1db92d1caeb930de860cbb831c|6.58|2014-11-24 16:04:00|1.4091206135396188|3|1600048037|182|0.6100726841846847|0|47|1251|-80.758228|12|34.95459|WHOLESOME COOKIES|0.0|1|FIBER ONE DBL CHOCOLATE COOKIE|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00016000480360|COOKIES|G1 GROCERY|-80.758228|1.4094969766762753|182|2
34.95459|53ba2a6f8e86ad00f71080151ebf700d3e882471|2.99|2015-02-08 21:04:00|1.4091206135396188|3|7007700107|182|0.6100726841846847|0|47|1279|-80.758228|48|34.95459|SINGLE SERVE FLAVOR|0.0|5|TAI-PEI CHICKEN FRIED RICE|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00070077001071|FROZEN MEALS|FROZEN|-80.758228|1.4094969766762753|182|1
34.95459|dcce7d12389ac032a09b5dea796be31373a39fab|19.99|2015-01-28 19:45:00|1.4091206135396188|3|1780013476|182|0.6100726841846847|0|47|156|-80.758228|24|34.95459|NFS-DOG FOOD-DRY|5.0|1|PURINA BENEFUL|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00017800134767|PET FOOD/SUPPLIES|G1 GROCERY|-80.758228|1.4094969766762753|182|1
34.95459|735e8333b29ed312d895b7e1237b330d28f7a4c9|10.99|2014-12-09 15:50:00|1.4091206135396188|3|2270012705|182|0.6100726841846847|0|47|3016|-80.758228|1000|34.95459|BRAND-COVER GIRL|0.0|17|CG LASHBLST FUSION MASC VRY BL|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00022700127047|COSMETICS|HBC|-80.758228|1.4094969766762753|182|1
34.95459|831b40dc7c0013c8a14eb27d2d52bbace4bc7ebd|10.99|2014-12-15 07:28:00|1.4091206135396188|3|2270012705|182|0.6100726841846847|0|47|3016|-80.758228|1000|34.95459|BRAND-COVER GIRL|0.0|17|CG LASHBLST FUSION MASC VRY BL|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00022700127047|COSMETICS|HBC|-80.758228|1.4094969766762753|182|1
34.95459|40f55d71813ab98f05d0cfd9512f338558fa620c|7.58|2014-11-15 16:13:00|1.4091206135396188|3|7774529186|182|0.6100726841846847|0|47|555|-80.758228|64|34.95459|PACKAGED SALADS|0.0|4|R.P. BISTRO BOWL COBB SALAD|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|0.61242566243833529|00077745291871|FRESH PRODUCE|PRODUCE|-80.758228|1.4094969766762753|182|2
34.95459|ac8e81d460b91d314d0fa5091a28c39493fa5af8|9.78|2015-02-21 22:21:00|80.762257539052428|3|7027223204|182|34.963046623339338|0|54|323|-80.699686|57|35.000049|TOPPINGS-REFRIGERATED|2.78|3|REDDI WIP EXTRA CREAMY|305be44309dab5499df1d365a54a6890c2b880ff|0.5843324101533035|34.983028186791387|00070272232089|MILK|DAIRY|-80.758228|80.758235622007263|249|2
35.23102|46f6b92e4a2e13e5e94f5354648eff393922cf24|2.49|2015-01-13 14:33:00|80.843945456961976|4|7203688048|205|35.234004274107683|0|59|526|-80.86175|64|35.40953|FRESH MUSHROOMS|0.0|4|HT SLICED BABY BELLAS|31798de1550bad9377eb2bf16d74f3b8febd773f|0.20620645804475607|35.232478750868765|00072036880482|FRESH PRODUCE|PRODUCE|-80.8438|80.843806476331721|209|1
35.23102|9053168fa36d373a58c68c4a1edf4cc9e0fa613e|3.99|2015-01-20 14:28:00|80.843945456961976|4|6055600161|205|35.234004274107683|0|59|556|-80.86175|64|35.40953|PACKAGED VEGETABLES|0.0|4|CUTBUTTERNUT SQUASH|31798de1550bad9377eb2bf16d74f3b8febd773f|0.20620645804475607|35.232478750868765|00640344020601|FRESH PRODUCE|PRODUCE|-80.8438|80.843806476331721|209|1
35.23102|23722be28817e1639bf0cdc3460ee223226777d3|1.89|2015-02-10 17:35:00|80.843945456961976|4|7680828008|205|35.234004274107683|0|59|149|-80.86175|23|35.40953|WHSE PASTA CORE|0.39|1|BARILLA PASTA ANGEL HAIR|31798de1550bad9377eb2bf16d74f3b8febd773f|0.20620645804475607|35.232478750868765|00076808501063|PASTA|G1 GROCERY|-80.8438|80.843806476331721|209|1
35.006282|01ed6dcf04325ad70cc2328b2132176a768d270b|11.98|2014-10-02 10:24:00|1.4091206135396188|4|7203695440|60|0.6109748797816256|0|47|1403|-80.562829|389|35.006282|THAW AND SELL PIES|3.0|14|"8"" SWEET POTATO PIE"|31ce379859a777e8d5ba1575058993b831f22977|0.4669838150754594|0.61242566243833529|00072036959362|PIES|BAKERY|-80.562829|1.4060866207711706|60|2
35.006282|f5b610104aaa79529b8d314a0242e3f59cc4b472|1.79|2014-10-26 13:45:00|1.4091206135396188|4|7142901230|60|0.6109748797816256|0|47|238|-80.562829|38|35.006282|RICE FLAVORED|0.79|1|ZATARAINS RICE SPANISH.|31ce379859a777e8d5ba1575058993b831f22977|0.4669838150754594|0.61242566243833529|00071429012271|RICE GRAINS AND BEANS|G1 GROCERY|-80.562829|1.4060866207711706|60|1
35.006282|2caac52816cb81b86dbe19993760bcf1b3b1a7d0|2.29|2014-10-03 11:14:00|1.4091206135396188|4|7203633079|60|0.6109748797816256|0|47|1244|-80.562829|21|35.006282|OTHER NUTS|0.29|1|HT DRY ROAST SUNFLOWER KERNEL|31ce379859a777e8d5ba1575058993b831f22977|0.4669838150754594|0.61242566243833529|00072036330796|NUTS|G1 GROCERY|-80.562829|1.4060866207711706|60|1
35.28326|d84c8787517f35a90c6ad2a8585dae7f45cef229|8.0|2015-01-29 19:06:00|1.4094857484078087|3||46|0.6158090578372145|0|26|511|-80.66939|64|35.28326|FRESH AVOCADOS|0.75|4|AVOCADOS, HASS XL 36CT|36462aa2eaa3d07ae740dc36bdebe3cbf48f3072|1.2330772300493043|0.61471665291522548|00204770000004|FRESH PRODUCE|PRODUCE|-80.66939|1.4079464610753885|46|4
35.28326|07e830b7a724e0b0515b8e35ac185cc6d7e4ed51|2.19|2015-01-27 21:29:00|1.4094857484078087|3|64420941200|46|0.6158090578372145|0|26|10|-80.66939|2|35.28326|LAYER CAKE MIX|0.0|1|D HINES SPICE CAKE MIX|36462aa2eaa3d07ae740dc36bdebe3cbf48f3072|1.2330772300493043|0.61471665291522548|00644209410606|BAKING MIXES|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|1d9f3ed4644b20ff8696d29794a16924aaa55406|10.58|2015-02-01 17:56:00|80.669414401537693|3|20895300000|46|35.301105445815907|0|19|977|-80.764523|201|35.341927|FRESH HT CHICKEN|0.0|2|HT FRESH BNLS CHICKEN BREAST|36462aa2eaa3d07ae740dc36bdebe3cbf48f3072|1.2330772300493043|35.305725790410776|00208953000003|POULTRY|MEAT|-80.66939|80.66939387625591|220|1
35.28326|b5ac16f75604c2a8980fe8481cc83e2c720f7c78|4.99|2015-02-13 09:07:00|1.4094857484078087|3|1117132944|46|0.6158090578372145|0|26|5606|-80.66939|1512|35.28326|BRUSH-KITCHEN|0.0|18|DAWN KITCHEN BRUSH|36462aa2eaa3d07ae740dc36bdebe3cbf48f3072|1.2330772300493043|0.61471665291522548|00011171329449|BROOMS/MOPS & BRUSHES|GM|-80.66939|1.4079464610753885|46|1
35.28326|a403cdbd8a8327b2d4e5ac5ec444abd290eb98b2|3.25|2014-11-14 12:32:00|1.4094857484078087|3|7203656080|46|0.6158090578372145|0|26|318|-80.66939|52|35.28326|SHREDDED/GRATED CHEESE|3.25|3|HT SHREDDED MOZZ/PROVLONE|36462aa2eaa3d07ae740dc36bdebe3cbf48f3072|1.2330772300493043|0.61471665291522548|00072036705174|CHEESE|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|a10d761cea2f1c4691c173f98b6481a7de6f0673|6.59|2015-01-08 20:06:00|1.4094857484078087|3|7940035291|46|0.6158090578372145|0|26|3814|-80.66939|1070|35.28326|INVISIBLE-FEMALE|0.0|17|DOVE WMN CARE NURISH AP/DEO|36462aa2eaa3d07ae740dc36bdebe3cbf48f3072|1.2330772300493043|0.61471665291522548|00079400352910|DEODORANT|HBC|-80.66939|1.4079464610753885|46|1
35.28326|ffd535938d50ad71876fe71e67b14815b4a6188c|12.99|2015-02-11 12:47:00|80.669414401537693|3|4460031182|46|35.301105445937949|0|19|385|-80.814133|65|35.333742|NFS-CHARCOAL|2.31|1|KINGSFORD CHARCOAL|36462aa2eaa3d07ae740dc36bdebe3cbf48f3072|1.2330772300493043|35.305725790410776|00044600304519|CHARCOAL/LOGS/ACCESSORIES|G1 GROCERY|-80.66939|80.66939291321043|472|1
35.28326|5257fdbd801fcd1bdb4ecb1533f45287e59da2d5|2.39|2015-03-04 19:33:00|1.4094857484078087|3|7203695175|46|0.6158090578372145|0|26|1607|-80.66939|371|35.28326|FROZEN DOUGH (BREAD)|0.0|14|FRESH LRG FRENCH BREAD|36462aa2eaa3d07ae740dc36bdebe3cbf48f3072|1.2330772300493043|0.61471665291522548|00072036951755|BREAD|BAKERY|-80.66939|1.4079464610753885|46|1
35.28326|43b41003eb3ecd726237881d112391de94eec881|5.29|2014-12-15 18:04:00|1.4094857484078087|3|4460030984|46|0.6158090578372145|0|26|385|-80.66939|65|35.28326|NFS-CHARCOAL|0.0|1|KINGSFORD SMOKEHOUSE BRIQUETS|36462aa2eaa3d07ae740dc36bdebe3cbf48f3072|1.2330772300493043|0.61471665291522548|00044600309842|CHARCOAL/LOGS/ACCESSORIES|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|811bec9def6e1de81e261c8c9b750254797d7832|4.89|2014-12-15 14:47:00|1.4094857484078087|3|5000030212|46|0.6158090578372145|0|26|144|-80.66939|229|35.28326|CEAMERS-POWDERED|0.0|1|COFFEE MATE REGULAR|36462aa2eaa3d07ae740dc36bdebe3cbf48f3072|1.2330772300493043|0.61471665291522548|00050000302123|COCOAS CREAMERS SYRUPS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|84f3c82810ace160af15121ae804b1bd90985dd3|5.89|2015-01-29 19:04:00|1.4094857484078087|3|5210000295|46|0.6158090578372145|0|26|1245|-80.66939|34|35.28326|SINGLE SPICES|0.0|1|MC GOURMET MILD CURRY POWDER|36462aa2eaa3d07ae740dc36bdebe3cbf48f3072|1.2330772300493043|0.61471665291522548|00052100002958|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|8dd2b5239dd9449c10fde856115384493fd1b855|4.99|2014-12-20 17:59:00|1.4094857484078087|3|7203688117|46|0.6158090578372145|0|26|583|-80.66939|136|35.28326|NUTS|0.0|4|HT FILBERTS IN SHELL 1LB|36462aa2eaa3d07ae740dc36bdebe3cbf48f3072|1.2330772300493043|0.61471665291522548|00072036881175|OTHER MERCHANDISE|PRODUCE|-80.66939|1.4079464610753885|46|1
35.28326|3fd5dd14e5d72349de8b9b60497d308e0f45e315|11.99|2015-01-10 13:37:00|1.4094857484078087|3|8858600177|46|0.6158090578372145|0|26|9949|-80.66939|886|35.28326|NFS-PREM-MERLOT|0.0|13|14 HANDS MERLOT|36462aa2eaa3d07ae740dc36bdebe3cbf48f3072|1.2330772300493043|0.61471665291522548|00088586001772|PREMIUM ($8-$10.99)|WINE|-80.66939|1.4079464610753885|46|1
35.28326|f46b087dcf5dd534d1155ce9be1598415e3379b0|0.79|2015-02-14 11:52:00|1.4094857484078087|3||46|0.6158090578372145|0|26|524|-80.66939|64|35.28326|FRESH PROD FRESH ONIONS|0.0|4|COO GREEN ONIONS|36462aa2eaa3d07ae740dc36bdebe3cbf48f3072|1.2330772300493043|0.61471665291522548|00204068000006|FRESH PRODUCE|PRODUCE|-80.66939|1.4079464610753885|46|1
35.140781|e328e2579f71441b22724b54bc27324ea9835ac2|2.85|2014-10-09 13:16:00|1.4091206135396188|3|4112907700|39|0.6133223301722653|0|47|1219|-80.62331|275|35.140781|PASTA SC CORE|0.85|1|CLASSICO SC ROASTED GARLIC|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|0.61242566243833529|00041129077825|PASTA SAUCES|G1 GROCERY|-80.62331|1.4071422133560694|39|1
35.140781|0f848734c3832d294971269f2621fd54b77b6a50|2.99|2014-09-25 12:36:00|1.4091206135396188|3|7203663104|39|0.6133223301722653|0|47|364|-80.62331|55|35.140781|ORGANIC AND CF EGGS|0.0|3|HTN NEST GRADE A LARGE EGG BRO|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|0.61242566243833529|00072036631046|EGGS FRESH|DAIRY|-80.62331|1.4071422133560694|39|1
35.140781|e1de03498c4df92d4cfa228306abb01e8d7f006a|2.99|2014-10-03 16:01:00|1.4091206135396188|3|7203663104|39|0.6133223301722653|0|47|364|-80.62331|55|35.140781|ORGANIC AND CF EGGS|0.0|3|HTN NEST GRADE A LARGE EGG BRO|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|0.61242566243833529|00072036631046|EGGS FRESH|DAIRY|-80.62331|1.4071422133560694|39|1
35.140781|84550d53536af32e70381ffa7de1af7f8eaee0d1|2.99|2014-10-28 14:17:00|80.632521683083056|3|7203663104|39|35.178576094200288|0|39|364|-80.654118|55|35.123768|ORGANIC AND CF EGGS|0.0|3|HTN NEST GRADE A LARGE EGG BRO|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|35.177497916598789|00072036631046|EGGS FRESH|DAIRY|-80.62331|80.623324668201946|473|1
35.140781|2e803f663fdbc8ba5215c67c19e460f3b154bfc4|2.99|2014-09-15 14:44:00|1.4091206135396188|3|7203663104|39|0.6133223301722653|0|47|364|-80.62331|55|35.140781|ORGANIC AND CF EGGS|0.0|3|HTN NEST GRADE A LARGE EGG BRO|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|0.61242566243833529|00072036631046|EGGS FRESH|DAIRY|-80.62331|1.4071422133560694|39|1
35.140781|ec2c72c3ba4fa50868b8bcdcbd17e36b41e2e22d|1.54|2014-11-27 12:32:00|1.4091206135396188|3|7203632360|39|0.6133223301722653|0|47|1441|-80.62331|274|35.140781|MAC AND CHEESE|0.54|1|HT DIN MAC CHEESE|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|0.61242566243833529|00072036323606|PREP FOODS DINNERS|G1 GROCERY|-80.62331|1.4071422133560694|39|2
35.140781|90f67c2bfe1d59205bc21ff9ebc629fb920b9765|6.67|2015-02-22 13:14:00|1.4091206135396188|3|7203612054|39|0.6133223301722653|0|47|189|-80.62331|29|35.140781|TUNA-POUCH|1.6700000000000002|1|HT CHUNK WHITE TUNA POUCH|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|0.61242566243833529|00072036120557|SEAFOOD-CANNED|G1 GROCERY|-80.62331|1.4071422133560694|39|5
35.140781|cd1c2fdc1317cb4481b671a02b38280e38be376e|2.5|2015-02-15 19:32:00|1.4091206135396188|3|7203697755|39|0.6133223301722653|0|47|81|-80.62331|9|35.140781|RTE CEREAL KIDS|0.53|1|HT CER FROSTED FLAKES|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|0.61242566243833529|00072036977557|CEREAL|G1 GROCERY|-80.62331|1.4071422133560694|39|1
35.140781|c7152c732c92dcf6dd27006b9b43329bcea916b3|1.99|2015-01-01 21:06:00|1.4091206135396188|3|7940002522|39|0.6133223301722653|0|47|3545|-80.62331|1045|35.140781|SHAMPOO-VALUE|0.4|17|SUAVE SHAMPOO CHERRY BLOSSOM|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|0.61242566243833529|00079400025227|HAIR & SCALP CARE|HBC|-80.62331|1.4071422133560694|39|1
35.140781|af6c7bbaae7f04f71e9ac1c56ca1cdcf1cba90cb|3.29|2015-02-27 15:28:00|1.4091206135396188|3|7468000388|39|0.6133223301722653|0|47|78|-80.62331|11|35.140781|MUSTARD|1.65|1|D WOEBERS DIP HONEY MUSTARD|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|0.61242566243833529|00074680003880|CONDIMENTS|G1 GROCERY|-80.62331|1.4071422133560694|39|1
35.140781|677a80671164c637859a335446be999a43551643|3.29|2015-01-14 21:03:00|1.4091206135396188|3|65724360508|39|0.6133223301722653|0|47|244|-80.62331|43|35.140781|BETTER-FOR-YOU NOVELTIES|1.64|5|SOBE LW PACIFIC COCONUT POPS|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|0.61242566243833529|00657243611083|FROZEN NOVELTIES|FROZEN|-80.62331|1.4071422133560694|39|1
35.140781|1aa8956a5b3b7976f4eddc2ca76f537eeff1fa64|5.99|2015-02-28 21:35:00|1.4091206135396188|3|78978501962|39|0.6133223301722653|0|47|244|-80.62331|43|35.140781|BETTER-FOR-YOU NOVELTIES|2.0|5|SKINNY COW LF VAN/CHOC I/C SDW|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|0.61242566243833529|00789785019628|FROZEN NOVELTIES|FROZEN|-80.62331|1.4071422133560694|39|1
35.140781|5147a07fc1bbfdcb68fc1c33d39872107bd25b30|5.34|2015-02-24 18:56:00|1.4091206135396188|3|7203698754|39|0.6133223301722653|0|47|1265|-80.62331|57|35.140781|ALMOND MILK|1.34|3|HT ALMOND DRINK UNSWT ORIGINAL|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|0.61242566243833529|00072036707352|MILK|DAIRY|-80.62331|1.4071422133560694|39|2
35.140781|0cfc914151d0a4f88f2cd284d5fcd84749950fb5|2.28|2015-02-02 18:17:00|1.4091206135396188|3||39|0.6133223301722653|0|47|522|-80.62331|64|35.140781|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|0.61242566243833529|00204664000004|FRESH PRODUCE|PRODUCE|-80.62331|1.4071422133560694|39|1
35.140781|c875c217df91d9101ddce2462c7104bae5a10419|3.67|2015-02-12 09:02:00|80.632521683083056|3|7203655019|39|35.178576048718369|0|39|332|-80.770346|52|35.052812|STRING/SNACK|0.0|3|HT TWISTARELLA STRING CHEESE|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|35.177497916598789|00072036550224|CHEESE|DAIRY|-80.62331|80.623383204155886|40|1
35.140781|1aca5984322d08749d49e385dad3044964d738a4|2.99|2014-11-21 08:56:00|80.632521683083056|3|3400000542|39|35.178576027226278|0|39|727|-80.8062|7|35.037115|SEASONAL CANDY-SINGLE FAC|0.49|1|I/O(C14)HRSY KISSES CANE|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|35.177497916598789|00034000005420|CANDY|G1 GROCERY|-80.62331|80.623398257881504|27|1
35.140781|cc69545507f2f12db097322a59fc2d61f832fc52|5.69|2015-03-01 19:26:00|1.4091206135396188|3|4956802016|39|0.6133223301722653|0|47|579|-80.62331|136|35.140781|SOY/MEATLESS PRODUCTS|0.0|4|FYH GRAPESEED OIL VEGENAISE|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|0.61242566243833529|00049568020167|OTHER MERCHANDISE|PRODUCE|-80.62331|1.4071422133560694|39|1
35.140781|3696148f00e54fc9f4d176846f7afb5cb7696b43|2.65|2014-11-25 13:24:00|80.632521683083056|3|4119680548|39|35.178576027226278|0|39|1201|-80.8062|33|35.037115|RTS CANNED|0.65|1|PROG HH SW BLK BEAN VEGETABLE|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|35.177497916598789|00041196458930|SOUP|G1 GROCERY|-80.62331|80.623398257881504|27|1
35.140781|2fbfd09c96560c89bc192ef4a45267b273e7cc2f|4.45|2014-09-30 15:52:00|1.4091206135396188|3|8087800218|39|0.6133223301722653|0|47|3536|-80.62331|1045|35.140781|SHAMPOO-PREMIUM|1.11|17|PANTENE SH DLY MOIS RENEWAL|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|0.61242566243833529|00080878171262|HAIR & SCALP CARE|HBC|-80.62331|1.4071422133560694|39|1
35.140781|bafaae56637803f1b5a44fea13b51500b09bf631|8.99|2014-10-20 21:00:00|80.632521683083056|3|7203695528|39|35.178576094200288|0|39|1659|-80.654118|381|35.123768|VARIETY SINGLE LAYER|0.0|14|SGL LYR DBL FUDGE CAKE.|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|35.177497916598789|00072036955289|CAKES|BAKERY|-80.62331|80.623324668201946|473|1
35.140781|b346e559abda625d7b260611e29adfa494aab392|1.29|2014-10-01 12:15:00|80.632521683083056|3|2200000899|39|35.178576093773735|0|39|48|-80.826724|7|35.195689|REGISTER GUM|0.29|1|EXTRA PEPPERMINT 15|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|35.177497916598789|00022000008916|CANDY|G1 GROCERY|-80.62331|80.623326229471132|412|1
35.140781|a3b6028f643b737ba6a9f64ef12ffe13f153aa67|1.67|2015-02-12 14:44:00|80.632521683083056|3|7062244101|39|35.178576027226278|0|39|53|-80.8062|7|35.037115|THEATER BOX|0.0|1|GOETZE'S CARAML THEATER BX|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|35.177497916598789|00070622441017|CANDY|G1 GROCERY|-80.62331|80.623398257881504|27|1
35.140781|a72ca5c90455394e06d7755380133ab8add6b015|2.99|2014-10-21 16:32:00|1.4091206135396188|3|73692100006|39|0.6133223301722653|0|47|364|-80.62331|55|35.140781|ORGANIC AND CF EGGS|0.0|3|NEST FRSH CAGE FR LG BROWN EGG|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|0.61242566243833529|00736921000064|EGGS FRESH|DAIRY|-80.62331|1.4071422133560694|39|1
35.140781|a67e25b68086d86ac0dfb95d8255d605d5b5810e|4.99|2015-02-15 19:37:00|1.4091206135396188|3|71575620002|39|0.6133223301722653|0|47|504|-80.62331|64|35.140781|FRESH BERRIES|2.5|4|STRAWBERRIES 1LB CLAM|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|0.61242566243833529|00812049005102|FRESH PRODUCE|PRODUCE|-80.62331|1.4071422133560694|39|1
35.140781|0044f3b35ae75c3355e54584a8190ff84393abde|5.99|2015-03-02 13:50:00|80.632521683083056|3|7116434316|39|35.178576027226278|0|39|3530|-80.8062|1045|35.037115|SHAMPOO-MID PRICE|2.0|17|HASK ARGAN OIL REPAIR SHAMPOO|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|35.177497916598789|00071164343166|HAIR & SCALP CARE|HBC|-80.62331|80.623398257881504|27|1
35.140781|b9057d848ad3fd8892157028d09a5ebd594ca870|3.49|2015-01-27 13:07:00|80.632521683083056|3|81547301440|39|35.178576027226278|0|39|1455|-80.8062|61|35.037115|DRINKABLE YOGURT|0.0|3|GO WILD BANANA&BRY DRINKABLE|384e52db900c098acaa1c11aa987401c50a0ba13|2.6115498688113523|35.177497916598789|00815473014412|YOGURT|DAIRY|-80.62331|80.623398257881504|27|1
35.318911|bb662d81fc7244b7107eba12977fdd5628f6af59|4.37|2015-02-04 10:43:00|80.780380710856576|4||167|35.368943495561737|0|48|523|-80.737839|64|35.297134|FRESH POTATOES|0.0|4|COO RUSSET POTATOES, BULK|3a6d37c41d9d7945f15a9cacdcd4ed45498dc1fd|3.45712462088821|35.351085445956379|00204072000009|FRESH PRODUCE|PRODUCE|-80.780702|80.780703937243814|258|1
35.412407|75660d8b3a9073505fa5475e58fcc889ea1dc696|4.19|2014-10-21 17:02:00|80.607132136635443|4|5210007086|68|35.471770183813732|0|9|217|-80.746334|34|35.41832|EXTRACTS FOOD COLORING|0.0|1|E  MCCORMICK VANILLA EXTRACT|3d07fbfbf67321f228a6d4bd8fd60c5e43e4a66e|4.10185285312355|35.47365851958088|00052100070865|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.662946|80.662969235415986|190|1
35.116751|bd7266b517185e3e5232734777755b394039036e|4.23|2014-11-02 20:29:00|80.825044058860698|2|20337400000|294|35.142129089089273|0|29|641|-80.85013|137|35.175855|PREMIUM PORK|1.93|2|PORK LOIN BNLS BUTTERFLY CHOPS|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00203382000006|PORK|MEAT|-80.824767|80.824782523149324|218|1
35.116751|b9670cd08a9f8fe53aedaf1de4b434ad6bbce4e8|2.18|2014-09-19 20:21:00|80.825044058860698|2||294|35.142129090503893|0|29|522|-80.825175|64|35.152722|FRESH TOMATOES|0.36|4|RED H/H TOMATOES, BULK|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00204799000009|FRESH PRODUCE|PRODUCE|-80.824767|80.824778559575378|160|1
35.116751|26d4564dd2183ba3119d3eb41f3009666cb918ab|7.64|2014-09-30 19:46:00|80.825044058860698|2|20943400000|294|35.142129083887333|0|29|883|-80.826724|145|35.195689|SHRIMP FARM RAISED|4.08|12|31/40 CT EZ PEEL WHITE SHRIMP|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00209434000000|SHRIMP|SEAFOOD|-80.824767|80.824792213096345|412|1
35.116751|d7c39fca3ffc40397e996ec5969ae6c15a65e48f|1.81|2014-09-23 12:52:00|80.825044058860698|2||294|35.142129090503893|0|29|523|-80.825175|64|35.152722|FRESH POTATOES|0.42|4|COO SWEET POTATOES, BULK|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00204091000004|FRESH PRODUCE|PRODUCE|-80.824767|80.824778559575378|160|1
35.116751|e06bdbc22972606c702966f932752e48c3e8975a|2.45|2014-10-29 20:35:00|80.825044058860698|2|7203663217|294|35.142129089089273|0|29|330|-80.85013|55|35.175855|EGGS|0.0|3|HT GRADE A LARGE EGGS 18 CT|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00072036632173|EGGS FRESH|DAIRY|-80.824767|80.824782523149324|218|1
35.116751|3cef66f7ca9b24784f930ec1f8b427a078662511|3.0|2014-10-21 19:22:00|80.825044058860698|2|7203655029|294|35.142129089089273|0|29|331|-80.85013|52|35.175855|NATURAL SLICED|1.33|3|HT SWISS 2% SLICES CHEESE|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00072036983954|CHEESE|DAIRY|-80.824767|80.824782523149324|218|1
35.116751|f39b540b2b6c299989d8a8ae72ea521745033f92|3.23|2014-09-30 16:02:00|1.4091206135396188|2||294|0.6129029275530112|0|47|536|-80.824767|64|35.116751|FRESH SQUASH|1.34|4|BUTTERNUT SQUASH|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|0.61242566243833529|00204759000001|FRESH PRODUCE|PRODUCE|-80.824767|1.4106583013072596|294|1
35.116751|8a82bbcaa0734695803fc7b02f03a572064bcda8|12.99|2014-10-25 10:11:00|80.825044058860698|2|20506300000|294|35.142129090503893|0|29|2020|-80.825175|505|35.152722|CHEESE SPECIALTIES|0.0|6|SPECIALITY CHEESE|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00205063000008|SPECIALTY CHEESE|DELI|-80.824767|80.824778559575378|160|1
35.116751|f61e3cf58a4893127664e9409da1f21eb2714a2a|2.5|2014-10-04 20:21:00|80.825044058860698|2|78142100610|294|35.142129090503893|0|29|1601|-80.825175|371|35.152722|BRANDED BREAD|0.51|14|LA BREA WHEAT BAGUETTE|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00781421521182|BREAD|BAKERY|-80.824767|80.824778559575378|160|1
35.116751|738041c14d2a9bca9ffb138eb21bbe38ead87eb9|2.45|2014-09-13 20:35:00|80.825044058860698|2|74759960724|294|35.142129090503893|0|29|62|-80.825175|7|35.152722|SPECIALTY BAR/BOX CHOCOLATE|0.0|1|GHIRARDELLI HAZELNUT DARK BAR|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00747599611742|CANDY|G1 GROCERY|-80.824767|80.824778559575378|160|1
35.116751|83661425e85b37f0ff0ac8057b66df979d5890a7|1.15|2014-10-07 15:35:00|80.825044058860698|2|7203624020|294|35.142129089089273|0|29|149|-80.85013|23|35.175855|WHSE PASTA CORE|0.0|1|HT PASTA RIGATONI|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00072036240255|PASTA|G1 GROCERY|-80.824767|80.824782523149324|218|1
35.116751|f4103679f803b54928dc79f3587e9925d7883bc2|5.99|2014-11-01 20:36:00|80.825044058860698|2|7365700252|294|35.142129089089273|0|29|152|-80.85013|24|35.175855|NFS-CAT FOOD DRY|0.0|1|EVOLVE ADULT CAT FOOD BONUS|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00073657002628|PET FOOD/SUPPLIES|G1 GROCERY|-80.824767|80.824782523149324|218|1
35.116751|d6f892fa618cade8b3945fb04bed43a8bdb14368|2.99|2014-11-22 20:39:00|80.825044058860698|2|4145811704|294|35.142129089089273|0|29|265|-80.85013|307|35.175855|FROZEN PIES|0.0|5|EDWARDS CHOC SUNDAE SINGLES|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00041458117049|DESSERTS FROZEN|FROZEN|-80.824767|80.824782523149324|218|1
35.116751|4c73c810e3bac2acaa4343f807f4d77eea6b8ff8|6.99|2014-09-20 10:20:00|80.825044058860698|2|3798202150|294|35.142129090503893|0|29|2023|-80.825175|505|35.152722|GOAT CHEESE|2.0|6|GOAT CHEESE ORIGINAL|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00037982021501|SPECIALTY CHEESE|DELI|-80.824767|80.824778559575378|160|1
35.116751|d1ab99cec92d8323a565b28e2c8b06baa5bc4764|9.99|2014-09-16 13:47:00|80.825044058860698|2|7203695109|294|35.142129089089273|0|29|2019|-80.85013|505|35.175855|PRESSED COOKED CHEESE|5.0|6|IMPTD GRATED PECORINO ROMANO|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00072036951090|SPECIALTY CHEESE|DELI|-80.824767|80.824782523149324|218|1
35.116751|edfe72ee03584a221769636ebf05f7a68f3a287d|2.99|2014-11-19 21:45:00|80.825044058860698|2|7261371099|294|35.142129089089273|0|29|1513|-80.85013|66|35.175855|NFS-LAUNDRY DETERGENT PODS|0.49|1|SUN LAUNDRY PACS 20CT|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00072613711000|DETERGENTS|G1 GROCERY|-80.824767|80.824782523149324|218|1
35.116751|c77226a4f14c281a487ce85baf09b9e850d63a1a|1.29|2014-09-29 09:58:00|80.825044058860698|2||294|35.142129089089273|0|29|501|-80.85013|64|35.175855|FRESH PEARS|0.19|4|BARTLETT PEARS|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00204409000009|FRESH PRODUCE|PRODUCE|-80.824767|80.824782523149324|218|1
35.116751|a4b1741c8eeb8282fe4adcd3fd81ba1786bf9bf6|1.5|2014-11-21 21:59:00|80.825044058860698|2|980012301|294|35.142129083887333|0|29|47|-80.826724|7|35.195689|REGISTER BARS|0.25|1|ROCHER|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00009800123018|CANDY|G1 GROCERY|-80.824767|80.824792213096345|412|1
35.116751|c308043af8ad3dce692f166c9ef7a10d82efef6e|5.99|2014-11-15 21:04:00|80.825044058860698|2|7203695897|294|35.142129083887333|0|29|1654|-80.826724|381|35.195689|DESSERT CAKES|0.0|14|2 CT. TIRAMISU|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00072036958976|CAKES|BAKERY|-80.824767|80.824792213096345|412|1
35.116751|6d6a0a7673f937b2e34fdb19eac1a9d5330df957|1.69|2014-11-03 10:04:00|80.825044058860698|2|7203617993|294|35.142129089089273|0|29|5618|-80.85013|1512|35.175855|RUBBER/HOUSEHOLD GLOVES|0.0|18|(PPL) HT LATEX GLOVES LARGE|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00072036179937|BROOMS/MOPS & BRUSHES|GM|-80.824767|80.824782523149324|218|1
35.116751|198e7452b409a8daa9f4d31cacbcdafe73e3e32b|2.87|2014-11-29 10:19:00|80.825044058860698|2||294|35.142129090503893|0|29|562|-80.825175|64|35.152722|FRESH CUT FRUIT|0.0|4|CANTALOUPE SLICES|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00204487000007|FRESH PRODUCE|PRODUCE|-80.824767|80.824778559575378|160|1
35.116751|987b3c622dac876ae6f4c7a9d9a8a0069ce1f310|1.39|2014-11-05 12:04:00|80.825044058860698|2|8265750067|294|35.142129089089273|0|29|31|-80.85013|4|35.175855|NON CARBONATED WATER|0.39|1|DEER PARK WATER 1LT|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00082657500676|BOTTLED WATER|G1 GROCERY|-80.824767|80.824782523149324|218|1
35.116751|a18b76245c2469d76b6dc3dd16ca53d1d8c088e8|1.39|2014-09-21 12:27:00|1.4091206135396188|2|8265750067|294|0.6129029275530112|0|47|31|-80.824767|4|35.116751|NON CARBONATED WATER|0.39|1|DEER PARK WATER 1LT|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|0.61242566243833529|00082657500676|BOTTLED WATER|G1 GROCERY|-80.824767|1.4106583013072596|294|1
35.116751|a11ae34912eea1dbfb9632eab18573d46f415b36|1.19|2014-11-14 10:10:00|80.825044058860698|2|8265778540|294|35.142129089089273|0|29|30|-80.85013|4|35.175855|CARBONATED WATER|0.19|1|DEER PRK SPARKLIN ORANGE 1L|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00082657785400|BOTTLED WATER|G1 GROCERY|-80.824767|80.824782523149324|218|1
35.116751|34f7c0499224367000516112af4a772b2b2c1388|1.19|2014-11-17 09:51:00|80.825044058860698|2|8265778540|294|35.142129089089273|0|29|30|-80.85013|4|35.175855|CARBONATED WATER|0.19|1|DEER PRK SPARKLIN ORANGE 1L|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00082657785400|BOTTLED WATER|G1 GROCERY|-80.824767|80.824782523149324|218|1
35.116751|42add628f8419ddcf47e94cb2fa0978e2da8c7d4|0.99|2014-10-06 10:05:00|80.825044058860698|2|3400000031|294|35.142129089089273|0|29|47|-80.85013|7|35.175855|REGISTER BARS|0.5|1|HERSHEY KIT KAT BAR|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00034000002467|CANDY|G1 GROCERY|-80.824767|80.824782523149324|218|1
35.116751|cec85b1124650da34b3d66e4f9d140329a08d706|10.95|2014-11-23 19:39:00|80.825044058860698|2|20689700000|294|35.142129083887333|0|29|2027|-80.826724|510|35.195689|SOMETHING CLASSIC|0.0|6|SOMETHING CLASSIC ENTREES|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00206897000004|SOMETHING CLASSIC|DELI|-80.824767|80.824792213096345|412|1
35.116751|c60377198fed32050631e21ae41b57563ef03ae0|2.65|2014-09-19 10:03:00|80.825044058860698|2|1600026460|294|35.142129089089273|0|29|42|-80.85013|6|35.175855|GRANOLA/YOGURT BARS|0.0|1|NV BAR CRN DARK CHOCOLATE|40c97c0124ac9bdf11f89a4efc6d4cccae4ef120|1.753564889602039|35.157881615307893|00016000413146|BREAKFAST FOODS|G1 GROCERY|-80.824767|80.824782523149324|218|1
35.603432|a3c292c5671c890e643cc54f4e2fea2dc76803d7|15.12|2014-11-12 14:33:00|1.4102725052409182|4||274|0.6213971134099097|0|1|500|-80.895009|64|35.603432|FRESH APPLES|5.68|4|HONEY CRISP APPLE|43fee264cd5fed551520d587df9ad4765178dc5e|4.615879203105908|0.61833652052202714|00233283000003|FRESH PRODUCE|PRODUCE|-80.895009|1.4118842554804456|274|1
35.43259|460ea79d584cc6da6245703f23580298841c80c7|2.09|2014-10-29 17:11:00|1.4057311447477159|4||202|0.6184153580092175|0|52|522|-80.605588|64|35.43259|FRESH TOMATOES|0.0|4|RED H/H TOMATOES, BULK|44c4b2d4dec22ac53ea4936fb3eaf8769c1d54c1|2.3630384249102026|0.6209993146566879|00204799000009|FRESH PRODUCE|PRODUCE|-80.605588|1.406832906106031|202|1
35.43259|c5272ef5fa80f9a2cc46e34361990d486b8cf3fe|2.42|2014-09-30 17:11:00|1.4057311447477159|4||202|0.6184153580092175|0|52|522|-80.605588|64|35.43259|FRESH TOMATOES|0.81|4|RED H/H TOMATOES, BULK|44c4b2d4dec22ac53ea4936fb3eaf8769c1d54c1|2.3630384249102026|0.6209993146566879|00204799000009|FRESH PRODUCE|PRODUCE|-80.605588|1.406832906106031|202|1
35.43259|b96aed7079d8bb2956372ed4941974c72ff361e8|3.69|2014-10-09 17:09:00|1.4057311447477159|4|7518500003|202|0.6184153580092175|0|52|1033|-80.605588|163|35.43259|HAMBURGER|0.0|7|MARTIN'S POTATO SANDWICH ROLLS|44c4b2d4dec22ac53ea4936fb3eaf8769c1d54c1|2.3630384249102026|0.6209993146566879|00075185000039|BUNS/ROLLS|COMMERCIAL BAKERY|-80.605588|1.406832906106031|202|1
35.43259|8ae72b1c3ee24684616386d4794c651c7f9a90df|4.58|2014-10-16 08:38:00|1.4057311447477159|4|7203633079|202|0.6184153580092175|0|52|1244|-80.605588|21|35.43259|OTHER NUTS|0.0|1|HT DRY ROAST SUNFLOWER KERNEL|44c4b2d4dec22ac53ea4936fb3eaf8769c1d54c1|2.3630384249102026|0.6209993146566879|00072036330796|NUTS|G1 GROCERY|-80.605588|1.406832906106031|202|2
34.977331|77e02932d8ff8d013b51bfcb118225294acbdcd2|8.49|2014-09-16 19:25:00|81.02739863253349|4|2301290136|149|35.025958324813416|0|14|1477|-80.764523|485|35.341927|SUSHI HYBRID|0.0|6|CRUNCHY ROLL SP|4565aaf21cc92cd3fd8fc3decb5a4e9cbe346a36|3.3600723792267364|35.014943729270243|00023012901363|SUSHI|DELI|-81.027334|81.027629635881169|220|1
35.096737|1fb901f97c60cfc490854509dc05eeedb7b7d8cb|3.75|2014-12-19 18:40:00|80.782094729586973|1|4610000012|30|35.109195257698694|0|27|318|-80.825175|52|35.152722|SHREDDED/GRATED CHEESE|0.0|3|SARGENTO OTB MOZZ TRAD CUT|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00046100000120|CHEESE|DAIRY|-80.78468|80.784686084205291|160|1
35.096737|5f7da2ca65c4622513a230cee133fd0f2dc9b4e8|6.78|2015-01-09 19:05:00|80.782094729586973|1|5000012734|30|35.109195257698694|0|27|341|-80.825175|57|35.152722|CREAMERS|1.78|3|COFFEEMATE SF FRENCH VANILLA|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00050000848119|MILK|DAIRY|-80.78468|80.784686084205291|160|2
35.096737|d06ca65d7e246a2742724eb900fb72207716da4c|3.39|2014-10-25 13:51:00|80.782094729586973|1|5000012734|30|35.109195258692949|0|27|341|-80.806073|57|35.106477|CREAMERS|0.89|3|COFFEEMATE SF FRENCH VANILLA|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00050000848119|MILK|DAIRY|-80.78468|80.784680070686093|4|1
35.096737|33aa90c80a023a7473bf57a237aca4e250db3d32|3.69|2014-09-29 18:14:00|80.782094729586973|1|5000012734|30|35.109195257698694|0|27|341|-80.825175|57|35.152722|CREAMERS|1.19|3|COFFEEMATE SF FRENCH VANILLA|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00050000848119|MILK|DAIRY|-80.78468|80.784686084205291|160|1
35.096737|805d9d3cc70b534a01c8264b0b9ac0cb6f54339a|3.39|2014-11-22 18:06:00|80.782094729586973|1|5000012734|30|35.109195257698694|0|27|341|-80.825175|57|35.152722|CREAMERS|0.89|3|COFFEEMATE SF FRENCH VANILLA|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00050000848119|MILK|DAIRY|-80.78468|80.784686084205291|160|1
35.096737|a110fefe71a81f183f5a9da50aa4f20a5c42ee33|4.19|2014-11-16 13:05:00|80.782094729586973|1|4812110208|30|35.109195258692949|0|27|1037|-80.806073|164|35.106477|ENGLISH MUFFINS|0.0|7|THOMAS ENG MUFFN ORIG 6 PK PP|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00048121102081|BREAKFAST|COMMERCIAL BAKERY|-80.78468|80.784680070686093|4|1
35.096737|955a5fead57721bbb820b95ada59ca4ba35c60b0|3.39|2014-12-12 18:04:00|80.782094729586973|1|5000012734|30|35.109195258692949|0|27|341|-80.806073|57|35.106477|CREAMERS|0.89|3|COFFEEMATE SF FRENCH VANILLA|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00050000848119|MILK|DAIRY|-80.78468|80.784680070686093|4|1
35.096737|882be22a08edea723a6dd789dae1df8d67cb061d|9.98|2014-11-23 13:32:00|80.782094729586973|1|7002500010|30|35.109195257698694|0|27|361|-80.825175|105|35.152722|BREAKFAST SAUSAGE|0.0|19|NEESE COUNTRY SAUSAGE HOT|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00070025000118|BREAKFAST SAUSAGE|CASE READY MEATS|-80.78468|80.784686084205291|160|2
35.096737|9b3675509779c1d35839a551a78f59dcedd29871|9.98|2014-12-24 10:03:00|80.782094729586973|1|7002500010|30|35.109195257698694|0|27|361|-80.825175|105|35.152722|BREAKFAST SAUSAGE|0.0|19|NEESE COUNTRY SAUSAGE HOT|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00070025000118|BREAKFAST SAUSAGE|CASE READY MEATS|-80.78468|80.784686084205291|160|2
35.096737|6b60de39e336375b14718e5613dd32863167b7eb|4.99|2015-02-16 16:22:00|80.782094729586973|1|7002500010|30|35.109195258285972|0|27|361|-80.771677|105|35.066546|BREAKFAST SAUSAGE|0.0|19|NEESE COUNTRY SAUSAGE HOT|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00070025000118|BREAKFAST SAUSAGE|CASE READY MEATS|-80.78468|80.784683892975522|45|1
35.096737|dcecef39a2ee53470fb75f2facd49b0213cb8c28|10.99|2014-12-28 12:26:00|80.782094729586973|1|7203683001|30|35.109195258692949|0|27|352|-80.806073|110|35.106477|IQF CHICKEN|2.51|19|HT 2.5 LB CHICKEN TENDR BRST|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00072036830029|FROZEN CASE MEAT|CASE READY MEATS|-80.78468|80.784680070686093|4|1
35.096737|c0017ec3d7a67fb68bf6e306f32334640521cc95|10.99|2015-01-25 12:49:00|80.782094729586973|1|7203683001|30|35.109195258692949|0|27|352|-80.806073|110|35.106477|IQF CHICKEN|0.0|19|HT 2.5 LB CHICKEN TENDR BRST|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00072036830029|FROZEN CASE MEAT|CASE READY MEATS|-80.78468|80.784680070686093|4|1
35.096737|0213bc56d3b308c72b6a371447dfffa29625966a|5.99|2014-11-08 20:11:00|1.4091206135396188|1|7203695511|30|0.612553617356517|0|47|1677|-80.78468|383|35.096737|INDIVIDUALS (PASTRY CASE)|0.0|14|2 CT. RICOTTA CHEESECAKE|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|0.61242566243833529|00072036955111|PASTRY CASE|BAKERY|-80.78468|1.4099586511700126|30|1
35.096737|c518025f4f609c66c140e86d74cafeb740fed31c|5.99|2015-02-24 18:16:00|80.782094729586973|1|7203695511|30|35.109195258285972|0|27|1677|-80.771677|383|35.066546|INDIVIDUALS (PASTRY CASE)|0.0|14|2 CT. RICOTTA CHEESECAKE|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00072036955111|PASTRY CASE|BAKERY|-80.78468|80.784683892975522|45|1
35.096737|4a887be6ae7d9b4cb0dde7f9fcb2f9dd6a438b03|4.89|2015-01-06 16:53:00|80.782094729586973|1|7203670830|30|35.109195258285972|0|27|31|-80.771677|4|35.066546|NON CARBONATED WATER|1.1|1|(U)HT PURIFIED WATER .5L 32 PK|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00072036708304|BOTTLED WATER|G1 GROCERY|-80.78468|80.784683892975522|45|1
35.096737|e0bc69fa9b8535f2ceef1ccb703bc30b09884d00|4.89|2015-02-23 16:18:00|80.782094729586973|1|7203670830|30|35.109195258285972|0|27|31|-80.771677|4|35.066546|NON CARBONATED WATER|1.1|1|(U)HT PURIFIED WATER .5L 32 PK|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00072036708304|BOTTLED WATER|G1 GROCERY|-80.78468|80.784683892975522|45|1
35.096737|b30daadf5f0b3188a7f0348d6b3adf0efb312ca1|9.78|2014-11-04 13:02:00|80.782094729586973|1|7203670830|30|35.109195258285972|0|27|31|-80.771677|4|35.066546|NON CARBONATED WATER|2.2|1|(U)HT PURIFIED WATER .5L 32 PK|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00072036708304|BOTTLED WATER|G1 GROCERY|-80.78468|80.784683892975522|45|2
35.096737|352b8e91cca4342307b43d196f907c398f1b01aa|3.99|2015-02-01 10:24:00|80.782094729586973|1|7835470843|30|35.109195258692949|0|27|317|-80.806073|52|35.106477|CHUNK AND BAR CHEESE|0.4|3|CABOT MONTEREY JACK|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00078354702185|CHEESE|DAIRY|-80.78468|80.784680070686093|4|1
35.096737|8616fba5c03abc982a1a43dbd2df09799c2c091d|8.99|2015-01-04 13:25:00|80.782094729586973|1|7940041649|30|35.109195258285972|0|27|3776|-80.771677|1070|35.066546|CLINICAL-MALE|0.0|17|DEGREE MEN CLINICAL CLEAN DEO|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00079400206961|DEODORANT|HBC|-80.78468|80.784683892975522|45|1
35.096737|dbfb74fca0a48cb1d540c32d751f5b50d70014dd|1.47|2014-12-08 16:18:00|80.782094729586973|1|7203613030|30|35.109195258285972|0|27|101|-80.771677|15|35.066546|FLOUR-ALL PURPOSE|0.0|1|HARRIS TEETER ALL PRPOSE FLOUR|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00072036130303|FLOUR|G1 GROCERY|-80.78468|80.784683892975522|45|1
35.096737|5d5011943fb98e160750d5d6924547c20a061465|2.99|2015-02-15 12:24:00|80.782094729586973|1|7203628064|30|35.109195258692949|0|27|160|-80.806073|25|35.106477|OLIVES|0.0|1|HT OLIVES SPANISH QUEEN STFD 7|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00072036280640|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.78468|80.784680070686093|4|1
35.096737|d3e0521ad7344817003577c9c948fa79990315d8|1.54|2014-12-01 19:30:00|80.782094729586973|1|7203636010|30|35.109195257698694|0|27|30|-80.825175|4|35.152722|CARBONATED WATER|0.0|1|HT SIMPLY CLEAR PEACH|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00072036360137|BOTTLED WATER|G1 GROCERY|-80.78468|80.784686084205291|160|2
35.096737|27c74baf7b579ab048a1f5ea2356708ae5005a50|1.54|2014-11-02 13:29:00|80.782094729586973|1|7203636010|30|35.109195257698694|0|27|30|-80.825175|4|35.152722|CARBONATED WATER|0.1|1|HT SIMPLY CLEAR PEACH|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00072036360137|BOTTLED WATER|G1 GROCERY|-80.78468|80.784686084205291|160|2
35.096737|bcfd048332ef6e3cd12d8c614b827d0475d31817|0.77|2015-01-31 14:54:00|80.782094729586973|1|7203636010|30|35.109195257698694|0|27|30|-80.825175|4|35.152722|CARBONATED WATER|0.0|1|HT SIMPLY CLEAR PEACH|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00072036360137|BOTTLED WATER|G1 GROCERY|-80.78468|80.784686084205291|160|1
35.096737|bdb0d1c766c609a935395d63450e7a11bdf93419|2.69|2014-09-14 13:14:00|80.782094729586973|1|7203663996|30|35.109195258692949|0|27|342|-80.806073|57|35.106477|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00072036631299|MILK|DAIRY|-80.78468|80.784680070686093|4|1
35.096737|28c2e31bf08a126679daf700175f77f96d528dd0|0.97|2014-12-22 16:17:00|80.782094729586973|1|7203670024|30|35.109195258285972|0|27|4876|-80.771677|1235|35.066546|RUBBING ALCOHOL|0.0|17|HT ISO ALCOHOL 70%  -70024|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00072036700247|FIRST AID|HBC|-80.78468|80.784683892975522|45|1
35.096737|8efd39a4a07957d91b3f3780019ab1c2e9186152|5.69|2014-11-01 16:26:00|80.782094729586973|1|7756725423|30|35.109195258285972|0|27|252|-80.771677|45|35.066546|PREMIUM ICE CREAM|2.84|5|BREYERS COOKIES N' CREAM I/C|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00077567254504|ICE CREAM|FROZEN|-80.78468|80.784683892975522|45|1
35.096737|756f7f43a404689beeec31ca979b2f186ae0935a|4.99|2015-02-19 14:30:00|80.782094729586973|1|7940026654|30|35.109195256964284|0|27|3548|-80.816172|1045|35.059823|HAIR CARE SHPOO 2 IN 1'S|0.0|17|DOVE MEN 2N1 FRESH CLEAN HAIR|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00079400266545|HAIR & SCALP CARE|HBC|-80.78468|80.784688022300642|66|1
35.096737|ff6e735ad35507313a586df28052fe19948705ee|5.99|2014-11-11 17:42:00|80.782094729586973|1|8066095401|30|35.109195258285972|0|27|459|-80.771677|83|35.066546|IMPORT BEER|0.0|16|CORONITA 6PK 7OZ BTL|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00080660954011|IMPORT BEER|BEER|-80.78468|80.784683892975522|45|1
35.096737|56a9d19abb73f8302d0f92e848027bf9641073e1|5.99|2014-11-13 14:19:00|1.4091206135396188|1|8066095401|30|0.612553617356517|0|47|459|-80.78468|83|35.096737|IMPORT BEER|0.0|16|CORONITA 6PK 7OZ BTL|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|0.61242566243833529|00080660954011|IMPORT BEER|BEER|-80.78468|1.4099586511700126|30|1
35.096737|7a1b6bbab7f056870e243cf87cb20b3e61e970a6|16.01|2014-12-31 17:53:00|80.782094729586973|1|20396500000|30|35.109195258285972|0|27|978|-80.771677|202|35.066546|SMOKED MEATS|2.29|2|HT BNLS QTR SPIRAL HONEY HAM|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00203965000003|SMOKED HAMS|MEAT|-80.78468|80.784683892975522|45|1
35.096737|160fc9d8330ebf42f3ad7d76e96f5529c29a80a6|3.99|2014-12-20 12:34:00|80.782094729586973|1|1090000015|30|35.109195257698694|0|27|440|-80.825175|76|35.152722|NFS-ALUMINUM FOIL|0.99|1|REYNOLDS FOIL 75 FT|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00010900000154|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.78468|80.784686084205291|160|1
35.096737|dbb4e515d0bc5d573f0e0831d5bde135e3766e56|3.0|2014-11-19 17:06:00|80.782094729586973|1|7203632016|30|35.109195258285972|0|27|195|-80.771677|30|35.066546|SALAD & COOKING OIL|0.5|1|HT VEGETABLE OIL|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00072036320223|SHORTENING/OIL|G1 GROCERY|-80.78468|80.784683892975522|45|1
35.096737|67269b9b268a75460e7c5cb82965769b24761487|2.99|2015-02-22 14:18:00|80.782094729586973|1|7231000123|30|35.109195258692949|0|27|233|-80.806073|37|35.106477|BLACK TEA|0.49|1|BIGELOW TEA BLK CINNAMON STICK|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00072310001787|TEA|G1 GROCERY|-80.78468|80.784680070686093|4|1
35.096737|59341969bb5b315cb447e318a62207a3f4b84a71|3.59|2014-12-04 16:41:00|1.4091206135396188|1|7203695890|30|0.612553617356517|0|47|1654|-80.78468|381|35.096737|DESSERT CAKES|0.0|14|GRANDE FINALE CAKE SLICE|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|0.61242566243833529|00072036958907|CAKES|BAKERY|-80.78468|1.4099586511700126|30|1
35.096737|e68847ad280168f7a375d83b6bce4540510ce8a7|12.99|2014-10-08 13:17:00|80.782094729586973|1|7203697003|30|35.109195257698694|0|27|751|-80.825175|87|35.152722|NFS-BOUQUETS|0.0|9|TRADITIONAL BQT #1|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00072036970039|FLORAL|FLORAL|-80.78468|80.784686084205291|160|1
35.096737|466d2756da871f610d931362ec141b8e6632ab55|12.99|2015-02-15 07:17:00|80.782094729586973|1|7023666334|30|35.109195256964284|0|27|1153|-80.816172|87|35.059823|NFS-FRESH CUT ARRANGE|0.0|9|PETITE EXPRESSION ARR.|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00070236663348|FLORAL|FLORAL|-80.78468|80.784688022300642|66|1
35.096737|bf9e3b0f20ef87d93e7940a1b5c100aa4a55cdb7|2.49|2014-12-24 18:20:00|80.782094729586973|1|7203697776|30|35.109195257698694|0|27|442|-80.825175|76|35.152722|NFS-COOKING-STORAGE BAGS|1.02|1|YH SLIDER STORAGE BAGS QUART|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00072036977755|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.78468|80.784686084205291|160|1
35.096737|f21d21299dc271a30478a7ea33b1a942bb356c07|2.49|2014-11-07 15:37:00|80.782094729586973|1|7203697776|30|35.109195257698694|0|27|442|-80.825175|76|35.152722|NFS-COOKING-STORAGE BAGS|1.02|1|YH SLIDER STORAGE BAGS QUART|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00072036977755|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.78468|80.784686084205291|160|1
35.096737|4ff5a2e3852e2711a9045e0e4020364666509c0a|4.49|2014-11-14 15:26:00|1.4091206135396188|1|7203695755|30|0.612553617356517|0|47|1647|-80.78468|379|35.096737|PACKAGED MUFFINS|1.99|14|12CT MINI BLUEBERRY MUFFINS|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|0.61242566243833529|00072036957559|MUFFINS|BAKERY|-80.78468|1.4099586511700126|30|1
35.096737|9a67fb6b08e1d0b70d8388cb60ac4b1a556b9f1d|6.99|2014-10-24 15:19:00|80.782094729586973|1|1130066079|30|35.109195257698694|0|27|727|-80.825175|7|35.152722|SEASONAL CANDY-SINGLE FAC|0.7|1|I/O(H14)TROLLI GUMMI MIX|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00011300660795|CANDY|G1 GROCERY|-80.78468|80.784686084205291|160|1
35.096737|1cec8e4c66d5a50d4b33cd3150e64fb85bced66e|3.99|2015-02-18 20:43:00|80.782094729586973|1|87694000404|30|35.109195258285972|0|27|155|-80.771677|24|35.066546|NFS-DOG TREATS|0.0|1|VARIETY PET CHICKN&POTATO BIS|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00876940004060|PET FOOD/SUPPLIES|G1 GROCERY|-80.78468|80.784683892975522|45|1
35.096737|e3048734f1692684f462e4bf756ade3839cd209e|7.99|2014-11-14 16:59:00|80.782094729586973|1|73468919002|30|35.109195258285972|0|27|7314|-80.771677|1600|35.066546|CHRSTMS TREE SKRT/STOCKG IMP|1.5|18|"17"" PLUSH ADULT HAT"|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00734689190027|SEASONAL MERCHANDISE|GM|-80.78468|80.784683892975522|45|1
35.096737|9067309d6cf5275b2e37f5bc22aa04f2337f1c15|12.99|2015-02-08 14:46:00|80.782094729586973|1|7023666335|30|35.109195258692949|0|27|751|-80.806073|87|35.106477|NFS-BOUQUETS|0.0|9|EASTER JOY BOUQUET|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00070236663355|FLORAL|FLORAL|-80.78468|80.784680070686093|4|1
35.096737|f6c3dd1109f26a657d60ac7d1e52b8a47ab02f6e|6.05|2015-01-18 13:35:00|80.782094729586973|1||30|35.109195258692949|0|27|566|-80.806073|64|35.106477|SERVICE BAR|0.42|4|HT 7 LAYER MEXICAN BEAN DIP|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00204506000001|FRESH PRODUCE|PRODUCE|-80.78468|80.784680070686093|4|1
35.096737|50bb5ab8da0688f3f8de9d0b51b9ace38087d7a7|1.99|2015-02-15 14:39:00|80.782094729586973|1|60322422423|30|35.109195257698694|0|27|533|-80.825175|64|35.152722|FRESH PEPPERS|0.0|4|MINI SWEET PEPPERS 1LB|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00603224224230|FRESH PRODUCE|PRODUCE|-80.78468|80.784686084205291|160|1
35.096737|a41ef7dc16e1ddf74a6c2df58915498ff7150d7b|3.39|2014-10-03 12:48:00|80.782094729586973|1|3700011086|30|35.109195257698694|0|27|725|-80.825175|66|35.152722|NFS-DISHWASHING LIQUID|0.0|1|JOY ULTRA LIQ DISH LEMON SCNT|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00037000110866|DETERGENTS|G1 GROCERY|-80.78468|80.784686084205291|160|1
35.096737|fe55561fc590c1079ce603b3b3e82898f70c9ce4|10.63|2015-03-09 08:48:00|80.782094729586973|1||30|35.109195257698694|0|27|562|-80.825175|64|35.152722|FRESH CUT FRUIT|0.0|4|BERRY BLAST|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00204873000000|FRESH PRODUCE|PRODUCE|-80.78468|80.784686084205291|160|1
35.096737|6fa56068626391f23199ce9855ce2aa4145ac3a2|1.85|2014-09-12 12:36:00|80.782094729586973|1|7203663216|30|35.109195256182112|0|27|330|-80.709466|55|35.124987|EGGS|0.0|3|HT GRADE A    LARGE BROWN EGGS|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00072036632166|EGGS FRESH|DAIRY|-80.78468|80.784689668234805|157|1
35.096737|bb759eefb027d0e15bb2b8f34696f6241a1f3e07|8.35|2014-12-18 15:11:00|80.782094729586973|1|76211188813|30|35.109195257698694|0|27|37|-80.825175|10|35.152722|PODS/CUPS/SINGLES|1.36|1|STARBUCKS SUMATRA KCUP|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00762111888181|COFFEE|G1 GROCERY|-80.78468|80.784686084205291|160|1
35.096737|57a752944dda00717c52f7a4a49d422ca1d0a180|4.49|2014-09-21 12:41:00|80.782094729586973|1|2840009217|30|35.109195257698694|0|27|1981|-80.825175|480|35.152722|CHIPS|0.0|6|STACY'S PITA CHIPS NAKED|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00028400092173|DRY GOODS|DELI|-80.78468|80.784686084205291|160|1
35.096737|6db8c5feeeeedfdcd4b46c35a566b1ca3b1c9a07|18.99|2015-01-24 13:51:00|80.782094729586973|1|20640400000|30|35.109195257698694|0|27|1654|-80.825175|381|35.152722|DESSERT CAKES|0.0|14|"SPEC ORDER CHC 8"" ROUND 3 LYR"|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00206404000008|CAKES|BAKERY|-80.78468|80.784686084205291|160|1
35.096737|8c30b9dedd39a678da78c8c946d89cf01e1d504b|6.0|2015-03-04 18:46:00|80.782094729586973|1|20527500000|30|35.109195257698694|0|27|1945|-80.825175|465|35.152722|SUPERFLAG CHEF CASE|0.0|6|$6.00 CUSTOM COLD MEAL|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00205275000001|COLD PREPARED FOODS|DELI|-80.78468|80.784686084205291|160|1
35.096737|2333d790d4367e6b7085a803d1541e5f9e217625|16.59|2015-02-15 14:29:00|80.782094729586973|1|20496000000|30|35.109195257698694|0|27|755|-80.825175|87|35.152722|NFS-BALLOONS|0.0|9|*BALLOONS|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00204960000005|FLORAL|FLORAL|-80.78468|80.784686084205291|160|1
35.096737|f3e4d579fbb9596ceef36fd129b8cbc10e9256ae|6.0|2014-11-11 17:49:00|80.782094729586973|1|20527500000|30|35.109195257698694|0|27|1945|-80.825175|465|35.152722|SUPERFLAG CHEF CASE|0.0|6|$6.00 CUSTOM COLD MEAL|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00205275000001|COLD PREPARED FOODS|DELI|-80.78468|80.784686084205291|160|1
35.096737|004e5a059540bc511e77f518f6e486c8744aca88|6.0|2015-02-11 19:04:00|80.782094729586973|1|20527500000|30|35.109195257698694|0|27|1945|-80.825175|465|35.152722|SUPERFLAG CHEF CASE|0.0|6|$6.00 CUSTOM COLD MEAL|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00205275000001|COLD PREPARED FOODS|DELI|-80.78468|80.784686084205291|160|1
35.096737|2b6a7f592d83352275c63721ea0db5a1b1a5cf95|20.99|2014-10-20 16:56:00|80.782094729586973|1|20496100000|30|35.109195257698694|0|27|754|-80.825175|87|35.152722|NFS-SGLE STEM CUT FLOWER|0.0|9|*SINGLE STEM CUT FLOWERS|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00204961000004|FLORAL|FLORAL|-80.78468|80.784686084205291|160|1
35.096737|cd22011204ca665f36d86f43e4d8095c26031d91|2.8|2014-12-08 12:34:00|80.782094729586973|1|20584900000|30|35.109195257698694|0|27|1945|-80.825175|465|35.152722|SUPERFLAG CHEF CASE|0.0|6|S/F KALE SALAD|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00205538000007|COLD PREPARED FOODS|DELI|-80.78468|80.784686084205291|160|2
35.096737|a531cb09e2028791b94eccd06661f0b05ee77401|9.69|2014-10-09 12:53:00|80.782094729586973|1|31254715020|30|35.109195258285972|0|27|4484|-80.771677|1210|35.066546|HEMORRHOIDAL|0.0|17|TUCKS PADS|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00312547150200|STOMACH REMEDIES|HBC|-80.78468|80.784683892975522|45|1
35.096737|88739b0ef4ba3e2a9d812643ab4a2adf9e761bc6|6.0|2015-01-27 14:13:00|80.782094729586973|1|20527500000|30|35.109195257698694|0|27|1945|-80.825175|465|35.152722|SUPERFLAG CHEF CASE|0.0|6|$6.00 CUSTOM COLD MEAL|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00205275000001|COLD PREPARED FOODS|DELI|-80.78468|80.784686084205291|160|1
35.096737|6f07322ae54457d8991fcd050620b906487a35ae|1.32|2015-01-13 15:11:00|80.782094729586973|1||30|35.109195258285972|0|27|524|-80.771677|64|35.066546|FRESH PROD FRESH ONIONS|0.0|4|COO WHITE ONIONS, XL|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00204663000005|FRESH PRODUCE|PRODUCE|-80.78468|80.784683892975522|45|1
35.096737|5a4f95b9d4da0d2f9919429c003ad084c7367037|1.89|2014-10-20 14:21:00|80.782094729586973|1|1300079630|30|35.109195258285972|0|27|69|-80.771677|26|35.066546|CANNED GRAVY|0.0|1|HEINZ HS PORK GRAVY|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00013000798907|PREPARED FOODS-DRY MIXES|G1 GROCERY|-80.78468|80.784683892975522|45|1
35.096737|e4df131e1cd1167b62416f549e4c09d9d7cf1a78|0.85|2014-10-12 12:56:00|80.782094729586973|1|7203663222|30|35.109195258692949|0|27|330|-80.806073|55|35.106477|EGGS|0.0|3|HT GRADE A    LARGE EGGS 6 CT.|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00072036632227|EGGS FRESH|DAIRY|-80.78468|80.784680070686093|4|1
35.096737|32117fc13c7ef1e29d299605cc41b2e854a0aa0b|3.58|2015-02-18 17:59:00|80.782094729586973|1|5100001047|30|35.109195258285972|0|27|212|-80.771677|33|35.066546|CONDENSED SOUP|0.54|1|CAMP COND KID CHICKEN NOODLE O|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00051000016218|SOUP|G1 GROCERY|-80.78468|80.784683892975522|45|2
35.096737|e0154e709b665ba001fd89999b27c00ae391d58c|0.5|2014-11-15 14:19:00|80.782094729586973|1||30|35.109195257732374|0|27|509|-80.770346|64|35.052812|FRESH CITRUS-REMAINING|0.0|4|COO LIMES, LRG|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00204048000002|FRESH PRODUCE|PRODUCE|-80.78468|80.784685980271831|40|1
35.096737|994510de000c5956120a3fe3394b74b944088ca5|29.98|2014-12-28 12:32:00|80.782094729586973|1|88582402833|30|35.109195258692949|0|27|7287|-80.806073|1600|35.106477|CHRISTMAS PLUSH IMP|11.24|18|"I/O 12.5"" SITTNG TEDDY W/RIBBN"|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00885824028337|SEASONAL MERCHANDISE|GM|-80.78468|80.784680070686093|4|2
35.096737|820b301ec33d0147c1316ad583fe5dc5d90bb1c1|7.99|2015-02-21 09:42:00|80.782094729586973|1|5200020805|30|35.109195258285972|0|27|171|-80.771677|20|35.066546|ISOTONIC DRINKS|2.99|1|GATORADE FRUIT PUNCH 8PK|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00052000208061|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.78468|80.784683892975522|45|1
35.096737|6198d292bafad2b875b36bb385549fc67757e5be|3.59|2014-09-14 09:26:00|80.782094729586973|1|7203670716|30|35.109195258285972|0|27|427|-80.771677|72|35.066546|NFS-TOILET TISSUE|0.0|1|YH BATH ULTRA STRONG 4DR|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00072036707178|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.78468|80.784683892975522|45|1
35.096737|4c0d811f7db79b5c27f6f7c235b2814435640263|12.59|2015-01-14 14:38:00|80.782094729586973|1|515|30|35.109195258285972|0|27|33|-80.771677|10|35.066546|COFFEE BULK|0.0|1|HT TRADER BULK COFFEE PLU|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00000000005150|COFFEE|G1 GROCERY|-80.78468|80.784683892975522|45|1
35.096737|5d40201e187b601c013794fe91aa30747fd827da|6.99|2014-12-01 14:49:00|80.782094729586973|1|5000025117|30|35.109195258285972|0|27|341|-80.771677|57|35.066546|CREAMERS|0.81|3|COFFEMATE FRENCH VANILLA 64 OZ|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00050000350223|MILK|DAIRY|-80.78468|80.784683892975522|45|1
35.096737|351fccc1aff592489716607ff6d3553b0a82b656|12.99|2014-11-02 10:14:00|80.782094729586973|1|7023666311|30|35.109195258285972|0|27|751|-80.771677|87|35.066546|NFS-BOUQUETS|0.0|9|$12.99 SUNNY DAY BOUQUET|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00070236663119|FLORAL|FLORAL|-80.78468|80.784683892975522|45|1
35.096737|2b81c74c6c787f2ae0555a181e8ad322e7e654e1|17.98|2014-10-13 17:45:00|80.782094729586973|1|8224201284|30|35.109195257698694|0|27|9917|-80.825175|891|35.152722|NFS-OTHER WINE|0.0|13|GNARLY HEAD AUTHENTIC BLACK|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00082242012843|WINE REMAINING|WINE|-80.78468|80.784686084205291|160|2
35.096737|611f5fbf07933a41e2a958d4167afad44c217b00|7.98|2014-11-21 18:12:00|80.782094729586973|1|3400021303|30|35.109195257698694|0|27|46|-80.825175|7|35.152722|PKG CHOC|0.5|1|HERSHEY'S NUGGETS SP DARK/ALMD|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00034000032105|CANDY|G1 GROCERY|-80.78468|80.784686084205291|160|2
35.096737|3dff4711e87cf9d2a8e345985d32c350cfd65ebb|20.940000000000005|2014-10-14 09:12:00|80.782094729586973|1|7203695201|30|35.109195257698694|0|27|1639|-80.825175|377|35.152722|BULK (DONUTS)|0.5|14|6CT FRESH GLAZED DONUTS|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00072036952011|DONUTS|BAKERY|-80.78468|80.784686084205291|160|6
35.096737|fdc25e22b3f6099201afe5ed40af04553a20441c|6.99|2014-12-09 15:05:00|80.782094729586973|1|902112006|30|35.109195257698694|0|27|1191|-80.825175|87|35.152722|NFS-SEASONAL ITEMS|0.0|9|"6"" POINSETTIA  5 RED/3 COLOR"|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00009021120063|FLORAL|FLORAL|-80.78468|80.784686084205291|160|1
35.096737|15b50cafb75c2f01a32a9ea77b4b06c3b594cf43|3.98|2015-02-24 18:19:00|80.782094729586973|1|7203626076|30|35.109195258285972|0|27|427|-80.771677|72|35.066546|NFS-TOILET TISSUE|0.4|1|HT WIPE ALOE VIT WIPE REFIL 42|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00072036260765|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.78468|80.784683892975522|45|2
35.096737|281ab04d885b5a254bd5383f8f6cf737c6c1023a|10.99|2014-11-10 18:15:00|80.782094729586973|1|20310500000|30|35.109195258285972|0|27|1153|-80.771677|87|35.066546|NFS-FRESH CUT ARRANGE|0.0|9|*BUDVASE|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00203105000009|FLORAL|FLORAL|-80.78468|80.784683892975522|45|1
35.096737|6584306c990ac201b36dd074b97fc0572bf54bc4|10.99|2014-10-11 15:33:00|80.782094729586973|1|8500001819|30|35.109195257698694|0|27|9955|-80.825175|886|35.152722|NFS-PREM-MALBEC|0.0|13|ALAMOS MENDOZA MALBEC|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00085000018194|PREMIUM ($8-$10.99)|WINE|-80.78468|80.784686084205291|160|1
35.096737|a92a6debd3cc8adcf85474039867ef7e509baa22|4.79|2014-10-15 12:12:00|80.782094729586973|1|3700023756|30|35.109195257698694|0|27|427|-80.825175|72|35.152722|NFS-TOILET TISSUE|0.0|1|CHARMIN FRESHMATES REFILL 80CT|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00037000237563|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.78468|80.784686084205291|160|1
35.096737|7de22868e6a9a4dc8863dc425828e3b3dead6dc8|3.49|2015-01-10 14:19:00|80.782094729586973|1|7080095048|30|35.109195258692949|0|27|357|-80.806073|104|35.106477|SMOKED SAUSAGE ROPES|1.02|19|SMITHFIELD KIELBASA LOOP|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00070800950126|DINNER SAUSAGE|CASE READY MEATS|-80.78468|80.784680070686093|4|1
35.096737|f40231a6a6f2c607189d123cfc3ee749a84307f5|3.99|2014-12-27 14:12:00|80.782094729586973|1|87694000404|30|35.109195256964284|0|27|155|-80.816172|24|35.059823|NFS-DOG TREATS|0.0|1|VARIETY PET HMESTYL BUFFET BIS|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00876940004077|PET FOOD/SUPPLIES|G1 GROCERY|-80.78468|80.784688022300642|66|1
35.096737|f8f07aab170d4747d507d4d65d8ccd91c5fd038b|18.99|2015-01-18 12:25:00|80.782094729586973|1|8088749023|30|35.109195257698694|0|27|9954|-80.825175|886|35.152722|NFS-PREM-ZINFANDEL|0.0|13|BOGLE PHANTOM|48e103cb3ffeaaccee868c5251f3e9701eac8fa6|0.8608355900745744|35.102887530186244|00080887490231|PREMIUM ($8-$10.99)|WINE|-80.78468|80.784686084205291|160|1
35.341927|f7f3f66a769c4d6cc8875b53cd999f58df03b301|1.5|2014-10-11 14:34:00|80.77969194620016|3|7203663107|220|35.344906363411056|0|20|1262|-80.8955|57|35.4437|HALF N HALF WHIPPING CREAM|0.0|3|HT HALF & HALF|4aed850a56b6f8280aca4aa73b8179c379e6cb15|0.20586683869129868|35.345012799095393|00072036632036|MILK|DAIRY|-80.764523|80.764524684436509|272|1
35.341927|e36b5be54e756b00213408e1dce33dfd8e81a701|0.97|2014-12-30 19:31:00|80.77969194620016|3|7203670024|220|35.344906363411056|0|20|4876|-80.8955|1235|35.4437|RUBBING ALCOHOL|0.0|17|HT ISO ALCOHOL 70%  -70024|4aed850a56b6f8280aca4aa73b8179c379e6cb15|0.20586683869129868|35.345012799095393|00072036700247|FIRST AID|HBC|-80.764523|80.764524684436509|272|1
35.341927|7307fa4d91203806cb6ebdc1e08b0f0198ae3595|33.98|2014-12-13 13:44:00|80.77969194620016|3|7199031600|220|35.344906363411056|0|20|455|-80.8955|82|35.4437|DOMESTIC PREMIUM 12PK&>|0.0|16|COORS LIGHT 24PK 12OZ CAN|4aed850a56b6f8280aca4aa73b8179c379e6cb15|0.20586683869129868|35.345012799095393|00071990316006|DOMESTIC BEER|BEER|-80.764523|80.764524684436509|272|2
35.341927|d5f0dae9e53cd82058e7dda31b59b71934ba09a4|1.39|2015-01-25 10:53:00|80.77969194620016|3|5210076069|220|35.344906363727695|0|20|80|-80.995484|34|35.444064|SEASONING PACKETS|0.39|1|MC G M BAJA CITRUS MARINADE|4aed850a56b6f8280aca4aa73b8179c379e6cb15|0.20586683869129868|35.345012799095393|00052100351889|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.764523|80.764523040507896|121|1
35.341927|93c1c5e179a126a1fd10ceef646487402b067ece|6.99|2015-01-05 16:53:00|80.77969194620016|3|4900002890|220|35.344906363411056|0|20|55|-80.8955|8|35.4437|REGULAR|2.0|23|SPRITE 12OZ 12PK FRIDGE CAN|4aed850a56b6f8280aca4aa73b8179c379e6cb15|0.20586683869129868|35.345012799095393|00049000028928|CARBONATED BEVERAGES|BEVERAGE|-80.764523|80.764524684436509|272|1
35.500972|297fdc95a39f6e72e0037741b0c068aa6001735f|15.42|2015-02-28 16:59:00|80.849735164501183|4|20194200000|268|35.545232268575077|0|11|299|-80.875654|49|35.585842|ANGUS BEEF|0.0|2|ANGUS BEEF BNLS SHORT RIBS|4eb8fbcd3b05731f3293e90ca0e6d1227e456e27|3.0582786745622825|35.604954314503821|00201942000008|BEEF|MEAT|-80.860108|80.860151993813133|99|1
35.082768|0d608c76d0f96f885ec6043246c506fde373af29|1.95|2014-10-31 12:06:00|80.732732175546019|1|1450001098|147|35.10602424815545|0|35|1272|-80.771677|50|35.066546|BAG VEG STEAM|0.0|5|BE STEAMFRESH CUT GRN BEANS|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00014500011015|VEGETABLES-FROZEN|FROZEN|-80.732725|80.732734814989655|45|1
35.082768|c24921ea982df0d162e88bbadc893866fdd561d2|1.77|2014-11-10 15:59:00|80.732732175546019|1|7203657031|147|35.10602424815545|0|35|322|-80.771677|53|35.066546|SOUR CREAM|0.52|3|HT SOUR CREAM|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00072036570314|CULTURES|DAIRY|-80.732725|80.732734814989655|45|1
35.082768|e52b46c5fd27df41adc8b01f05d7708e72fb8a20|1.69|2014-09-16 12:44:00|80.732732175546019|1|7680828073|147|35.10602424815545|0|35|149|-80.771677|23|35.066546|WHSE PASTA CORE|0.69|1|BARILLA PASTA ROTINI|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00076808280982|PASTA|G1 GROCERY|-80.732725|80.732734814989655|45|1
35.082768|1a081fb0b639c25a220611423bbc169c7d5ad65a|5.29|2014-12-03 13:27:00|1.4091206135396188|1|7203670704|147|0.6123098123133061|0|47|252|-80.732725|45|35.082768|PREMIUM ICE CREAM|2.29|5|I/OHT ALL NATURAL PEPP BARK IC|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|0.61242566243833529|00072036707055|ICE CREAM|FROZEN|-80.732725|1.409051865357139|147|1
35.082768|d493dfa7f79269b46c21ff0787f1050d1f03f648|26.82|2014-11-17 12:49:00|80.732732175546019|1|20007200000|147|35.10602424815545|0|35|975|-80.771677|201|35.066546|POULTRY-FROZEN|10.12|2|16 X 20 H T PREMIUM TURKEY|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00200072000001|POULTRY|MEAT|-80.732725|80.732734814989655|45|1
35.082768|3e46b58cc3940fd7dbe961dbc2bb68fe346c6687|4.0|2014-11-26 11:14:00|80.732732175546019|1|65780295163|147|35.106024241539274|0|35|1165|-80.848528|87|35.053394|NFS-FRESH CONSUMER BUNCH|0.0|9|BUNCH- ALSTROEMERIA   RIVERD|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00657802951636|FLORAL|FLORAL|-80.732725|80.732748579853592|11|1
35.082768|5dc9db702b1c8aee87485e2c20dd3d0af3f838d7|1.5|2015-02-22 17:37:00|80.732732175546019|1||147|35.10602424815545|0|35|523|-80.771677|64|35.066546|FRESH POTATOES|0.3|4|COO SWEET POTATOES, BULK|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00204091000004|FRESH PRODUCE|PRODUCE|-80.732725|80.732734814989655|45|1
35.082768|4fc20bda904b3e7c768cae0bb7d8a9652130bd67|0.85|2015-01-02 11:40:00|80.732732175546019|1||147|35.106024249541903|0|35|523|-80.7007|64|35.06858|FRESH POTATOES|0.26|4|COO SWEET POTATOES, BULK|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00204091000004|FRESH PRODUCE|PRODUCE|-80.732725|80.732725080415094|273|1
35.082768|f795bda8b8e15f131c7d6c188ab75a17d12da729|3.99|2014-12-04 09:50:00|1.4091206135396188|1|7203695676|147|0.6123098123133061|0|47|1656|-80.732725|381|35.082768|CUP CAKES|0.0|14|FFM MINI VANILLA CUPCAKES|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|0.61242566243833529|00072036956767|CAKES|BAKERY|-80.732725|1.409051865357139|147|1
35.082768|58b42959f3621c64f1cd214cfe69d47900e58dad|1.69|2014-09-28 17:22:00|80.732732175546019|1|7203688003|147|35.10602424815545|0|35|527|-80.771677|64|35.066546|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00072036880031|FRESH PRODUCE|PRODUCE|-80.732725|80.732734814989655|45|1
35.082768|dd5d6058340520afa10e26a50e7799b8f387b515|6.99|2014-10-15 12:57:00|1.4091206135396188|1||147|0.6123098123133061|0|47|1347|-80.732725|64|35.082768|PUMPKINS|1.99|4|CARVING PUMPKINS, LARGE|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|0.61242566243833529|00204737000009|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|1
35.082768|f0d6f428eb338a0e6a0ece7573754bc04639a839|2.19|2014-09-26 10:51:00|80.732732175546019|1|64420941200|147|35.10602424815545|0|35|10|-80.771677|2|35.066546|LAYER CAKE MIX|0.0|1|D HINES SPICE CAKE MIX|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00644209410606|BAKING MIXES|G1 GROCERY|-80.732725|80.732734814989655|45|1
35.082768|c90be45ba739cfeb4cdf79113c04fa95ef6ccc74|4.99|2014-12-19 12:59:00|80.732732175546019|1|7403006610|147|35.10602424815545|0|35|332|-80.771677|52|35.066546|STRING/SNACK|2.5|3|SORRENTO CHEDDAR STICKSTERS|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00074030069207|CHEESE|DAIRY|-80.732725|80.732734814989655|45|1
35.082768|baf3a474f4b74286aa308b2cb982048bd04314f6|27.96|2015-01-26 12:00:00|1.4091206135396188|1|7203670967|147|0.6123098123133061|0|47|37|-80.732725|10|35.082768|PODS/CUPS/SINGLES|7.96|1|HT HOUSE BLEND DECAF K-CUPS|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|0.61242566243833529|00072036709691|COFFEE|G1 GROCERY|-80.732725|1.409051865357139|147|4
35.082768|cbe13fba771c2b49d8148bcc13276615ca646de9|5.18|2014-11-24 11:43:00|80.732732175546019|1|7173000720|147|35.10602424815545|0|35|150|-80.771677|23|35.066546|NOODLES/DUMPLINGS-DRY|1.29|1|NO YOLKS DUMPLINGS|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00071730007201|PASTA|G1 GROCERY|-80.732725|80.732734814989655|45|2
35.082768|00f042b21d5cdf58c8852dafb22989e319bef8bb|13.98|2015-02-13 14:38:00|80.732732175546019|1|7203670967|147|35.10602424815545|0|35|37|-80.771677|10|35.066546|PODS/CUPS/SINGLES|3.98|1|HT HOUSE BLEND DECAF K-CUPS|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00072036709691|COFFEE|G1 GROCERY|-80.732725|80.732734814989655|45|2
35.082768|e94ecf2217090d190a08eacf8ee1a0a442a912a1|3.89|2015-01-30 12:54:00|80.732732175546019|1|4812113545|147|35.10602424815545|0|35|1036|-80.771677|164|35.066546|BREAKFAST BAGELS|1.95|7|THOMAS 100% WHEAT BGL THIN PP|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00048121135461|BREAKFAST|COMMERCIAL BAKERY|-80.732725|80.732734814989655|45|1
35.082768|591c3e15af4975f25cd05b6520ee3707971db9b3|0.54|2015-03-06 18:01:00|1.4091206135396188|1||147|0.6123098123133061|0|47|522|-80.732725|64|35.082768|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|0.61242566243833529|00204664000004|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|1
35.082768|82a0b708c52cc20db68d5478f808324bdce5db0c|12.23|2014-09-21 13:52:00|80.732732175546019|1|20895300000|147|35.10602424815545|0|35|977|-80.771677|201|35.066546|FRESH HT CHICKEN|6.12|2|HT FRESH BNLS CHICKEN BREAST|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00208953000003|POULTRY|MEAT|-80.732725|80.732734814989655|45|1
35.082768|991367151471dd23dc32904b6ff858066f7356c5|5.19|2014-12-09 10:23:00|80.732732175546019|1|30573055807|147|35.10602424815545|0|35|4484|-80.771677|1210|35.066546|HEMORRHOIDAL|0.0|17|PREPARATION H MED. WIPES-55607|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00305730558075|STOMACH REMEDIES|HBC|-80.732725|80.732734814989655|45|1
35.082768|3e54e140cf1af18ec136ddb7a05effa9c7efc35d|8.79|2014-12-06 12:14:00|80.732732175546019|1|30573288310|147|35.10602424815545|0|35|4484|-80.771677|1210|35.066546|HEMORRHOIDAL|0.0|17|PREPARATION H SUPP-88310|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00305732883106|STOMACH REMEDIES|HBC|-80.732725|80.732734814989655|45|1
35.082768|214b968c30c3762d3e30692aba5b44475822a662|22.98|2015-01-09 13:14:00|1.4091206135396188|1|3700086344|147|0.6123098123133061|0|47|1205|-80.732725|67|35.082768|NFS-JUMBO DIAPERS|5.0|1|PAMP SWADDLER JUMBO PK SIZE 4|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|0.61242566243833529|00037000863458|DISPOSABLE DIAPERS|G1 GROCERY|-80.732725|1.409051865357139|147|2
35.082768|247ddc57ec665dc213b1528fb75e471e8fa00c3d|3.18|2014-09-24 13:53:00|1.4091206135396188|1|7090050126|147|0.6123098123133061|0|47|1221|-80.732725|275|35.082768|PASTA SC VALUE|0.68|1|DEI FRTLI PIZZA SAUCE|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|0.61242566243833529|00070900501266|PASTA SAUCES|G1 GROCERY|-80.732725|1.409051865357139|147|2
35.082768|b5dcebbd9fdfe2e1319b58a43727520014593944|2.2|2014-10-09 11:17:00|1.4091206135396188|1||147|0.6123098123133061|0|47|500|-80.732725|64|35.082768|FRESH APPLES|0.0|4|RED DEL APPLE, WA  48|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|0.61242566243833529|00233284000002|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|1
35.082768|c14ee73eadee615234a331754c5ffa49d13c2a70|4.19|2015-01-15 18:26:00|1.4091206135396188|1|5215900001|147|0.6123098123133061|0|47|690|-80.732725|61|35.082768|ORGANIC|0.0|3|STONYFIELD ORGANIC WM PLAIN|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|0.61242566243833529|00052159000011|YOGURT|DAIRY|-80.732725|1.409051865357139|147|1
35.082768|9be93efb714730c2f92fdba2f6855fd68a9fcd6b|2.29|2014-10-12 18:05:00|80.732732175546019|1|1800000260|147|35.10602424815545|0|35|325|-80.771677|54|35.066546|BISCUITS-REFRIGERATED|0.79|3|GRANDS BUTTERMILK BISCUITS|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00018000001828|DOUGH PRODUCTS|DAIRY|-80.732725|80.732734814989655|45|1
35.082768|f8b16a83f64133728110c793dd1b1d073e939b50|6.59|2014-12-08 13:06:00|80.732732175546019|1|7192196239|147|35.10602424815545|0|35|284|-80.771677|892|35.066546|SUPER PREMIUM PIZZA|1.59|5|DIGIORNO 12in TC PEPPERONI|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00071921006594|FROZEN PIZZA|FROZEN|-80.732725|80.732734814989655|45|1
35.082768|219908a8912bb039cfd5154312233ae7f12f8379|6.79|2014-12-29 16:32:00|80.732732175546019|1|4900002890|147|35.106024249541903|0|35|54|-80.7007|8|35.06858|DIET|1.8|23|FRESCA 12OZ 12PK FRIDGEPACK CN|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00049000031058|CARBONATED BEVERAGES|BEVERAGE|-80.732725|80.732725080415094|273|1
35.082768|086f3fa9d3aee37375b91bb73109a47234560581|8.58|2014-11-09 14:26:00|80.732732175546019|1|4400002747|147|35.10602424815545|0|35|91|-80.771677|13|35.066546|SPRAYED BUTTER CRACKERS|2.15|1|RITZ CRACKERS|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00044000031114|CRACKERS|G1 GROCERY|-80.732725|80.732734814989655|45|2
35.082768|441d62d4dc8798be8b901a8e8f18c2ebedbe4444|7.98|2014-10-18 13:45:00|80.732732175546019|1|4000015140|147|35.10602424815545|0|35|46|-80.771677|7|35.066546|PKG CHOC|0.98|1|SNICKERS FUN SIZE|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00040000151401|CANDY|G1 GROCERY|-80.732725|80.732734814989655|45|2
35.082768|48cc9513763b35eb7f76163b2027ef502180de8a|1.17|2014-09-25 12:19:00|80.732732175546019|1|7203690021|147|35.10602424815545|0|35|1033|-80.771677|163|35.066546|HAMBURGER|0.0|7|H T HAMBURGER BUNS|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00072036900210|BUNS/ROLLS|COMMERCIAL BAKERY|-80.732725|80.732734814989655|45|1
35.082768|d9c2368c73673b9a91dd7e365261db0e1e19bff6|1.94|2014-11-26 13:31:00|1.4091206135396188|1|7203671102|147|0.6123098123133061|0|47|1025|-80.732725|162|35.082768|WHITE|0.0|7|HT OLD FASHIONED BREAD|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|0.61242566243833529|00072036711021|SLICED BREAD|COMMERCIAL BAKERY|-80.732725|1.409051865357139|147|2
35.082768|caab40e9e83ddcc6b19b4b9e1c5850683d218bd8|4.69|2014-10-07 11:54:00|80.732732175546019|1|7203695754|147|35.10602424815545|0|35|1603|-80.771677|371|35.066546|PRIVATE LABEL BREAD|0.0|14|BAND OF BAKERS ROASTED GARLIC|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00072036957542|BREAD|BAKERY|-80.732725|80.732734814989655|45|1
35.082768|33e240a0726ef5cb24a88cee32e55b604451e93d|8.58|2014-12-13 13:47:00|80.732732175546019|1|2840015938|147|35.10602424815545|0|35|201|-80.771677|31|35.066546|POTATO CHIPS|3.58|1|XXL RUFFLES SR CRM & ONION|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00028400159630|SNACKS|G1 GROCERY|-80.732725|80.732734814989655|45|2
35.082768|70260e5316a068cc379fd386e37e3469e39b5102|0.94|2014-12-20 11:45:00|1.4091206135396188|1|7248600220|147|0.6123098123133061|0|47|11|-80.732725|2|35.082768|MUFFIN MIXES|0.0|1|JIFFY CORN MUFFIN MIX|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|0.61242566243833529|00072486002205|BAKING MIXES|G1 GROCERY|-80.732725|1.409051865357139|147|2
35.082768|81cdd64062607a06282cabdaf4fb7ddbf7e0864b|2.29|2015-03-02 15:33:00|80.732732175546019|1|7203663996|147|35.10602424815545|0|35|342|-80.771677|57|35.066546|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00072036631299|MILK|DAIRY|-80.732725|80.732734814989655|45|1
35.082768|e020546754cdba28f5566bcf44deabe2520d8646|4.58|2015-02-03 18:23:00|1.4091206135396188|1|7203663996|147|0.6123098123133061|0|47|342|-80.732725|57|35.082768|FRESH MILK|0.82|3|HARRIS TEETER FF SKIM MILK|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|0.61242566243833529|00072036631299|MILK|DAIRY|-80.732725|1.409051865357139|147|2
35.082768|60a61e90ca1b33fba0174c743c0ea60bce2b2422|3.99|2014-12-02 12:08:00|80.732732175546019|1|7203663995|147|35.10602424815545|0|35|342|-80.771677|57|35.066546|FRESH MILK|1.52|3|HARRIS TEETER FF SKIM MILK|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00072036631282|MILK|DAIRY|-80.732725|80.732734814989655|45|1
35.082768|9d67873092f8ab2296caad30755cbeeaacb1a419|8.99|2014-10-29 14:05:00|1.4091206135396188|1|2301290142|147|0.6123098123133061|0|47|1477|-80.732725|485|35.082768|SUSHI HYBRID|0.0|6|CRUNCHY DRAGON ROLL SP|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|0.61242566243833529|00023012901424|SUSHI|DELI|-80.732725|1.409051865357139|147|1
35.082768|ade3140fa349f509e528693db4d7a206b7504f62|7.18|2015-01-16 14:05:00|80.732732175546019|1|4000024906|147|35.106024246084409|0|35|46|-80.709466|7|35.124987|PKG CHOC|2.12|1|M&M DARK CHOC PEANUT|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00040000236153|CANDY|G1 GROCERY|-80.732725|80.73274049919165|157|2
35.082768|efb8f7c8ff3b58aaaa131fccd8d5ed814f644e91|7.38|2014-10-07 19:27:00|80.732732175546019|1|71514172928|147|35.106024249541903|0|35|330|-80.7007|55|35.06858|EGGS|0.0|3|EGGLAND BEST GRADE A EX-LG EGG|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00715141729283|EGGS FRESH|DAIRY|-80.732725|80.732725080415094|273|2
35.082768|a843e439610787695ebfbd024c85ebbe3bb034b0|1.79|2015-02-18 13:36:00|80.732732175546019|1|7056097906|147|35.10602424815545|0|35|1272|-80.771677|50|35.066546|BAG VEG STEAM|0.0|5|PCTSWT STEAMABLES GRN PEAS|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00070560979016|VEGETABLES-FROZEN|FROZEN|-80.732725|80.732734814989655|45|1
35.082768|a24826388f9f81d1c63d628d6b7f455c0fcd99fd|4.89|2014-12-22 15:56:00|1.4091206135396188|1|74236526435|147|0.6123098123133061|0|47|345|-80.732725|57|35.082768|ORGANIC MILK|0.0|3|HORIZON WHOLE  DHA|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|0.61242566243833529|00742365264474|MILK|DAIRY|-80.732725|1.409051865357139|147|1
35.082768|482802079a7b358a7b0cb0aa6f2f416ecd9826a9|3.99|2014-11-14 11:29:00|80.732732175546019|1|7835470843|147|35.10602424815545|0|35|317|-80.771677|52|35.066546|CHUNK AND BAR CHEESE|1.49|3|CABOT SERIOUSLY SHARP|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00078354708439|CHEESE|DAIRY|-80.732725|80.732734814989655|45|1
35.082768|6d8e9fb575681740b337bd3fd5581a1489091277|6.78|2014-10-07 19:29:00|80.732732175546019|1|71514150349|147|35.106024249541903|0|35|330|-80.7007|55|35.06858|EGGS|1.78|3|EGGLAND BEST GRADE A LARGE EGG|51b93baff4d94658190ffcf3da631d9c8470e01d|1.606950681519739|35.101032182271901|00715141503494|EGGS FRESH|DAIRY|-80.732725|80.732725080415094|273|2
35.23102|72772f52bd92a92ca42d7bd43ca86f357be4987e|3.99|2014-12-09 22:25:00|80.843809562956082|4|4300095117|205|35.269468301924427|0|37|209|-80.737839|20|35.297134|POWDERED SOFT DRINKS|0.0|1|COUNTRY TIME LEMONADE (8QT)|535f7cc5ecefc0811c442203aa3d123f287c49f4|2.656686627400627|35.255745041786184|00043000951170|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.8438|80.843855014934022|258|1
35.103409|db625d395bc937ece331766129c7404b3d16be1d|4.69|2015-01-02 11:53:00|1.4132775322775095|4|1600043779|88|0.6126700657242101|0|58|1433|-80.992182|9|35.103409|GRANOLA|0.0|1|NV PROTEIN GRANOLA OATS HONEY|544677dfe1fc7c550335646875c3a6b360c70bf6|5.844925944913263|0.61177642288969325|00016000437791|CEREAL|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|445bd02fdfee14ba4e6e5da316c021843b8aa03c|11.07|2014-10-09 13:24:00|1.4132775322775095|4|1630015352|88|0.6126700657242101|0|58|139|-80.992182|20|35.103409|REMAINING SHELF STABLE JUICES|0.0|1|DD UNSWEET ORANGE JUICE 6PK|544677dfe1fc7c550335646875c3a6b360c70bf6|5.844925944913263|0.61177642288969325|00016300153520|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.992182|1.413580244274486|88|3
35.103409|bef038b9ea9beca084293356d045bfd4087536b0|5.38|2015-02-27 14:43:00|80.992238315890603|4|7203688023|88|35.187998347416219|0|22|555|-81.027334|64|34.977331|PACKAGED SALADS|0.0|4|HT CURLY SPINACH,PKG|544677dfe1fc7c550335646875c3a6b360c70bf6|5.844925944913263|35.131650835559327|00072036880239|FRESH PRODUCE|PRODUCE|-80.992182|80.992334061404662|149|2
35.103409|bcae5239b3588cb45794b34de07bc57284ae0599|5.38|2015-01-23 14:21:00|80.992238315890603|4|7203688023|88|35.187998347416219|0|22|555|-81.027334|64|34.977331|PACKAGED SALADS|0.0|4|HT CURLY SPINACH,PKG|544677dfe1fc7c550335646875c3a6b360c70bf6|5.844925944913263|35.131650835559327|00072036880239|FRESH PRODUCE|PRODUCE|-80.992182|80.992334061404662|149|2
35.103409|ffc62b2ce57431e87ee4c14ef9d661f9d5fc41cc|4.98|2014-09-20 16:06:00|1.4132775322775095|4|7203688048|88|0.6126700657242101|0|58|526|-80.992182|64|35.103409|FRESH MUSHROOMS|0.49|4|HT SLICED BABY BELLAS|544677dfe1fc7c550335646875c3a6b360c70bf6|5.844925944913263|0.61177642288969325|00072036880482|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|2
35.103409|176a21685c67027c2953f9e72e399aa933d24cb1|9.98|2015-01-19 11:53:00|80.992238315890603|4|4082201114|88|35.18799840660671|0|22|1878|-80.806073|435|35.106477|HUMMUS|2.49|6|HUMMUS W/ ROASTED PINE NUTS|544677dfe1fc7c550335646875c3a6b360c70bf6|5.844925944913263|35.131650835559327|00040822011747|SALADS|DELI|-80.992182|80.992272254348734|4|2
35.103409|3e5e9f4289235064f0cb9c6086eb4a748f0b8a0c|6.26|2014-10-30 13:11:00|1.4132775322775095|4|20598500000|88|0.6126700657242101|0|58|1821|-80.992182|410|35.103409|BH TURKEY|0.0|6|BOARS HEAD NO SALT TURKE|544677dfe1fc7c550335646875c3a6b360c70bf6|5.844925944913263|0.61177642288969325|00205985000001|BH MEAT|DELI|-80.992182|1.413580244274486|88|1
35.103409|48d4508d9516bd09d3d47f445a7a7d1ae73ec37c|5.99|2014-12-01 12:08:00|80.992238315890603|4|5440000004|88|35.187998347416219|0|22|76|-81.027334|11|34.977331|MEAT SAUCES|0.0|1|A1 STEAK SAUCE 15 OZ|544677dfe1fc7c550335646875c3a6b360c70bf6|5.844925944913263|35.131650835559327|00054400000047|CONDIMENTS|G1 GROCERY|-80.992182|80.992334061404662|149|1
35.103409|118e05b3afc10c4f747fb77afe1bb662eed038e0|9.99|2014-11-20 15:58:00|80.992238315890603|4|8992427896|88|35.187998430429687|0|22|455|-80.994596|82|35.061685|DOMESTIC PREMIUM 12PK&>|0.0|16|YUENGLING LAGER 12PK 12OZ BTL|544677dfe1fc7c550335646875c3a6b360c70bf6|5.844925944913263|35.131650835559327|00089924278962|DOMESTIC BEER|BEER|-80.992182|80.992228021476535|475|1
35.103409|333c40e28efce55ce96044ac2be2ebfd2042f242|5.49|2014-10-20 15:43:00|1.4132775322775095|4|2301290003|88|0.6126700657242101|0|58|1483|-80.992182|485|35.103409|SUSHI ROLL AND WRAP|0.0|6|avocado salad roll|544677dfe1fc7c550335646875c3a6b360c70bf6|5.844925944913263|0.61177642288969325|00023012900038|SUSHI|DELI|-80.992182|1.413580244274486|88|1
35.103409|f2605482a3368662b45f31f0c2febed3e891440a|4.29|2015-01-12 13:50:00|1.4132775322775095|4|2840015938|88|0.6126700657242101|0|58|201|-80.992182|31|35.103409|POTATO CHIPS|2.15|1|RUFFLES REGULAR|544677dfe1fc7c550335646875c3a6b360c70bf6|5.844925944913263|0.61177642288969325|00028400159388|SNACKS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|237fa65279d38f4cac31054432161f55607ca857|3.55|2014-12-04 16:41:00|1.4132775322775095|4|7433610102|88|0.6126700657242101|0|58|342|-80.992182|57|35.103409|FRESH MILK|0.0|3|HIGHLAND CREST 2% REDUCE FAT|544677dfe1fc7c550335646875c3a6b360c70bf6|5.844925944913263|0.61177642288969325|00074336101021|MILK|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|a70cb57414c8a368b321a571d982b3bb00fd0112|2.69|2014-12-08 16:40:00|80.992238315890603|4|7225001739|88|35.187998347416219|0|22|1025|-81.027334|162|34.977331|WHITE|0.5|7|NATOWN WHITEWHEAT RTOP BRD|544677dfe1fc7c550335646875c3a6b360c70bf6|5.844925944913263|35.131650835559327|00072250017398|SLICED BREAD|COMMERCIAL BAKERY|-80.992182|80.992334061404662|149|1
35.103409|1236a0188e732c41ab3fa357eb39d2c163035feb|8.59|2014-11-08 16:57:00|1.4132775322775095|4|76211120604|88|0.6126700657242101|0|58|36|-80.992182|10|35.103409|PREMIUM GROUND|1.6|1|STARBUCKS CAFFE VERONA GROUND|544677dfe1fc7c550335646875c3a6b360c70bf6|5.844925944913263|0.61177642288969325|00762111622877|COFFEE|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|33b1a0f4edde7ba87e4bad2aa878f9444b692d42|10.49|2015-03-05 15:43:00|1.4132775322775095|4|20956600000|88|0.6126700657242101|0|58|664|-80.992182|145|35.103409|SHRIMP WILD CAUGHT|0.0|12|WC E. COAST SHRIMP MEDIUM (US)|544677dfe1fc7c550335646875c3a6b360c70bf6|5.844925944913263|0.61177642288969325|00209566000008|SHRIMP|SEAFOOD|-80.992182|1.413580244274486|88|1
34.95459|31ffdc0cb5b4a46185c666342927d7049e9bfa6c|8.99|2015-01-07 13:12:00|80.801203185414451|4|3160404104|182|35.221009130224346|0|24|4612|-80.816172|1215|35.059823|VITAMIN-MINERALS|4.5|17|VITAMELTS ZINC 15 MG|558f4ba59498ff0fafe33132786933463393e619|18.408924957971134|35.194272495053255|00031604041045|VITAMINS & SUPPLEMENTS|HBC|-80.758228|80.758500311755526|66|1
34.95459|978f7e1be3c9c502133d27cd995c8ac3e2492dfa|3.59|2014-10-15 10:40:00|80.801203185414451|4|7940018420|182|35.221009171710413|0|24|3816|-80.848528|1070|35.053394|INVISIBLE-MALE|0.0|17|DEGREE COOL COMFORT INV SOLID|558f4ba59498ff0fafe33132786933463393e619|18.408924957971134|35.194272495053255|00079400205704|DEODORANT|HBC|-80.758228|80.758430828110022|11|1
35.024332|eba6925e31773b99584b3afe8f6363902c950854|7.96|2015-01-10 15:11:00|80.805842308733688|4|20896500000|343|35.040147321607122|0|49|977|-80.837892|201|34.937113|FRESH HT CHICKEN|0.0|2|HT FRESH CHICKEN DRUMMETTES|592d68633407db752e5164652722ae9032819632|1.0928013930929041|35.053350220983141|00208965000008|POULTRY|MEAT|-80.760919|80.760943269058956|372|2
35.585842|e5490caa2d56ae01e80f68b110c8d1b4573a098f|3.89|2014-09-13 16:47:00|80.891462859624312|4|3800039125|99|35.645628106177277|0|45|74|-80.762919|9|35.442529|RTE CEREAL ALL FAMILY|1.95|1|KELLOGG RICE KRISPIES 9|5a19733e1f25571ceca2f85371f78e8ac927c20a|4.131077513560516|35.636605227883024|00038000318443|CEREAL|G1 GROCERY|-80.875654|80.875725547906455|471|1
35.585842|0ddbe0b642eb2ff949b47b387f7c3774a7d6b04b|2.18|2014-10-10 18:54:00|1.4102725052409182|4||99|0.6210901099944839|0|1|522|-80.875654|64|35.585842|FRESH TOMATOES|1.46|4|RED H/H TOMATOES, BULK|5a19733e1f25571ceca2f85371f78e8ac927c20a|4.131077513560516|0.61833652052202714|00204799000009|FRESH PRODUCE|PRODUCE|-80.875654|1.411546447003722|99|1
35.603432|15648004a2c223d5e2635aa094a8934ea5754480|6.49|2014-10-20 17:54:00|80.895431304315082|4|7703401130|274|35.810634030515281|0|10|141|-80.661096|21|35.172688|TRAIL MIXES AND BLENDS|0.0|1|SECOND NATURE WHLSOME MEDLEY|5b435b9eb052a62467d2e2d72f83b612a56ec667|14.317243366459325|35.810118468028598|00077034011302|NUTS|G1 GROCERY|-80.895009|80.89588013995828|474|1
35.603432|771e028ccbc8aa5b752462ff070401b3067c65fe|3.85|2015-02-08 16:19:00|80.895431304315082|4|4812127620|274|35.810634771696044|0|10|1037|-80.764523|164|35.341927|ENGLISH MUFFINS|0.0|7|THOMAS LITE MULTIGRAIN EM PP|5b435b9eb052a62467d2e2d72f83b612a56ec667|14.317243366459325|35.810118468028598|00048121276201|BREAKFAST|COMMERCIAL BAKERY|-80.895009|80.895550347478832|220|1
35.603432|4ff12f1ce7d70b3969cdccdeb17d15d8e9486457|1.72|2015-02-22 18:20:00|80.895431304315082|4||274|35.810634030515281|0|10|523|-80.661096|64|35.172688|FRESH POTATOES|0.35|4|COO SWEET POTATOES, BULK|5b435b9eb052a62467d2e2d72f83b612a56ec667|14.317243366459325|35.810118468028598|00204091000004|FRESH PRODUCE|PRODUCE|-80.895009|80.89588013995828|474|1
35.603432|af02bcfd5b82bebd7f23e6ff56bc52027a43c6c4|29.98|2015-01-14 20:03:00|80.895431304315082|4|75444108251|274|35.810634607837422|0|10|663|-80.737839|154|35.297134|FISH FILLETS/STEAKS PKGD|10.04|12|TILAPIA FILLETS|5b435b9eb052a62467d2e2d72f83b612a56ec667|14.317243366459325|35.810118468028598|00754441082513|FISH FILLETS/STEAKS|SEAFOOD|-80.895009|80.895638318215589|258|2
35.603432|e3f2c7d48ddbe4038c5f45be40b3102cfb18a243|2.99|2015-01-24 14:12:00|80.895431304315082|4|20443000000|274|35.810633469783859|0|10|510|-80.709466|64|35.124987|FRESH PINEAPPLE|0.0|4|GOLD PINEAPPLES|5b435b9eb052a62467d2e2d72f83b612a56ec667|14.317243366459325|35.810118468028598|00643126072003|FRESH PRODUCE|PRODUCE|-80.895009|80.896063182198972|157|1
35.603432|428f55129e96a5a367cffc524f209d8383b929e3|29.98|2014-12-07 09:23:00|80.895431304315082|4|75444108251|274|35.810634607837422|0|10|663|-80.737839|154|35.297134|FISH FILLETS/STEAKS PKGD|5.02|12|TILAPIA FILLETS|5b435b9eb052a62467d2e2d72f83b612a56ec667|14.317243366459325|35.810118468028598|00754441082513|FISH FILLETS/STEAKS|SEAFOOD|-80.895009|80.895638318215589|258|2
35.603432|ee55a907070f87d1a66f1e5401812edf5e498c81|1.89|2014-11-23 10:30:00|80.895431304315082|4|2000000065|274|35.810634030515281|0|10|1272|-80.661096|50|35.172688|BAG VEG STEAM|0.89|5|GG BOIL IN BAG ROSEMARY|5b435b9eb052a62467d2e2d72f83b612a56ec667|14.317243366459325|35.810118468028598|00020000481821|VEGETABLES-FROZEN|FROZEN|-80.895009|80.89588013995828|474|1
35.603432|19c0534564cbf79f94b270a9f1b91d628cb5ce3f|14.97|2014-10-05 11:48:00|80.895431304315082|4|20943300000|274|35.810634030515281|0|10|664|-80.661096|145|35.172688|SHRIMP WILD CAUGHT|4.3|12|WC P & D ARGENTINA PINK SHRMP|5b435b9eb052a62467d2e2d72f83b612a56ec667|14.317243366459325|35.810118468028598|00209433000001|SHRIMP|SEAFOOD|-80.895009|80.89588013995828|474|1
35.603432|944179fe6e61e8db4f317220618a421989b4d714|14.940000000000001|2014-11-09 15:26:00|80.895431304315082|4|20496100000|274|35.810632982565878|0|10|754|-80.64817|87|35.04711|NFS-SGLE STEM CUT FLOWER|0.0|9|*SINGLE STEM CUT FLOWERS|5b435b9eb052a62467d2e2d72f83b612a56ec667|14.317243366459325|35.810118468028598|00204961000004|FLORAL|FLORAL|-80.895009|80.896199593126511|129|6
35.603432|5df63fb6eeaea1e8112103c3d4455b5f39d755fa|13.99|2014-10-12 18:14:00|80.895431304315082|4|20943300000|274|35.810634030515281|0|10|664|-80.661096|145|35.172688|SHRIMP WILD CAUGHT|4.02|12|WC P & D ARGENTINA PINK SHRMP|5b435b9eb052a62467d2e2d72f83b612a56ec667|14.317243366459325|35.810118468028598|00209433000001|SHRIMP|SEAFOOD|-80.895009|80.89588013995828|474|1
35.603432|2c5955cebbf831df81f0a1034a20267eef0b11d9|28.26|2014-09-28 16:30:00|80.895431304315082|4|20943300000|274|35.810634030515281|0|10|664|-80.661096|145|35.172688|SHRIMP WILD CAUGHT|8.12|12|WC P & D ARGENTINA PINK SHRMP|5b435b9eb052a62467d2e2d72f83b612a56ec667|14.317243366459325|35.810118468028598|00209433000001|SHRIMP|SEAFOOD|-80.895009|80.89588013995828|474|1
35.603432|59e11b6ae55d92ea1d549eb27d76e82fd60bcf6e|14.86|2014-12-07 09:23:00|80.895431304315082|4|20889500000|274|35.810634607837422|0|10|648|-80.737839|154|35.297134|FISH FLTS/STK FARM RAISD|3.43|12|FR TILAPIA FILLET|5b435b9eb052a62467d2e2d72f83b612a56ec667|14.317243366459325|35.810118468028598|00208895000000|FISH FILLETS/STEAKS|SEAFOOD|-80.895009|80.895638318215589|258|1
35.603432|56788378767cca4a05a4dc2394dc20522a3ef48e|6.49|2014-11-20 19:39:00|80.895431304315082|4|3807520530|274|35.810634625013428|0|10|9983|-80.814133|889|35.333742|NFS-SPARKLING|0.0|13|VERDI RASPBERRY|5b435b9eb052a62467d2e2d72f83b612a56ec667|14.317243366459325|35.810118468028598|00038075205303|SPARKLING|WINE|-80.895009|80.895629682194382|472|1
35.603432|d1cb50ba3f81c6721ae8b43b89269065c7443a23|3.89|2015-01-29 19:09:00|80.895431304315082|4|2265530615|274|35.810634607837422|0|10|487|-80.737839|105|35.297134|PRECOOKED B/FAST SAUSAGE|0.92|19|BUTTERBALL COOKED TURK PATTIES|5b435b9eb052a62467d2e2d72f83b612a56ec667|14.317243366459325|35.810118468028598|00022655306160|BREAKFAST SAUSAGE|CASE READY MEATS|-80.895009|80.895638318215589|258|1
35.603432|4a6b7d14297972ebc6df5b9ab01d3feda333ee50|3.49|2014-11-04 17:34:00|80.895431304315082|4|7146426040|274|35.810634030515281|0|10|577|-80.661096|136|35.172688|OTHER MERCH FR MSC JUICE|0.0|4|BOLTHOUSE GREEN GOODNESS|5b435b9eb052a62467d2e2d72f83b612a56ec667|14.317243366459325|35.810118468028598|00071464240400|OTHER MERCHANDISE|PRODUCE|-80.895009|80.89588013995828|474|1
35.603432|92757035fe03615bf0f41b9ddedceb98c28909a4|3.79|2014-12-24 14:13:00|80.895431304315082|4|6414408004|274|35.810634030515281|0|10|60|-80.661096|9|35.172688|HOT CEREAL|0.0|1|WHEATENA HOT CEREAL|5b435b9eb052a62467d2e2d72f83b612a56ec667|14.317243366459325|35.810118468028598|00064144080045|CEREAL|G1 GROCERY|-80.895009|80.89588013995828|474|1
35.603432|1a6491987476fcb4e9f241a9e023d32641b220a9|4.99|2014-10-27 18:35:00|80.895431304315082|4|71575620002|274|35.810634030515281|0|10|504|-80.661096|64|35.172688|FRESH BERRIES|2.5|4|STRAWBERRIES 1LB CLAM|5b435b9eb052a62467d2e2d72f83b612a56ec667|14.317243366459325|35.810118468028598|00071430007525|FRESH PRODUCE|PRODUCE|-80.895009|80.89588013995828|474|1
35.23102|ce50502f861b976e68d467582e928de123410264|1.69|2014-10-08 18:55:00|1.4094857484078087|2|7680828073|205|0.6148972978359727|0|26|149|-80.8438|23|35.23102|WHSE PASTA CORE|0.31|1|BARILLA PASTA RIGATONI|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00076808502947|PASTA|G1 GROCERY|-80.8438|1.4109904898237917|205|1
35.23102|994a46969c486ff1dec68e0fdbf1044e88ad5355|3.19|2014-12-23 18:02:00|1.4094857484078087|2|7203655010|205|0.6148972978359727|0|26|317|-80.8438|52|35.23102|CHUNK AND BAR CHEESE|0.0|3|HT NY SHARP WHT CHEDDAR CHEESE|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00072036705082|CHEESE|DAIRY|-80.8438|1.4109904898237917|205|1
35.23102|db27c09de4a015b2659ecf03f82945fc7b5296b6|2.99|2015-02-14 17:56:00|80.843809562956082|2|7231000145|205|35.259238867051259|0|37|235|-80.810056|37|35.219587|GREEN TEA|0.49|1|BIGELOW TEA GREEN|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|35.255745041786184|00072310008472|TEA|G1 GROCERY|-80.8438|80.84380117605744|401|1
35.23102|588f1e5c8f466d55ba20ba565a32838d2d695b49|1.5|2014-10-29 17:43:00|80.843809562956082|2|7940038057|205|35.259238865964448|0|37|4121|-80.844274|1085|35.204336|DEODORANT|0.0|17|DOVE AP/DEO COOL ESSNTL TRAVEL|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|35.255745041786184|00079400380579|TRIAL SIZE|HBC|-80.8438|80.843809661522258|61|1
35.23102|c0d20ec25e548fe892106c9bf8d021956182b62f|2.19|2015-01-20 17:55:00|80.843809562956082|2|7418226090|205|35.259238865964448|0|37|722|-80.844274|73|35.204336|NFS-HAND SOAPS|1.19|1|SS HAND COUNTRY DESIGNS|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|35.255745041786184|00074182260125|PERSONAL SOAP/BATH ADDITIVES|G1 GROCERY|-80.8438|80.843809661522258|61|1
35.23102|f1b063fd6ae305f0e683dda954ff7a36a11e2fde|1.5|2014-11-13 18:16:00|80.843809562956082|2|7940038057|205|35.259238865964448|0|37|4121|-80.844274|1085|35.204336|DEODORANT|0.0|17|DOVE AP/DEO COOL ESSNTL TRAVEL|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|35.255745041786184|00079400380579|TRIAL SIZE|HBC|-80.8438|80.843809661522258|61|1
35.23102|a6ce347362b82d33dc21fdecef5c12531315dd95|1.5|2014-12-17 19:01:00|80.843809562956082|2|8680000015|205|35.259238867051259|0|37|4139|-80.810056|1085|35.219587|HAND & BODY LOTION|0.0|17|NEUTROGN HAND CRM TRIAL/TRAVEL|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|35.255745041786184|00086800000150|TRIAL SIZE|HBC|-80.8438|80.84380117605744|401|1
35.23102|945e0ad3c535579b6c3ec4904d13acc2d77b396a|3.99|2014-09-13 13:19:00|1.4094857484078087|2|4114305160|205|0.6148972978359727|0|26|119|-80.8438|17|35.23102|RAISINS|0.0|1|SUN MAID GOLDEN RAISINS|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00041143051603|FRUIT-DRIED|G1 GROCERY|-80.8438|1.4109904898237917|205|1
35.23102|0ec8237a8a803c7532b5911a1541be2f04061ecf|2.99|2015-02-25 16:33:00|80.843809562956082|2|3915310140|205|35.259238867051259|0|37|214|-80.810056|33|35.219587|BROTH|0.49|1|RACHAEL RAY CHCK LOW SOD STOCK|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|35.255745041786184|00039153101449|SOUP|G1 GROCERY|-80.8438|80.84380117605744|401|1
35.23102|b943e14e29ad45a10e589ebfc3a2cbcc03c120ad|2.29|2014-10-15 16:58:00|1.4094857484078087|2|4000040145|205|0.6148972978359727|0|26|62|-80.8438|7|35.23102|SPECIALTY BAR/BOX CHOCOLATE|0.0|1|DOVE MILK CHOC BAR|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00040000401452|CANDY|G1 GROCERY|-80.8438|1.4109904898237917|205|1
35.23102|75a8fa23e4261184e766ee4a1214253fe5ea8ed1|4.84|2014-09-30 19:13:00|1.4094857484078087|2|20596200000|205|0.6148972978359727|0|26|1821|-80.8438|410|35.23102|BH TURKEY|0.88|6|BOARS HEAD MAPLE HONEY TURKEY|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00205962000000|BH MEAT|DELI|-80.8438|1.4109904898237917|205|1
35.23102|1199a2647e109cf5d9611e35cd8997d9e078d569|3.63|2014-12-21 13:33:00|1.4094857484078087|2|20596200000|205|0.6148972978359727|0|26|1821|-80.8438|410|35.23102|BH TURKEY|0.0|6|BOARS HEAD MAPLE HONEY TURKEY|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00205962000000|BH MEAT|DELI|-80.8438|1.4109904898237917|205|1
35.23102|46c85958a6f9d38e6955337fc46295e8d1f9dd75|3.38|2015-01-01 14:26:00|1.4094857484078087|2|73801577715|205|0.6148972978359727|0|26|545|-80.8438|64|35.23102|FRESH SPROUTS|0.38|4|BLACK-EYED PEAS, PKG|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00738015777159|FRESH PRODUCE|PRODUCE|-80.8438|1.4109904898237917|205|2
35.23102|f5f7821e1c2a6df14058bae4781c459874f7389f|3.14|2014-12-20 17:18:00|80.843809562956082|2||205|35.259238865880455|0|37|500|-80.826724|64|35.195689|FRESH APPLES|0.53|4|HONEY CRISP APPLE|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|35.255745041786184|00233283000003|FRESH PRODUCE|PRODUCE|-80.8438|80.843810022625746|412|1
35.23102|ad2677efd60590eb3251965ddf0165e8078f4075|1.04|2015-03-09 18:55:00|1.4094857484078087|2||205|0.6148972978359727|0|26|523|-80.8438|64|35.23102|FRESH POTATOES|0.0|4|COO RUSSET POTATOES, BULK|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00204072000009|FRESH PRODUCE|PRODUCE|-80.8438|1.4109904898237917|205|1
35.23102|75b7271ee0bac5d707589f4a03376cfe997e2c19|1.9|2014-12-14 17:23:00|80.843809562956082|2|61300871771|205|35.259238865964448|0|37|99|-80.844274|32|35.204336|LIQUID TEA|0.0|1|ARIZONA ARNOLD PALMER HALF/HAL|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|35.255745041786184|00613008719302|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.8438|80.843809661522258|61|2
35.23102|477e14da8d90065ca28558f74fddec220bf7bd62|1.9|2014-12-30 15:09:00|1.4094857484078087|2|61300871771|205|0.6148972978359727|0|26|99|-80.8438|32|35.23102|LIQUID TEA|0.15|1|ARIZONA ARNOLD PALMER HALF/HAL|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00613008719302|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.8438|1.4109904898237917|205|2
35.23102|ba13e80f4ab854652a01e4d5e56a85bafc4dfe7d|2.19|2015-02-15 15:10:00|80.843809562956082|2|64420931131|205|35.259238865964448|0|37|8|-80.844274|2|35.204336|BROWNIE MIXES|0.94|1|D HINES DARK CHOC FUDGE BRWNIE|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|35.255745041786184|00644209420957|BAKING MIXES|G1 GROCERY|-80.8438|80.843809661522258|61|1
35.23102|7dc223880f2bf4ba88fb9257a6d81835236d27a9|0.95|2014-10-04 19:12:00|80.843809562956082|2|61300871771|205|35.259238863556888|0|37|99|-80.945176|32|35.323246|LIQUID TEA|0.0|1|ARIZONA ARNOLD PALMER HALF/HAL|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|35.255745041786184|00613008719302|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.8438|80.843817235540442|166|1
35.23102|998bf4c68da513a9c4d2ebf9418781bdabc6d1a1|1.9|2014-10-02 18:00:00|80.843809562956082|2|61300871771|205|35.259238867051259|0|37|99|-80.810056|32|35.219587|LIQUID TEA|0.0|1|ARIZONA ARNOLD PALMER HALF/HAL|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|35.255745041786184|00613008719302|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.8438|80.84380117605744|401|2
35.23102|2881212eb281f547209559edb66408f30333fe87|0.97|2015-02-23 16:42:00|80.843809562956082|2|7203637031|205|35.259238867051259|0|37|212|-80.810056|33|35.219587|CONDENSED SOUP|0.0|1|HT SP HLTHY CRM MUSHROOM|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|35.255745041786184|00072036370389|SOUP|G1 GROCERY|-80.8438|80.84380117605744|401|1
35.23102|c14c71dcce4240c3aea2a0d63ea6629602c62170|5.99|2015-01-23 17:18:00|1.4094857484078087|2|76108880157|205|0.6148972978359727|0|26|1939|-80.8438|465|35.23102|COLD PREP FOODS SIDES|0.0|6|YUKON GOLD MASHED POTATOES|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00761088801575|COLD PREPARED FOODS|DELI|-80.8438|1.4109904898237917|205|1
35.23102|b8f71553408b75682529aa6eb989b952c33a2da1|2.59|2014-11-19 17:42:00|1.4094857484078087|2|7203695296|205|0.6148972978359727|0|26|1654|-80.8438|381|35.23102|DESSERT CAKES|0.0|14|RED VELVET CAKE SLICE|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00072036952967|CAKES|BAKERY|-80.8438|1.4109904898237917|205|1
35.23102|b41ddeb8ed2e1e0d5704e89a583b0565d7f5e419|3.29|2014-09-16 15:15:00|1.4094857484078087|2|7203698583|205|0.6148972978359727|0|26|67|-80.8438|10|35.23102|SOLUBLE INSTANT|0.0|1|HT DECAF INSTANT COFFEE|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00072036985835|COFFEE|G1 GROCERY|-80.8438|1.4109904898237917|205|1
35.23102|e788380364b48dd7a1363fb25325ad1d1fac236a|3.89|2015-02-01 16:36:00|1.4094857484078087|2|8411410812|205|0.6148972978359727|0|26|201|-80.8438|31|35.23102|POTATO CHIPS|0.0|1|KETTLE LIGHT CHIPS|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00084114108128|SNACKS|G1 GROCERY|-80.8438|1.4109904898237917|205|1
35.23102|f8a79a1453d3ca8e412c0c95c19d90dbb938d056|1.19|2015-01-15 18:06:00|1.4094857484078087|2|3940001747|205|0.6148972978359727|0|26|242|-80.8438|39|35.23102|CANNED BEANS|0.19|1|BUSH BEAN KIDNEY DK|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00039400017349|VEGETABLES-CAN/JAR|G1 GROCERY|-80.8438|1.4109904898237917|205|1
35.23102|c03448909f862c3d9f827ad294db4a986d504541|1.19|2014-10-22 18:24:00|1.4094857484078087|2|3940001747|205|0.6148972978359727|0|26|242|-80.8438|39|35.23102|CANNED BEANS|0.19|1|BUSH BEAN KIDNEY DK|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00039400017349|VEGETABLES-CAN/JAR|G1 GROCERY|-80.8438|1.4109904898237917|205|1
35.23102|40bf8e1ad23e2a500152fd6833a7b7cbf0097ef5|2.39|2014-10-13 17:02:00|1.4094857484078087|2|4127102562|205|0.6148972978359727|0|26|341|-80.8438|57|35.23102|CREAMERS|0.0|3|ITNAT'L DELIGHT FRNCH VANILLA|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00041271025620|MILK|DAIRY|-80.8438|1.4109904898237917|205|1
35.23102|fb4bb061f3b87c3038fd05f260209f4ddc57c7da|2.39|2014-11-08 17:57:00|1.4094857484078087|2|4127102562|205|0.6148972978359727|0|26|341|-80.8438|57|35.23102|CREAMERS|0.0|3|ITNAT'L DELIGHT FRNCH VANILLA|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00041271025620|MILK|DAIRY|-80.8438|1.4109904898237917|205|1
35.23102|683a858b6ef512d089401db396f008869a98cbae|8.39|2014-12-02 15:47:00|1.4094857484078087|2|20899300000|205|0.6148972978359727|0|26|1419|-80.8438|201|35.23102|SMART CHICKEN ORGANIC|0.0|2|SMART ORGANIC BNLS CHICK BRST|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00208993000001|POULTRY|MEAT|-80.8438|1.4109904898237917|205|1
35.23102|51687996871745888d8196e62b84a9e25bbe3c7d|5.95|2014-09-11 18:17:00|1.4094857484078087|2|20689900000|205|0.6148972978359727|0|26|2027|-80.8438|510|35.23102|SOMETHING CLASSIC|0.0|6|SOMETHING CLASSIC SANDWICHES|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00206899000002|SOMETHING CLASSIC|DELI|-80.8438|1.4109904898237917|205|1
35.23102|fbb858f58f2a8f952062c06711fa8419da109cad|0.96|2015-01-17 16:32:00|80.843809562956082|2||205|35.259238865880455|0|37|524|-80.826724|64|35.195689|FRESH PROD FRESH ONIONS|0.0|4|COO SHALLOTS, BULK|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|35.255745041786184|00204662000006|FRESH PRODUCE|PRODUCE|-80.8438|80.843810022625746|412|1
35.23102|5d9fb9980ddb3fc3ba95e72ed2ba9e4f7f75daa0|3.99|2014-10-31 17:29:00|80.843809562956082|2|4000015140|205|35.259238865964448|0|37|46|-80.844274|7|35.204336|PKG CHOC|0.99|1|3 MUSKETEER FUN SIZE|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|35.255745041786184|00040000151227|CANDY|G1 GROCERY|-80.8438|80.843809661522258|61|1
35.23102|ee04a4f2d3d4ace3ed0dc2ff9a3784c3ec4f79a4|3.99|2015-01-04 19:02:00|1.4094857484078087|2|7203695283|205|0.6148972978359727|0|26|1663|-80.8438|381|35.23102|CREME CAKE|0.0|14|FFM SLICED POUND CAKE|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00072036952752|CAKES|BAKERY|-80.8438|1.4109904898237917|205|1
35.23102|e96ae0bd7a4d9997c85e43fea86ed4d2325317c3|5.38|2014-09-28 17:10:00|80.843809562956082|2|5000032822|205|35.259238867051259|0|37|341|-80.810056|57|35.219587|CREAMERS|0.0|3|COFFEE-MATE HAZLENUT|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|35.255745041786184|00050000328222|MILK|DAIRY|-80.8438|80.84380117605744|401|2
35.23102|b9725034c9d23c12b2bf3b945983bfa07feb8e48|3.0|2015-02-08 13:40:00|1.4094857484078087|2|61300873089|205|0.6148972978359727|0|26|99|-80.8438|32|35.23102|LIQUID TEA|0.0|1|PP ARIZONA ARNOLD PALMER|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00613008730895|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.8438|1.4109904898237917|205|3
35.23102|788998df8d3d0865bc25999028bdca44c4d689a0|6.0|2015-03-03 18:28:00|80.843809562956082|2|89470001004|205|35.259238867051259|0|37|685|-80.810056|61|35.219587|GREEK|0.0|3|CHOBANI SEASONAL GREEN TEA|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|35.255745041786184|00818290013866|YOGURT|DAIRY|-80.8438|80.84380117605744|401|5
35.23102|79fae890aa0cf87974ad45440be387773cfd1020|3.99|2014-12-01 11:55:00|1.4094857484078087|2|3120000455|205|0.6148972978359727|0|26|130|-80.8438|20|35.23102|CRANBERRY JUICE/DRINKS-SHELF|0.0|1|OS SPARKLING CRANBERY DIET 4PK|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00031200003461|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.8438|1.4109904898237917|205|1
35.23102|d2400d692f93347ca81159dee8bae06b6639b7b9|5.49|2015-01-30 16:57:00|1.4094857484078087|2|7203695136|205|0.6148972978359727|0|26|1687|-80.8438|385|35.23102|THAW & SELL (SWEET GOODS)|0.0|14|FUDGE ICED BROWNIE|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00072036951359|SWEET GOODS|BAKERY|-80.8438|1.4109904898237917|205|1
35.23102|cda5234821054f4c038c09068b60d584c33d267e|1.99|2014-10-09 16:13:00|1.4094857484078087|2|4430005462|205|0.6148972978359727|0|26|247|-80.8438|39|35.23102|VEGETABLES-FLANKER|0.0|1|AUNT NELLIE BEETS ONION PICKL|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00044300054684|VEGETABLES-CAN/JAR|G1 GROCERY|-80.8438|1.4109904898237917|205|1
35.23102|2ab550ee2d6507a387d00f6d0b7bd54f3f1235d5|2.19|2014-09-20 17:39:00|80.843809562956082|2||205|35.259238865880455|0|37|536|-80.826724|64|35.195689|FRESH SQUASH|0.0|4|COO ZUCCHINI SQUASH, FANCY|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|35.255745041786184|00204067000007|FRESH PRODUCE|PRODUCE|-80.8438|80.843810022625746|412|1
35.23102|e3c771ba898fab7b8135146fd35bbfe57ea8ae24|5.63|2014-10-20 10:45:00|1.4094857484078087|2|27082900000|205|0.6148972978359727|0|26|973|-80.8438|201|35.23102|FRESH PERDUE CHICKEN|0.0|2|PERDUE BNLS CHICKEN BREAST|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00270829000004|POULTRY|MEAT|-80.8438|1.4109904898237917|205|1
35.23102|d2ab168fdded54d8bad4f9e174f99981cf74e29b|0.99|2014-10-02 18:04:00|80.843809562956082|2|4000000435|205|35.259238867051259|0|37|47|-80.810056|7|35.219587|REGISTER BARS|0.0|1|(FE)DOVE MILK CHOC SINGLES|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|35.255745041786184|00040000459842|CANDY|G1 GROCERY|-80.8438|80.84380117605744|401|1
35.23102|d3b51a83613b804b050649b794e13be27ea6f6f9|2.59|2014-12-10 16:50:00|1.4094857484078087|2|7203695278|205|0.6148972978359727|0|26|1654|-80.8438|381|35.23102|DESSERT CAKES|0.0|14|DOUBLE FUDGE CAKE SLICE|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00072036952783|CAKES|BAKERY|-80.8438|1.4109904898237917|205|1
35.23102|45bdbd29f72f70dc56494861fe1dd53e80b6b8b0|12.78|2014-10-20 10:50:00|1.4094857484078087|2|4154800385|205|0.6148972978359727|0|26|252|-80.8438|45|35.23102|PREMIUM ICE CREAM|3.2|5|EDY'S SLOW CHURNED FRENCH VA|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|0.61471665291522548|00041548737867|ICE CREAM|FROZEN|-80.8438|1.4109904898237917|205|2
35.23102|9990aecafaba4bd88342388e261df215a0554bf8|1.89|2014-10-31 17:20:00|80.843809562956082|2|2000000065|205|35.259238865964448|0|37|1275|-80.844274|50|35.204336|BOX VEG|0.0|5|GG HONEY GLAZED CARROTS|5c60b0621d4a13fc5ba9772d3afe836b40777918|1.9498555682467458|35.255745041786184|00020000125688|VEGETABLES-FROZEN|FROZEN|-80.8438|80.843809661522258|61|1
35.059823|4a060cd58331fa50ce22d1693dc09339d838c6a0|2.99|2014-11-27 01:11:00|1.4091206135396188|4|7203698444|66|0.6119093465164359|0|47|266|-80.816172|307|35.059823|SHELLS AND PIE CRUSTS|0.99|5|HT PIE CRUSTS DEEP DISH|5cb11b1d487f6f06fe4089321738c2ce39450bb1|0.6144447802952047|0.61242566243833529|00072036984449|DESSERTS FROZEN|FROZEN|-80.816172|1.4105082902580508|66|1
35.059823|14e026243cbafa945f296c2cf96123e2daa267c2|14.89|2015-01-26 22:39:00|80.816179662140996|4|36761830050|66|35.06871542027168|0|41|4502|-80.848528|1210|35.053394|LAXATIVE-STIMULANT|2.0|17|JHK) SENOKOT TABLETS|5cb11b1d487f6f06fe4089321738c2ce39450bb1|0.6144447802952047|35.070508771677183|00367618300503|STOMACH REMEDIES|HBC|-80.816172|80.816174314867041|11|1
35.059823|4663a707484fb9f43442ea225b0b68f7fd0bfd9c|4.79|2014-11-17 21:46:00|1.4091206135396188|4|18685200031|66|0.6119093465164359|0|47|275|-80.816172|45|35.059823|SUPER PREMIUM ICE CREAM|0.0|5|TALENTI CARIBB COCONUT GELATO|5cb11b1d487f6f06fe4089321738c2ce39450bb1|0.6144447802952047|0.61242566243833529|00186852000327|ICE CREAM|FROZEN|-80.816172|1.4105082902580508|66|1
35.059823|989ff2e8e717bee5ef58e17a1b8e28374dc4bc25|13.99|2014-11-27 11:58:00|1.4091206135396188|4|7289010016|66|0.6119093465164359|0|47|459|-80.816172|83|35.059823|IMPORT BEER|0.0|16|AMSTEL LIGHT 12PK 12OZ BOTTLES|5cb11b1d487f6f06fe4089321738c2ce39450bb1|0.6144447802952047|0.61242566243833529|00072890100160|IMPORT BEER|BEER|-80.816172|1.4105082902580508|66|1
35.059823|21d2f06e57df81133201f98ce6f4960b0622771b|5.36|2015-02-01 16:27:00|1.4091206135396188|4||66|0.6119093465164359|0|47|566|-80.816172|64|35.059823|SERVICE BAR|0.37|4|HT 7 LAYER MEXICAN BEAN DIP|5cb11b1d487f6f06fe4089321738c2ce39450bb1|0.6144447802952047|0.61242566243833529|00204506000001|FRESH PRODUCE|PRODUCE|-80.816172|1.4105082902580508|66|1
35.059823|5114c6de62a2050301b199b20790f81071e98732|1.29|2014-11-26 00:26:00|80.816179662140996|4||66|35.068715419239624|0|41|527|-80.78468|64|35.096737|FRESH CARROTS|0.0|4|COO CARROTS, BUNCHED|5cb11b1d487f6f06fe4089321738c2ce39450bb1|0.6144447802952047|35.070508771677183|00204094000001|FRESH PRODUCE|PRODUCE|-80.816172|80.816177723293578|30|1
35.059823|4f77be1c9c256fb5985ee9381248a838b8b57712|6.0|2015-03-07 19:51:00|1.4091206135396188|4|2400001738|66|0.6119093465164359|0|47|257|-80.816172|39|35.059823|TOMATOES|0.2|1|DEL MONTE TOMATO STEWD ITALIAN|5cb11b1d487f6f06fe4089321738c2ce39450bb1|0.6144447802952047|0.61242566243833529|00024000019381|VEGETABLES-CAN/JAR|G1 GROCERY|-80.816172|1.4105082902580508|66|5
35.059823|404a4959b1d48930b93ea66b02fad633ce58d725|3.75|2015-03-03 21:35:00|80.816179662140996|4|4138309010|66|35.068715419239624|0|41|1263|-80.78468|57|35.096737|GOOD FOR YOU MILK|0.0|3|LACTAID 100 REDUCED FAT MILK|5cb11b1d487f6f06fe4089321738c2ce39450bb1|0.6144447802952047|35.070508771677183|00041383090103|MILK|DAIRY|-80.816172|80.816177723293578|30|1
35.059823|33bab94c8e692e236db503dacced81181399acbe|8.99|2014-09-21 15:45:00|1.4091206135396188|4|18195400002|66|0.6119093465164359|0|47|459|-80.816172|83|35.059823|IMPORT BEER|0.0|16|PERONI 6PK LNNR|5cb11b1d487f6f06fe4089321738c2ce39450bb1|0.6144447802952047|0.61242566243833529|00181954000022|IMPORT BEER|BEER|-80.816172|1.4105082902580508|66|1
35.059823|d5af32e15d231cd472637ba77c4a4091b9bc201b|2.58|2015-01-20 14:55:00|1.4091206135396188|4|2700039014|66|0.6119093465164359|0|47|257|-80.816172|39|35.059823|TOMATOES|0.0|1|HUNTS TOMATO SAUCE 15|5cb11b1d487f6f06fe4089321738c2ce39450bb1|0.6144447802952047|0.61242566243833529|00027000390146|VEGETABLES-CAN/JAR|G1 GROCERY|-80.816172|1.4105082902580508|66|2
35.059823|756a9bb0473eae7036d3971cf12373802145b8de|4.39|2014-10-20 09:52:00|1.4091206135396188|4|1313006025|66|0.6119093465164359|0|47|60|-80.816172|9|35.059823|HOT CEREAL|0.0|1|CREAM OF WHEAT INST ORIGINAL|5cb11b1d487f6f06fe4089321738c2ce39450bb1|0.6144447802952047|0.61242566243833529|00013130060257|CEREAL|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|a53e7cf82e5245a372cadb8da49eae5ffac97299|34.99|2015-02-14 16:04:00|1.4091206135396188|4|7203696867|66|0.6119093465164359|0|47|740|-80.816172|87|35.059823|NFS-ROSE BQT|5.0|9|PREMIUM DZ ROSE BOUQUET|5cb11b1d487f6f06fe4089321738c2ce39450bb1|0.6144447802952047|0.61242566243833529|00072036968678|FLORAL|FLORAL|-80.816172|1.4105082902580508|66|1
35.172688|14516e6238a5c6c2eff7fca8483347ad8cb7ab39|2.85|2015-02-23 14:16:00|1.4094857484078087|4|7203604237|474|0.6138792123766993|0|26|41|-80.661096|6|35.172688|BREAKFAST BARS|0.88|1|HT BAR CEREAL APPLE LF|5cea8d928d67ff4fedaff56216d5691b730c0a8b|4.150707219205793|0.61471665291522548|00072036042385|BREAKFAST FOODS|G1 GROCERY|-80.661096|1.407801703467228|474|1
35.172688|5d37cffef865102b0e2b59cfd7e7ece302607d11|3.34|2014-09-29 13:47:00|1.4094857484078087|4|7203643010|474|0.6138792123766993|0|26|252|-80.661096|45|35.172688|PREMIUM ICE CREAM|0.84|5|HT PREM CHOCOLATE IC|5cea8d928d67ff4fedaff56216d5691b730c0a8b|4.150707219205793|0.61471665291522548|00072036430113|ICE CREAM|FROZEN|-80.661096|1.407801703467228|474|1
35.172688|5068261fd653810bd3269aa25838f4a5b9a9e3c4|4.99|2014-09-12 16:55:00|1.4094857484078087|4|2840015297|474|0.6138792123766993|0|26|204|-80.661096|31|35.172688|TORTILLA CHIPS|1.0|1|DORITOS NACHO CHEES PARTY SIZE|5cea8d928d67ff4fedaff56216d5691b730c0a8b|4.150707219205793|0.61471665291522548|00028400152976|SNACKS|G1 GROCERY|-80.661096|1.407801703467228|474|1
35.172688|d386acd18719ba9b4452536e0098ef86b62744bd|1.9|2014-12-20 16:39:00|1.4094857484078087|4|4600028869|474|0.6138792123766993|0|26|77|-80.661096|272|35.172688|HISP SAUCES/SEASONINGS|0.0|1|E  OEP SEASONING TACO|5cea8d928d67ff4fedaff56216d5691b730c0a8b|4.150707219205793|0.61471665291522548|00046000288697|HISPANIC PREP. FOODS|G1 GROCERY|-80.661096|1.407801703467228|474|2
35.172688|a7db16bbf4c61f62d2659bcbe202adbd8e1b2721|1.99|2015-02-19 14:03:00|1.4094857484078087|4|7127915102|474|0.6138792123766993|0|26|555|-80.661096|64|35.172688|PACKAGED SALADS|0.0|4|F.E. GREEN LEAF SHREDS|5cea8d928d67ff4fedaff56216d5691b730c0a8b|4.150707219205793|0.61471665291522548|00071279151021|FRESH PRODUCE|PRODUCE|-80.661096|1.407801703467228|474|1
35.172688|85e6171bdbe013b3c2b0bac079291ff570e6b07f|1.5|2015-01-27 14:14:00|1.4094857484078087|4|7203663107|474|0.6138792123766993|0|26|1262|-80.661096|57|35.172688|HALF N HALF WHIPPING CREAM|0.0|3|HT HALF & HALF|5cea8d928d67ff4fedaff56216d5691b730c0a8b|4.150707219205793|0.61471665291522548|00072036632036|MILK|DAIRY|-80.661096|1.407801703467228|474|1
35.172688|a67000790ed94da0f48acb020d83848528eaedfd|8.99|2014-12-04 12:45:00|80.632521683083056|4|7017786268|474|35.232758219847241|0|39|1247|-80.70901|37|35.17335|SINGLES PODS CUPS TEA|2.0|1|I/O TWININGS K CUP CHRISTMAS|5cea8d928d67ff4fedaff56216d5691b730c0a8b|4.150707219205793|35.177497916598789|00070177862688|TEA|G1 GROCERY|-80.661096|80.661111490811336|174|1
35.43259|e51d3c19f92a937c6ca3976f89e48ce7782ed1d7|2.69|2014-09-13 18:12:00|1.4057311447477159|4|7225001739|202|0.6184153580092175|0|52|1025|-80.605588|162|35.43259|WHITE|0.0|7|NATOWN WHITEWHEAT RTOP BRD|5e72859ad4956d2afd344ad160f7c661d4d97781|6.875442647461331|0.6209993146566879|00072250017398|SLICED BREAD|COMMERCIAL BAKERY|-80.605588|1.406832906106031|202|1
35.297134|274da622a3f1bcf7ab90c4be223a37e493536251|11.54|2015-03-04 20:18:00|80.728244613218536|4|7203698516|258|35.309302352083094|0|5|426|-80.814133|72|35.333742|NFS-PAPER TOWELS|0.0|1|YH TOWEL 8RL PRINT|5f379bb125b099a8ddd709053c34c5f11eafa577|0.8408037439038158|35.296297200616316|00072036985163|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.737839|80.737839504004725|472|2
35.297134|d3c89001731ba9a68f125a3ef266273ad9dd73da|2.29|2014-09-21 01:13:00|80.728244613218536|4|7203636049|258|35.309302352083975|0|5|30|-80.780702|4|35.318911|CARBONATED WATER|0.62|1|HT SIMPLY WHT GRAPE 4 PK|5f379bb125b099a8ddd709053c34c5f11eafa577|0.8408037439038158|35.296297200616316|00072036360489|BOTTLED WATER|G1 GROCERY|-80.737839|80.737839470807501|167|1
35.297134|624e30999aadb67a5eb4aee6d9ab4d61225ebc44|3.39|2014-12-06 13:06:00|80.728244613218536|4|7203620985|258|35.309302351368686|0|5|130|-80.764523|20|35.341927|CRANBERRY JUICE/DRINKS-SHELF|0.39|1|HT CRANBERRY CHERRY COCKTAIL|5f379bb125b099a8ddd709053c34c5f11eafa577|0.8408037439038158|35.296297200616316|00072036200945|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.737839|80.737844134036735|220|1
35.297134|a4be33e8723a1992667a2e145ee09d37cc7c6684|3.49|2015-01-27 19:05:00|80.728244613218536|4|2265530605|258|35.309302351368686|0|5|357|-80.764523|104|35.341927|SMOKED SAUSAGE ROPES|0.99|19|BBALL HOT & SPICY SMKD SAUSAGE|5f379bb125b099a8ddd709053c34c5f11eafa577|0.8408037439038158|35.296297200616316|00022655306139|DINNER SAUSAGE|CASE READY MEATS|-80.737839|80.737844134036735|220|1
35.297134|7cc8e09a086975362490674bef61a288676b27d3|3.89|2014-10-03 18:00:00|80.728244613218536|4|7261345171|258|35.309302352083094|0|5|417|-80.814133|71|35.333742|NFS-FABRIC SOFTENERS|0.89|1|SNUGGLE LIQ FAB SOFT PUR FUSIO|5f379bb125b099a8ddd709053c34c5f11eafa577|0.8408037439038158|35.296297200616316|00072613451746|LAUNDRY SUPPLIES|G1 GROCERY|-80.737839|80.737839504004725|472|1
35.297134|2e958093edcb4f83c17afcf82b41937d70787617|2.99|2014-09-13 10:15:00|80.728244613218536|4|7203655010|258|35.309302352083094|0|5|317|-80.814133|52|35.333742|CHUNK AND BAR CHEESE|0.0|3|HT EXTRA SHARP CHEDDAR CHEESE|5f379bb125b099a8ddd709053c34c5f11eafa577|0.8408037439038158|35.296297200616316|00072036559951|CHEESE|DAIRY|-80.737839|80.737839504004725|472|1
35.297134|be0339435655c6b492bcadb5d09256bbf4b57429|5.0|2014-10-16 12:51:00|80.728244613218536|4|20491700000|258|35.309302291131971|0|5|562|-80.992182|64|35.103409|FRESH CUT FRUIT|0.0|4|POM/BLUEBERRY (IN-STORE)|5f379bb125b099a8ddd709053c34c5f11eafa577|0.8408037439038158|35.296297200616316|00204917000003|FRESH PRODUCE|PRODUCE|-80.737839|80.73788619541844|88|1
35.297134|8d5bcad12c7713688947e6b2a57ee4fefae77bfe|3.99|2014-09-30 21:22:00|80.728244613218536|4|7684010015|258|35.309302352083094|0|5|275|-80.814133|45|35.333742|SUPER PREMIUM ICE CREAM|0.0|5|BEN & JERRY KARMEL SUTRA|5f379bb125b099a8ddd709053c34c5f11eafa577|0.8408037439038158|35.296297200616316|00076840101542|ICE CREAM|FROZEN|-80.737839|80.737839504004725|472|1
35.297134|9ce7d43c3273e991ea346465b47e08e16b0ad848|13.47|2014-12-24 18:58:00|80.728244613218536|4|76352830903|258|35.309302352083975|0|5|339|-80.780702|57|35.318911|EGGNOGS/DRINKS|0.5|3|I/O PROMISE LAND EGG NOG|5f379bb125b099a8ddd709053c34c5f11eafa577|0.8408037439038158|35.296297200616316|00763528309030|MILK|DAIRY|-80.737839|80.737839470807501|167|3
35.323246|56ee10b794811ef9a4a051eb7c6c14e61f5cad11|8.58|2014-10-04 13:31:00|1.4102725052409182|4|2840016014|166|0.6165069451919168|0|1|201|-80.945176|31|35.323246|POTATO CHIPS|2.15|1|LAYS CLASSIC|5f7d00aa6518e90eb42a5b17beba6616f838ff9c|2.060807865397842|0.61833652052202714|00028400160148|SNACKS|G1 GROCERY|-80.945176|1.4127598348062935|166|2
35.323246|ea7e1aba5bc2b82ec54173ee6ba6739766072ac8|8.58|2014-11-22 20:05:00|1.4102725052409182|4|2840016014|166|0.6165069451919168|0|1|201|-80.945176|31|35.323246|POTATO CHIPS|2.14|1|LAYS CLASSIC|5f7d00aa6518e90eb42a5b17beba6616f838ff9c|2.060807865397842|0.61833652052202714|00028400160148|SNACKS|G1 GROCERY|-80.945176|1.4127598348062935|166|2
35.323246|2a255011739427fb3021759af4bab807d0a2bcf8|13.49|2014-09-13 18:31:00|1.4102725052409182|4|36382455020|166|0.6165069451919168|0|1|4236|-80.945176|1200|35.323246|DEX ADULT/CHILDREN|0.0|17|MUCINEX FSTMX ADLT NTTME CAPLT|5f7d00aa6518e90eb42a5b17beba6616f838ff9c|2.060807865397842|0.61833652052202714|00363824550206|COUGH/COLD/SINUS|HBC|-80.945176|1.4127598348062935|166|1
35.219587|a66125773d4436d3c04cf45e2cf725f75610ae15|3.99|2014-10-26 13:15:00|1.4094857484078087|4|7203663995|401|0.6146977543425921|0|26|342|-80.810056|57|35.219587|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|5f7f00198fe8c1d13c009c301012d7d18b9584e9|3.119268612967971|0.61471665291522548|00072036631282|MILK|DAIRY|-80.810056|1.4104015459209989|401|1
35.219587|4b38fe2854e7332f1317b40988cacca437b0311b|8.45|2014-10-26 13:14:00|1.4094857484078087|4|7680828073|401|0.6146977543425921|0|26|149|-80.810056|23|35.219587|WHSE PASTA CORE|0.0|1|BARILLA PASTA PENNE RIGATE|5f7f00198fe8c1d13c009c301012d7d18b9584e9|3.119268612967971|0.61471665291522548|00076808280739|PASTA|G1 GROCERY|-80.810056|1.4104015459209989|401|5
35.219587|d94bc5e7948caffa74299dcdf225e3a6f3a3247f|1.89|2014-10-27 19:10:00|80.810069425230125|4|4000000432|401|35.264729917825605|0|23|47|-80.737839|7|35.297134|REGISTER BARS|0.0|1|E  SNICKERS KING SIZE BAR|5f7f00198fe8c1d13c009c301012d7d18b9584e9|3.119268612967971|35.240679762029046|00040000002635|CANDY|G1 GROCERY|-80.810056|80.810118708832604|258|1
35.219587|5ecdc981afadfb4994005a59e214a24200a8a5f0|1.89|2014-10-27 19:09:00|80.810069425230125|4|4000000432|401|35.264729917825605|0|23|47|-80.737839|7|35.297134|REGISTER BARS|0.0|1|E  SNICKERS KING SIZE BAR|5f7f00198fe8c1d13c009c301012d7d18b9584e9|3.119268612967971|35.240679762029046|00040000002635|CANDY|G1 GROCERY|-80.810056|80.810118708832604|258|1
34.977331|883ceb474eafda1905a4a5699e0936397df5e7fe|4.29|2014-10-20 13:03:00|1.41290891556208|2|2840016014|149|0.6104695895098807|0|33|201|-81.027334|31|34.977331|POTATO CHIPS|1.29|1|LAYS WAVY REGULAR|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00028400160209|SNACKS|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|5f1180b2d1ea7adacfe8473bda0979be873fe78b|17.97|2014-12-09 14:11:00|1.41290891556208|2|1834175105|149|0.6104695895098807|0|33|9934|-81.027334|885|34.977331|NFS POP CHARDONNAY|0.0|13|CB-BAREFOOT CHARDONNAY|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00018341751055|POPULAR (4-$7.99)|WINE|-81.027334|1.4141937624131469|149|3
34.977331|98ef767343a2c2928d174d38bd0c04437367524f|11.98|2014-10-10 10:26:00|1.41290891556208|2|1834175105|149|0.6104695895098807|0|33|9934|-81.027334|885|34.977331|NFS POP CHARDONNAY|2.02|13|CB-BAREFOOT CHARDONNAY|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00018341751055|POPULAR (4-$7.99)|WINE|-81.027334|1.4141937624131469|149|2
34.977331|d5c966e1c95d0042cbd2fe1cd157f1e3f3fe403b|4.29|2014-12-24 10:12:00|1.41290891556208|2|2840016014|149|0.6104695895098807|0|33|201|-81.027334|31|34.977331|POTATO CHIPS|2.15|1|LAYS WAVY REGULAR|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00028400160209|SNACKS|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|5ba8dc70304783638b450b05eae469c828df6ce0|9.0|2014-12-10 13:50:00|1.41290891556208|2|1834175105|149|0.6104695895098807|0|33|9934|-81.027334|885|34.977331|NFS POP CHARDONNAY|0.0|13|CB-BAREFOOT CHARDONNAY|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00018341751055|POPULAR (4-$7.99)|WINE|-81.027334|1.4141937624131469|149|2
34.977331|df77179d0a4db4c5bd473bacc33847758de4c9aa|15.0|2015-02-05 10:08:00|1.41290891556208|2|1834175105|149|0.6104695895098807|0|33|9934|-81.027334|885|34.977331|NFS POP CHARDONNAY|0.0|13|CB-BAREFOOT CHARDONNAY|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00018341751055|POPULAR (4-$7.99)|WINE|-81.027334|1.4141937624131469|149|3
34.977331|24a957a26e7e1f66529ffc8fb6d7628b8a3fd0ba|9.0|2014-12-26 15:59:00|1.41290891556208|2|1834175105|149|0.6104695895098807|0|33|9934|-81.027334|885|34.977331|NFS POP CHARDONNAY|0.0|13|CB-BAREFOOT CHARDONNAY|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00018341751055|POPULAR (4-$7.99)|WINE|-81.027334|1.4141937624131469|149|2
34.977331|dc1102d819e9a58e2672ff421fd475e768056d61|2.38|2014-10-27 15:34:00|1.41290891556208|2|20895000000|149|0.6104695895098807|0|33|977|-81.027334|201|34.977331|FRESH HT CHICKEN|0.0|2|HT FRESH CHICKEN DRUMSTICKS|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00208950000006|POULTRY|MEAT|-81.027334|1.4141937624131469|149|2
34.977331|036729a0ac8cabd38e69ba0b7361e47475210d32|10.02|2014-11-26 12:23:00|1.41290891556208|2|20551900000|149|0.6104695895098807|0|33|2022|-81.027334|505|34.977331|BLUE VEINED CHEESE|0.0|6|BLUE STILTON (FC)|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00205519000002|SPECIALTY CHEESE|DELI|-81.027334|1.4141937624131469|149|1
34.977331|c9cea04d22d789cf3325ac457db3959a48d8a389|3.16|2014-12-16 12:03:00|1.41290891556208|2|20895000000|149|0.6104695895098807|0|33|977|-81.027334|201|34.977331|FRESH HT CHICKEN|0.0|2|HT FRESH CHICKEN DRUMSTICKS|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00208950000006|POULTRY|MEAT|-81.027334|1.4141937624131469|149|1
34.977331|adec3051e2ccb415e42965556ba6dff0255aa9b2|4.19|2014-09-12 11:27:00|1.41290891556208|2|4812127620|149|0.6104695895098807|0|33|1037|-81.027334|164|34.977331|ENGLISH MUFFINS|2.1|7|THOMAS SEASONAL EM PP|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00048121221003|BREAKFAST|COMMERCIAL BAKERY|-81.027334|1.4141937624131469|149|1
34.977331|a85ccff7b86a6de262b9c12e49630a156a616ebb|3.75|2015-01-05 15:03:00|1.41290891556208|2|4610000094|149|0.6104695895098807|0|33|318|-81.027334|52|34.977331|SHREDDED/GRATED CHEESE|1.25|3|SARGENTO CB FOUR STATE CHEDDAR|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00046100011065|CHEESE|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|d39f393704828ad3f5827d625b5d34c3e0a1d0fb|3.65|2014-10-31 11:27:00|1.41290891556208|2|4610000094|149|0.6104695895098807|0|33|318|-81.027334|52|34.977331|SHREDDED/GRATED CHEESE|0.0|3|SARGENTO CB FOUR STATE CHEDDAR|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00046100011065|CHEESE|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|82b97adbec08778c1860abda3c8fde5b590dd9a8|5.78|2014-12-13 11:11:00|1.41290891556208|2|3760007060|149|0.6104695895098807|0|33|714|-81.027334|274|34.977331|MICROWAVE MEALS|0.78|1|DINTY MOORE CMPL BEEF STEW|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00037600070607|PREP FOODS DINNERS|G1 GROCERY|-81.027334|1.4141937624131469|149|2
34.977331|6d95f33d99f9c4a69464a004ca48bf547c0d2774|4.19|2014-11-09 11:36:00|1.41290891556208|2|4125875120|149|0.6104695895098807|0|33|211|-81.027334|33|34.977331|BOUILLON|0.0|1|WYLERS BOUILLON BEEF GRANULES|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00041258751191|SOUP|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|fa3083f4e9407deab61a79082dcc15dd130e3984|17.81|2014-10-02 20:22:00|81.02739863253349|2|20895300000|149|35.035533123585651|0|14|977|-80.992182|201|35.103409|FRESH HT CHICKEN|0.0|2|HT FRESH BNLS CHICKEN BREAST|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|35.014943729270243|00208953000003|POULTRY|MEAT|-81.027334|81.027438431055117|88|2
34.977331|529336217c2a607aabd7e7ec87543247fcfe2a59|2.59|2014-11-03 14:34:00|1.41290891556208|2|7203663996|149|0.6104695895098807|0|33|342|-81.027334|57|34.977331|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00072036631299|MILK|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|9ee7e863e134538045d43848bb40ee2316453865|5.89|2014-09-17 12:14:00|1.41290891556208|2|20600100000|149|0.6104695895098807|0|33|1802|-81.027334|400|34.977331|FFM HAM|2.36|6|VIRGINIA BAKED HAM|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00206001000005|FFM MEAT|DELI|-81.027334|1.4141937624131469|149|1
34.977331|74854b196332ea36d769b9e33faf5e732c6dec2f|11.98|2015-01-13 11:06:00|1.41290891556208|2|8981900171|149|0.6104695895098807|0|33|9934|-81.027334|885|34.977331|NFS POP CHARDONNAY|0.0|13|BERINGER CHARDONNAY|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00089819001712|POPULAR (4-$7.99)|WINE|-81.027334|1.4141937624131469|149|2
34.977331|2bceb1c6b0826c78a2c8a66bfb59d09ffb148686|5.09|2015-01-15 19:59:00|1.41290891556208|2|20600100000|149|0.6104695895098807|0|33|1802|-81.027334|400|34.977331|FFM HAM|0.0|6|VIRGINIA BAKED HAM|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00206001000005|FFM MEAT|DELI|-81.027334|1.4141937624131469|149|1
34.977331|5c3d5a3059b392fba18e978afbb88d7c99d53ad6|1.99|2015-02-06 13:49:00|1.41290891556208|2|60322422423|149|0.6104695895098807|0|33|533|-81.027334|64|34.977331|FRESH PEPPERS|0.0|4|MINI SWEET PEPPERS 1LB|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00603224224230|FRESH PRODUCE|PRODUCE|-81.027334|1.4141937624131469|149|1
34.977331|6e212126aed21746ddb7fd3656f040a1e13878fa|5.39|2015-02-22 19:02:00|1.41290891556208|2|20600200000|149|0.6104695895098807|0|33|1802|-81.027334|400|34.977331|FFM HAM|2.7|6|HONEY CURED HAM|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00206002000004|FFM MEAT|DELI|-81.027334|1.4141937624131469|149|1
34.977331|aac83b6539b1001ea960da3f58dbbb676844e7e3|5.49|2014-12-02 12:38:00|1.41290891556208|2|7203695136|149|0.6104695895098807|0|33|1687|-81.027334|385|34.977331|THAW & SELL (SWEET GOODS)|0.0|14|FUDGE BROWNIE|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00072036951366|SWEET GOODS|BAKERY|-81.027334|1.4141937624131469|149|1
34.977331|54e93b38718b528db5c5adefdacf95b758795366|1.69|2014-12-07 14:16:00|1.41290891556208|2|7203688003|149|0.6104695895098807|0|33|527|-81.027334|64|34.977331|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00072036880031|FRESH PRODUCE|PRODUCE|-81.027334|1.4141937624131469|149|1
34.977331|9c8a988cc374529dbc2801edf1f71f49dba77ee0|6.79|2014-12-06 18:54:00|1.41290891556208|2|7203000314|149|0.6104695895098807|0|33|1685|-81.027334|385|34.977331|ENTENMANNS (SWEET GOODS)|3.39|14|ENT CHS DANISH TWIST PP|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00072030003146|SWEET GOODS|BAKERY|-81.027334|1.4141937624131469|149|1
34.977331|f97b7375bdba94a7d2a7d6f7ddf44ae255f120e6|9.99|2014-09-27 11:26:00|1.41290891556208|2|7203661033|149|0.6104695895098807|0|33|666|-81.027334|145|34.977331|PACKAGED COOKED|0.0|12|HT COOKED SHRIMP RING 10OZ|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00072036610331|SHRIMP|SEAFOOD|-81.027334|1.4141937624131469|149|1
34.977331|28d71a676a3d95e7418f5d36c35c8fee5a259256|2.59|2014-10-23 14:49:00|1.41290891556208|2|7203663996|149|0.6104695895098807|0|33|342|-81.027334|57|34.977331|FRESH MILK|0.0|3|HARRIS TEETER 2%   MILK|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00072036639998|MILK|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|016bbee2806bdff06febdaccbf921ea1d8171be2|2.69|2014-12-23 14:01:00|1.41290891556208|2|7225001125|149|0.6104695895098807|0|33|1025|-81.027334|162|34.977331|WHITE|0.0|7|MERITA OLD FASHIONED 20 OZ|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00072250011259|SLICED BREAD|COMMERCIAL BAKERY|-81.027334|1.4141937624131469|149|1
34.977331|1192261cf9a91ba89ded3b3892c67669b2e74d8c|3.69|2014-10-15 11:47:00|1.41290891556208|2|1380015173|149|0.6104695895098807|0|33|1279|-81.027334|48|34.977331|SINGLE SERVE FLAVOR|0.0|5|STOUFFER PEPP FRENCH BRD PIZZA|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00013800151735|FROZEN MEALS|FROZEN|-81.027334|1.4141937624131469|149|1
34.977331|9900b5d7e9a66ce079d61b263276a38079dfdd79|3.18|2014-09-29 13:40:00|1.41290891556208|2|2400016299|149|0.6104695895098807|0|33|247|-81.027334|39|34.977331|VEGETABLES-FLANKER|0.0|1|DEL MONTE SAUERKRAUT|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00024000163145|VEGETABLES-CAN/JAR|G1 GROCERY|-81.027334|1.4141937624131469|149|2
34.977331|a50487ea022515afc60c084b3f82ecb821bc417d|4.79|2015-03-04 12:54:00|1.41290891556208|2|1200000514|149|0.6104695895098807|0|33|54|-81.027334|8|34.977331|DIET|0.79|23|DT PEPSI 16.9OZ 6PK|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00012000504068|CARBONATED BEVERAGES|BEVERAGE|-81.027334|1.4141937624131469|149|1
34.977331|5e0044a55170f62d18b1953431634eb7a41585ee|5.38|2014-10-03 12:28:00|1.41290891556208|2|1480000034|149|0.6104695895098807|0|33|128|-81.027334|20|34.977331|APPLE JUICE-SHELF|0.0|1|MOTTS 100% PURE APPLE JUICE|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00014800000344|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-81.027334|1.4141937624131469|149|2
34.977331|902409e9fdb705776512dcc9ec5975d7b08d410d|5.59|2014-09-11 12:51:00|1.41290891556208|2|20165900000|149|0.6104695895098807|0|33|297|-81.027334|49|34.977331|GROUND BEEF|1.6|2|GROUND BEEF 93% LEAN|6150df3f32f775df5ea632c145c5f67b2ac3e8f2|4.021630529911472|0.61055446569467375|00201659000001|BEEF|MEAT|-81.027334|1.4141937624131469|149|1
35.43259|b744489eceda30b111cc70a25de77f2d29bc7f7b|1.79|2015-02-21 11:04:00|80.606823361882718|3|5100001047|202|35.49048122497333|0|57|212|-80.662946|33|35.412407|CONDENSED SOUP|0.54|1|CAMP COND NEW ENG CLAM CHOWDER|6540bca0a640122cd53d6500abeea4a65d0fefa4|4.00014428878895|35.500309569604553|00051000013675|SOUP|G1 GROCERY|-80.605588|80.605621541959607|68|1
35.43259|740996160522260feb646e3f5ea7b375e430004d|1.79|2014-10-25 11:46:00|1.4057311447477159|3|5100001047|202|0.6184153580092175|0|52|212|-80.605588|33|35.43259|CONDENSED SOUP|0.79|1|CAMP COND NEW ENG CLAM CHOWDER|6540bca0a640122cd53d6500abeea4a65d0fefa4|4.00014428878895|0.6209993146566879|00051000013675|SOUP|G1 GROCERY|-80.605588|1.406832906106031|202|1
35.43259|4c002f4157c6b8b32db0eba655122361311c8bd1|8.35|2015-02-07 09:09:00|80.606823361882718|3|76211188813|202|35.49048122497333|0|57|37|-80.662946|10|35.412407|PODS/CUPS/SINGLES|1.36|1|STARBUCKS CAFFEE VERONA KCUPS|6540bca0a640122cd53d6500abeea4a65d0fefa4|4.00014428878895|35.500309569604553|00762111930255|COFFEE|G1 GROCERY|-80.605588|80.605621541959607|68|1
35.43259|460b798123c1f36622ba9fb02cbc4c301a91c4da|6.949999999999999|2014-10-04 13:31:00|80.606823361882718|3|3940001606|202|35.49048122497333|0|57|243|-80.662946|39|35.412407|BAKED BEANS|1.9500000000000002|1|BUSH BKD BEAN EZO VEG|6540bca0a640122cd53d6500abeea4a65d0fefa4|4.00014428878895|35.500309569604553|00039400016304|VEGETABLES-CAN/JAR|G1 GROCERY|-80.605588|80.605621541959607|68|5
35.43259|dffb990123b3a86dd46ecefb948f1d4c18995d9e|1.89|2014-11-09 12:01:00|1.4057311447477159|3|4600086031|202|0.6184153580092175|0|52|77|-80.605588|272|35.43259|HISP SAUCES/SEASONINGS|0.0|1|OEP ENCHILADA SC MILD|6540bca0a640122cd53d6500abeea4a65d0fefa4|4.00014428878895|0.6209993146566879|00046000860312|HISPANIC PREP. FOODS|G1 GROCERY|-80.605588|1.406832906106031|202|1
35.43259|9fbb12382f1635fcb07b442c72590d4340103b93|1.89|2014-11-08 15:00:00|1.4057311447477159|3|4600086031|202|0.6184153580092175|0|52|77|-80.605588|272|35.43259|HISP SAUCES/SEASONINGS|0.0|1|OEP ENCHILADA SC MILD|6540bca0a640122cd53d6500abeea4a65d0fefa4|4.00014428878895|0.6209993146566879|00046000860312|HISPANIC PREP. FOODS|G1 GROCERY|-80.605588|1.406832906106031|202|1
35.43259|0eb09ca806be422c5b6b5e9cca174c55a8557d84|14.7|2014-11-15 09:44:00|80.606823361882718|3|4470002268|202|35.49048122497333|0|57|358|-80.662946|100|35.412407|REGULAR BACON|3.68|19|OSCAR MAYER SLICED BACON|6540bca0a640122cd53d6500abeea4a65d0fefa4|4.00014428878895|35.500309569604553|00044700019887|BACON|CASE READY MEATS|-80.605588|80.605621541959607|68|2
35.43259|fa8c8da73bb2e84c1cfef68c79062b95e4554698|4.13|2014-11-02 10:58:00|80.606823361882718|3||202|35.49048122497333|0|57|500|-80.662946|64|35.412407|FRESH APPLES|0.0|4|RED DEL APPLE, WA  48|6540bca0a640122cd53d6500abeea4a65d0fefa4|4.00014428878895|35.500309569604553|00233284000002|FRESH PRODUCE|PRODUCE|-80.605588|80.605621541959607|68|1
35.43259|080f664bf04c986ebc9746638b1547e0810a76e3|4.23|2014-12-14 12:41:00|1.4057311447477159|3||202|0.6184153580092175|0|52|500|-80.605588|64|35.43259|FRESH APPLES|0.0|4|RED DEL APPLE, WA  48|6540bca0a640122cd53d6500abeea4a65d0fefa4|4.00014428878895|0.6209993146566879|00233284000002|FRESH PRODUCE|PRODUCE|-80.605588|1.406832906106031|202|1
35.43259|7731c18622c555e06186edc8afcfeef6f2407df8|2.45|2014-09-27 11:30:00|1.4057311447477159|3|7203663217|202|0.6184153580092175|0|52|330|-80.605588|55|35.43259|EGGS|0.45|3|HT GRADE A LARGE EGGS 18 CT|6540bca0a640122cd53d6500abeea4a65d0fefa4|4.00014428878895|0.6209993146566879|00072036632173|EGGS FRESH|DAIRY|-80.605588|1.406832906106031|202|1
35.43259|3acc964e122fa3c300c08937b8cc42263cd2486f|5.38|2015-03-07 12:17:00|80.606823361882718|3|7203663217|202|35.49048122497333|0|57|330|-80.662946|55|35.412407|EGGS|1.38|3|HT GRADE A LARGE EGGS 18 CT|6540bca0a640122cd53d6500abeea4a65d0fefa4|4.00014428878895|35.500309569604553|00072036632173|EGGS FRESH|DAIRY|-80.605588|80.605621541959607|68|2
35.43259|6c5e71541678766f72cb69dc350acda431ac5d3f|2.79|2015-01-01 13:29:00|80.606823361882718|3|61611227958|202|35.49048122497333|0|57|581|-80.662946|136|35.412407|FRESH SALSA|0.29|4|WHOLLY GUACAMOLE CLASSIC 8OZ|6540bca0a640122cd53d6500abeea4a65d0fefa4|4.00014428878895|35.500309569604553|00616112279588|OTHER MERCHANDISE|PRODUCE|-80.605588|80.605621541959607|68|1
35.43259|a7a7296f237ce579aac7ce46f43fbe2086365912|0.97|2015-01-24 10:03:00|1.4057311447477159|3|7203671102|202|0.6184153580092175|0|52|1025|-80.605588|162|35.43259|WHITE|0.0|7|HT OLD FASHIONED BREAD|6540bca0a640122cd53d6500abeea4a65d0fefa4|4.00014428878895|0.6209993146566879|00072036711021|SLICED BREAD|COMMERCIAL BAKERY|-80.605588|1.406832906106031|202|1
35.43259|1e02e0cd034ddbbdf473666b782ca9d85dd99e80|0.97|2014-09-20 10:55:00|80.606823361882718|3|7203671102|202|35.49048122497333|0|57|1025|-80.662946|162|35.412407|WHITE|0.0|7|HT OLD FASHIONED BREAD|6540bca0a640122cd53d6500abeea4a65d0fefa4|4.00014428878895|35.500309569604553|00072036711021|SLICED BREAD|COMMERCIAL BAKERY|-80.605588|80.605621541959607|68|1
35.43259|384d1e6bd983d430c7073b02820ebf9259731f60|0.97|2015-01-10 11:59:00|80.606823361882718|3|7203671102|202|35.49048122497333|0|57|1025|-80.662946|162|35.412407|WHITE|0.0|7|HT OLD FASHIONED BREAD|6540bca0a640122cd53d6500abeea4a65d0fefa4|4.00014428878895|35.500309569604553|00072036711021|SLICED BREAD|COMMERCIAL BAKERY|-80.605588|80.605621541959607|68|1
35.43259|319f1b8337a351f437adf8e0a886f8d196cdcb03|0.97|2014-12-20 10:42:00|80.606823361882718|3|7203671102|202|35.49048122497333|0|57|1025|-80.662946|162|35.412407|WHITE|0.0|7|HT OLD FASHIONED BREAD|6540bca0a640122cd53d6500abeea4a65d0fefa4|4.00014428878895|35.500309569604553|00072036711021|SLICED BREAD|COMMERCIAL BAKERY|-80.605588|80.605621541959607|68|1
35.43259|1048b8fe399bc17dab31b58b2093d43ec78a750f|3.75|2014-11-14 12:48:00|80.606823361882718|3|7203698557|202|35.490480944828782|0|57|424|-80.810056|72|35.219587|NFS-FACIAL TISSUE|0.75|1|HT FACIAL TISSUE LOTION|6540bca0a640122cd53d6500abeea4a65d0fefa4|4.00014428878895|35.500309569604553|00072036985583|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.605588|80.605811644558685|401|3
35.43259|a0a31b0774e6e8e418720c362653b6a8af0e3d0e|1.99|2014-12-04 18:36:00|1.4057311447477159|3|7203698434|202|0.6184153580092175|0|52|3992|-80.605588|1080|35.43259|DENTAL FLOSSER|0.0|17|(JHK) HT DENTAL FLOSSERS MINT|6540bca0a640122cd53d6500abeea4a65d0fefa4|4.00014428878895|0.6209993146566879|00072036984340|ORAL HYGIENE|HBC|-80.605588|1.406832906106031|202|1
35.43259|f5b5640087d7a0a012b0d64e2a62d1539b88d276|1.89|2014-11-29 10:08:00|80.606823361882718|3|1300079630|202|35.49048122497333|0|57|69|-80.662946|26|35.412407|CANNED GRAVY|0.55|1|HEINZ GRAVY TURKEY HOMESTYLE|6540bca0a640122cd53d6500abeea4a65d0fefa4|4.00014428878895|35.500309569604553|00013000799102|PREPARED FOODS-DRY MIXES|G1 GROCERY|-80.605588|80.605621541959607|68|1
35.43259|cb96b0b7eb58c21aa4da3d4439680967a50c606a|25.98|2015-01-31 12:21:00|80.606823361882718|3|78615000014|202|35.49048122497333|0|57|459|-80.662946|83|35.412407|IMPORT BEER|0.0|16|STELLA ARTOIS 12PK BOTTLES|6540bca0a640122cd53d6500abeea4a65d0fefa4|4.00014428878895|35.500309569604553|00786150000144|IMPORT BEER|BEER|-80.605588|80.605621541959607|68|2
35.43259|77036f150ebd984cbb245452a8bdcc7860ab5873|28.96|2015-02-01 16:48:00|80.606823361882718|3|3410057243|202|35.49048122497333|0|57|455|-80.662946|82|35.412407|DOMESTIC PREMIUM 12PK&>|0.0|16|MILLER LITE HIGH GRAPHICS 24PK|6540bca0a640122cd53d6500abeea4a65d0fefa4|4.00014428878895|35.500309569604553|00034100572433|DOMESTIC BEER|BEER|-80.605588|80.605621541959607|68|2
35.43259|a38ccf8b73804951f91f515235381d5694f98dcf|14.99|2014-11-26 13:56:00|80.606823361882718|3|3410057243|202|35.49048122497333|0|57|455|-80.662946|82|35.412407|DOMESTIC PREMIUM 12PK&>|0.0|16|MILLER LITE HIGH GRAPHICS 24PK|6540bca0a640122cd53d6500abeea4a65d0fefa4|4.00014428878895|35.500309569604553|00034100572433|DOMESTIC BEER|BEER|-80.605588|80.605621541959607|68|1
35.124987|5f410c27f3882e1df306bdcb9eb8f648604f1dac|3.99|2014-11-09 17:29:00|80.709550101431233|3|8043210346|157|35.16598669365937|0|43|462|-80.737839|84|35.297134|WINE COOLERS SPRITZER|0.0|16|SEAGRAMS JAMAICAN ME HAPPY 4PK|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00080432103463|SPECIALTY|BEER|-80.709466|80.709549397642547|258|1
35.124987|31be5deb4f20bdc1bdbc4428863084332e51530c|2.0|2014-12-21 18:48:00|80.709550101431233|3||157|35.16598669365937|0|43|511|-80.737839|64|35.297134|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00204770000004|FRESH PRODUCE|PRODUCE|-80.709466|80.709549397642547|258|1
35.124987|4bd88004ad45dbf467b47e6d57f85f94ea7dae8c|2.0|2014-11-04 20:07:00|80.709550101431233|3||157|35.16598669365937|0|43|511|-80.737839|64|35.297134|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00204770000004|FRESH PRODUCE|PRODUCE|-80.709466|80.709549397642547|258|1
35.124987|5402a38c98e18f5020267904ad03d8a914628871|2.0|2014-09-21 17:24:00|80.709550101431233|3||157|35.165986691485259|0|43|511|-80.780702|64|35.318911|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00204770000004|FRESH PRODUCE|PRODUCE|-80.709466|80.709550981167098|167|1
35.124987|222f2d84b217705715136e04fcdf26ba8f9c74e8|2.0|2014-11-16 17:28:00|80.709550101431233|3||157|35.16598669365937|0|43|511|-80.737839|64|35.297134|FRESH AVOCADOS|0.21|4|AVOCADOS, HASS XL 36CT|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00204770000004|FRESH PRODUCE|PRODUCE|-80.709466|80.709549397642547|258|1
35.124987|b93b0ad9352c0e1bfad5db0130644fa41eeeb347|2.0|2015-01-11 19:42:00|80.709550101431233|3||157|35.16598669365937|0|43|511|-80.737839|64|35.297134|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00204770000004|FRESH PRODUCE|PRODUCE|-80.709466|80.709549397642547|258|1
35.124987|dea92f497eb0a9100f11921b776f8b42ab2db0ec|2.0|2014-12-27 20:13:00|80.709550101431233|3||157|35.16598669365937|0|43|511|-80.737839|64|35.297134|FRESH AVOCADOS|0.75|4|AVOCADOS, HASS XL 36CT|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00204770000004|FRESH PRODUCE|PRODUCE|-80.709466|80.709549397642547|258|1
35.124987|aae8b7503e92d2f5f3ce000d7ac0577f1e28659e|1.14|2015-01-02 19:32:00|80.709550101431233|3||157|35.16598669365937|0|43|523|-80.737839|64|35.297134|FRESH POTATOES|0.0|4|COO RUSSET POTATOES, BULK|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00204072000009|FRESH PRODUCE|PRODUCE|-80.709466|80.709549397642547|258|1
35.124987|6168e53bac458e2ef81c54cb57abc63961184014|2.0|2014-11-23 15:47:00|80.709550101431233|3||157|35.16598669365937|0|43|511|-80.737839|64|35.297134|FRESH AVOCADOS|0.11|4|AVOCADOS, HASS XL 36CT|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00204770000004|FRESH PRODUCE|PRODUCE|-80.709466|80.709549397642547|258|1
35.124987|af154ecc332b5a6a3497ca81622d8f48e295de3e|2.0|2014-09-10 19:36:00|80.709550101431233|3||157|35.16598669365937|0|43|511|-80.737839|64|35.297134|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00204770000004|FRESH PRODUCE|PRODUCE|-80.709466|80.709549397642547|258|1
35.124987|490f7d46ca27126c00dea23ce323d744e389005d|2.0|2014-09-11 16:12:00|80.709550101431233|3||157|35.16598669365937|0|43|511|-80.737839|64|35.297134|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00204770000004|FRESH PRODUCE|PRODUCE|-80.709466|80.709549397642547|258|1
35.124987|c11a007e8b8dc7f4c239175ddb411ca60f8f1ef2|2.0|2014-11-13 19:32:00|80.709550101431233|3||157|35.16598669365937|0|43|511|-80.737839|64|35.297134|FRESH AVOCADOS|0.21|4|AVOCADOS, HASS XL 36CT|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00204770000004|FRESH PRODUCE|PRODUCE|-80.709466|80.709549397642547|258|1
35.124987|8da17ccd40c7f03227af2eefb4647e32b0b861b9|2.0|2014-10-10 17:53:00|80.709550101431233|3||157|35.16598669365937|0|43|511|-80.737839|64|35.297134|FRESH AVOCADOS|0.5|4|AVOCADOS, HASS XL 36CT|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00204770000004|FRESH PRODUCE|PRODUCE|-80.709466|80.709549397642547|258|1
35.124987|c2a80558ac20c6c6a20529437d20430c4df21e17|2.0|2014-12-07 15:02:00|80.709550101431233|3||157|35.16598669365937|0|43|511|-80.737839|64|35.297134|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00204770000004|FRESH PRODUCE|PRODUCE|-80.709466|80.709549397642547|258|1
35.124987|461c4fcfadd5a4ca7e493e5a29eccf1c2489d933|2.0|2014-09-25 18:49:00|80.709550101431233|3||157|35.16598669365937|0|43|511|-80.737839|64|35.297134|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00204770000004|FRESH PRODUCE|PRODUCE|-80.709466|80.709549397642547|258|1
35.124987|3ee3137a463cb70bfb934d7c7a2e55df42cdd9b3|2.0|2015-01-31 17:42:00|80.709550101431233|3||157|35.165986691485259|0|43|511|-80.780702|64|35.318911|FRESH AVOCADOS|0.75|4|AVOCADOS, HASS XL 36CT|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00204770000004|FRESH PRODUCE|PRODUCE|-80.709466|80.709550981167098|167|1
35.124987|c751791d925643c6d7da32df1361d9865e38e4ce|3.5|2014-12-07 18:34:00|80.709550101431233|3|7203603041|157|35.165986691485259|0|43|220|-80.780702|34|35.318911|PEPPER|1.0|1|E  HT BLACK PEPPER|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00072036030412|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.709466|80.709550981167098|167|1
35.124987|8ce247178a041263bca2497b6267fd3efa6f2cdb|3.99|2015-01-11 20:05:00|80.709550101431233|3|7127927100|157|35.16598669365937|0|43|555|-80.737839|64|35.297134|PACKAGED SALADS|0.0|4|F.E. BABY SPINACH|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00071279271002|FRESH PRODUCE|PRODUCE|-80.709466|80.709549397642547|258|1
35.124987|916c1cecd1e1f93df950e8f1bbddb31c702f54c1|0.84|2015-02-15 17:03:00|80.709550101431233|3||157|35.16598669365937|0|43|524|-80.737839|64|35.297134|FRESH PROD FRESH ONIONS|0.0|4|COO SHALLOTS, BULK|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00204662000006|FRESH PRODUCE|PRODUCE|-80.709466|80.709549397642547|258|1
35.124987|e50c7140c5be547a9026f8727f569bdc90109075|5.03|2014-09-25 19:15:00|80.709550101431233|3|20927000000|157|35.16598669365937|0|43|668|-80.737839|146|35.297134|LEGS/CLUSTERS|2.53|12|ROCK CRAB CLUSTERS (CA)|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00209270000004|CRAB|SEAFOOD|-80.709466|80.709549397642547|258|1
35.124987|16eca134da0aff33e08067402a5515b2cee5fba1|0.95|2014-10-09 18:36:00|80.709550101431233|3|4600028869|157|35.16598669365937|0|43|77|-80.737839|272|35.297134|HISP SAUCES/SEASONINGS|0.0|1|OEP SEASONING TACO HOT & SPICY|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00046000288758|HISPANIC PREP. FOODS|G1 GROCERY|-80.709466|80.709549397642547|258|1
35.124987|1424c13bf4a79720e38837dc038571587c245635|1.79|2014-12-26 19:54:00|80.709550101431233|3|7203688032|157|35.16598669365937|0|43|555|-80.737839|64|35.297134|PACKAGED SALADS|0.0|4|HT SHREDDED ICEBERG LETTUCE|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00072036880321|FRESH PRODUCE|PRODUCE|-80.709466|80.709549397642547|258|1
35.124987|f4366d67493ce459d9907e446adaefe8842aaf4a|3.29|2015-03-09 15:30:00|80.709550101431233|3|2840014741|157|35.16598669365937|0|43|205|-80.737839|31|35.297134|REMAINING SNACKS|0.29|1|SUNCHIPS REGULAR|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00028400147415|SNACKS|G1 GROCERY|-80.709466|80.709549397642547|258|1
35.124987|35e6615ce609398fb153d35b67106d92893f2214|6.79|2015-01-01 12:20:00|80.709550101431233|3|4850001833|157|35.16598669365937|0|43|335|-80.737839|56|35.297134|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA HOMESTYLE|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00048500018293|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.709466|80.709549397642547|258|1
35.124987|7c198002c4dadf5a15f661de54395f52d774d82d|4.29|2015-03-08 16:49:00|80.709550101431233|3|4178000011|157|35.16598669365937|0|43|201|-80.737839|31|35.297134|POTATO CHIPS|1.3|1|UTZ RED HOT CHIP|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00041780001887|SNACKS|G1 GROCERY|-80.709466|80.709549397642547|258|1
35.124987|8423020811a7631b51efe0c0a9b52d631d4a5da8|4.29|2015-02-05 16:22:00|80.709550101431233|3|4178000011|157|35.165986691485259|0|43|201|-80.780702|31|35.318911|POTATO CHIPS|1.3|1|UTZ RED HOT CHIP|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00041780001887|SNACKS|G1 GROCERY|-80.709466|80.709550981167098|167|1
35.124987|547ac78e86579eeab96972713bbfa493310f76f9|11.98|2014-12-28 19:20:00|80.709550101431233|3|20931700000|157|35.16598669365937|0|43|676|-80.737839|148|35.297134|TAILS|0.0|12|WC LOBSTER TAILS 4.2 OZ  (CA)|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00209317000004|LOBSTERS|SEAFOOD|-80.709466|80.709549397642547|258|1
35.124987|d1ac9fa006b9ee2caf07b6b86fe08c139bae0c13|2.99|2014-11-01 17:52:00|80.709550101431233|3|2858800400|157|35.16598669365937|0|43|5846|-80.737839|1538|35.297134|KITCHEN GADGETS BARWARE|0.6|18|OENO. PICNIC CORKSCREW|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00028588004005|KITCHEN GADGETS|GM|-80.709466|80.709549397642547|258|1
35.124987|914c1860ff64c9672bf20d38677dc4de2d60c7bf|4.29|2014-09-17 10:02:00|80.709550101431233|3|7343500004|157|35.16598669365937|0|43|1631|-80.737839|373|35.297134|THAW & SELL (ROLLS)|0.0|14|KING'S HAWAIIAN 12CT ROLLS|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00073435000044|ROLLS|BAKERY|-80.709466|80.709549397642547|258|1
35.124987|253db27dcc57b35e2445dac0300ca59b07dca09a|1.69|2014-10-21 17:46:00|80.709550101431233|3|7680828008|157|35.16598669365937|0|43|149|-80.737839|23|35.297134|WHSE PASTA CORE|0.31|1|BARILLA PASTA LINGUINI|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00076808280173|PASTA|G1 GROCERY|-80.709466|80.709549397642547|258|1
35.124987|c4a93fa62cae86ad1cbd1532df96bcfe7928fa64|2.49|2015-02-04 19:24:00|80.709550101431233|3|7203688213|157|35.16598669365937|0|43|555|-80.737839|64|35.297134|PACKAGED SALADS|0.0|4|HT BABY SPINACH|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00072036882134|FRESH PRODUCE|PRODUCE|-80.709466|80.709549397642547|258|1
35.124987|0b01b054b455b2413dec5880cf6befc80935f506|4.49|2014-10-12 13:52:00|80.709550101431233|3|71575620002|157|35.16598669365937|0|43|504|-80.737839|64|35.297134|FRESH BERRIES|0.5|4|STRAWBERRIES 1LB CLAM|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00665290001184|FRESH PRODUCE|PRODUCE|-80.709466|80.709549397642547|258|1
35.124987|645dd7359b327a406810baa38fc593680c42f221|1.79|2015-01-12 19:27:00|80.709550101431233|3|2830000089|157|35.16598669365937|0|43|1134|-80.737839|57|35.297134|CARTON MILK|0.0|3|SHAMROCK FARMS 2% MILK|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00028300000902|MILK|DAIRY|-80.709466|80.709549397642547|258|1
35.124987|947873ed0574a4e89c9f18143637efa8bbc8eca5|1.25|2014-11-25 10:04:00|80.709550101431233|3|4900005537|157|35.16598669365937|0|43|55|-80.737839|8|35.297134|REGULAR|0.26|23|SPRITE 1.25 LITER BOTTLE|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00049000055450|CARBONATED BEVERAGES|BEVERAGE|-80.709466|80.709549397642547|258|1
35.124987|d7bf965bf1a3aff80939fe20c087d6da5be7f66b|0.79|2014-11-09 17:26:00|80.709550101431233|3||157|35.16598669365937|0|43|532|-80.737839|64|35.297134|FRESH CUCUMBERS|0.2|4|COO CUCUMBERS S/S|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00204062000002|FRESH PRODUCE|PRODUCE|-80.709466|80.709549397642547|258|1
35.124987|b122ce38e787feb8f8bc539ce7b61f928f92eea8|9.99|2014-12-05 22:25:00|80.709550101431233|3|3410057509|157|35.16598669365937|0|43|455|-80.737839|82|35.297134|DOMESTIC PREMIUM 12PK&>|0.0|16|MILLER LITE 12PK 12OZ BTL|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00034100575090|DOMESTIC BEER|BEER|-80.709466|80.709549397642547|258|1
35.124987|27b70f405b85d44d946d415242798d3ca4719a2d|2.15|2014-12-23 20:23:00|80.709550101431233|3|7142909849|157|35.16598669365937|0|43|238|-80.737839|38|35.297134|RICE FLAVORED|0.16|1|ZAT RICE RED BEANS|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00071429098497|RICE GRAINS AND BEANS|G1 GROCERY|-80.709466|80.709549397642547|258|1
35.124987|e5a82ae37959e268549f2f64c30187ea825faac4|9.98|2014-10-26 19:03:00|80.709550101431233|3|71575620002|157|35.16598669365937|0|43|504|-80.737839|64|35.297134|FRESH BERRIES|2.49|4|STRAWBERRIES 1LB CLAM|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00071430007525|FRESH PRODUCE|PRODUCE|-80.709466|80.709549397642547|258|2
35.124987|2d3d08d4fd4e4f3554f3403bfa860c9e38f72e60|1.79|2015-01-12 19:36:00|80.709550101431233|3|5200033875|157|35.16598669365937|0|43|171|-80.737839|20|35.297134|ISOTONIC DRINKS|0.41|1|GATORADE AM TROPICAL MANGO|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00052000322132|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.709466|80.709549397642547|258|1
35.124987|b2fbaf197e121ec30c2d1c940109de0e3208e701|4.29|2014-10-21 17:53:00|80.709550101431233|3|2100061531|157|35.16598669365937|0|43|333|-80.737839|52|35.297134|PARMESAN CHEESE|0.79|3|KRAFT GRATED PARMESAN CHEESE|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00021000615315|CHEESE|DAIRY|-80.709466|80.709549397642547|258|1
35.124987|00dbdecf0530b545658f3ffa3c1703305e064edf|14.97|2015-01-31 17:57:00|80.709550101431233|3|20931900000|157|35.16598669365937|0|43|676|-80.737839|148|35.297134|TAILS|0.0|12|WC LOBSTER TAILS 2/3 OZ  (CA)|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00209319000002|LOBSTERS|SEAFOOD|-80.709466|80.709549397642547|258|1
35.124987|197e9b3eeab1b56160834daffaa416f38271dfda|1.89|2014-10-15 19:50:00|80.709550101431233|3|7203663202|157|35.16598669365937|0|43|1262|-80.737839|57|35.297134|HALF N HALF WHIPPING CREAM|0.0|3|HT HEAVY WHIPPING CREAM|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00072036631268|MILK|DAIRY|-80.709466|80.709549397642547|258|1
35.124987|1520b65818d73b901796c36d92284a844d248813|1.89|2014-10-15 20:35:00|80.709550101431233|3|7203663202|157|35.16598669365937|0|43|1262|-80.737839|57|35.297134|HALF N HALF WHIPPING CREAM|0.0|3|HT HEAVY WHIPPING CREAM|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00072036631268|MILK|DAIRY|-80.709466|80.709549397642547|258|1
35.124987|ded37e1499a64ff5e98bbf7781e6f6b2b3e447f2|1.99|2014-10-09 19:12:00|80.709550101431233|3|4600081101|157|35.16598669365937|0|43|1213|-80.737839|272|35.297134|HISP DINNERS/SHELLS|0.0|1|OEP SHELL TACO 12CT|67a8d72d162b7928ffeb1670921799526cf5a786|2.832983739829059|35.165986692693096|00046000811017|HISPANIC PREP. FOODS|G1 GROCERY|-80.709466|80.709549397642547|258|1
35.667941|46f70dad6b893512462276ad998264b977c4e6eb|3.29|2015-02-27 17:01:00|1.4057311447477159|4|7410814498|178|0.6225230078570788|0|52|3650|-80.497332|1060|35.667941|COMB|0.0|17|CNR COMB 3PK ASST PRO STYLE|6866a4386ace8338ae5d257b0a2761ad443fa407|2.6513195023021012|0.6209993146566879|00074108144980|HAIR CARE ACCESSORIES|HBC|-80.497332|1.4049434824709919|178|1
35.667941|063499bcb73c3b4de747952df8d767ce1a2c6a0b|1.69|2014-10-27 18:15:00|80.497482303704658|4|4900000044|178|35.706311386212505|0|6|54|-80.746334|8|35.41832|DIET|0.0|23|CB COKE ZERO 20 OZ|6866a4386ace8338ae5d257b0a2761ad443fa407|2.6513195023021012|35.699188602026126|00049000040869|CARBONATED BEVERAGES|BEVERAGE|-80.497332|80.497508367172784|190|1
35.667941|f5b52d771545780e0b24a9e51a2c3d4f37b8a32c|1.69|2014-11-22 15:20:00|1.4057311447477159|4|1200000129|178|0.6225230078570788|0|52|55|-80.497332|8|35.667941|REGULAR|0.0|23|CB PEPSI COLA 20 0Z|6866a4386ace8338ae5d257b0a2761ad443fa407|2.6513195023021012|0.6209993146566879|00012000001291|CARBONATED BEVERAGES|BEVERAGE|-80.497332|1.4049434824709919|178|1
35.667941|8b3fc447eb59213d15b14ec3d70109627613a801|3.29|2014-10-03 18:01:00|1.4057311447477159|4|7203698555|178|0.6225230078570788|0|52|427|-80.497332|72|35.667941|NFS-TOILET TISSUE|0.5|1|HT 1000 SHEET BATHTISSUE 4 RL|6866a4386ace8338ae5d257b0a2761ad443fa407|2.6513195023021012|0.6209993146566879|00072036985552|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|8117ccbad19c8967478378b198ef87a522eccd96|2.91|2014-10-01 09:33:00|1.4057311447477159|4|7203603070|178|0.6225230078570788|0|52|29|-80.497332|3|35.667941|REMAINING BAKING SUPPLIES|0.0|1|HT PURE CORN STRCH|6866a4386ace8338ae5d257b0a2761ad443fa407|2.6513195023021012|0.6209993146566879|00072036030702|BAKING SUPPLIES|G1 GROCERY|-80.497332|1.4049434824709919|178|3
35.667941|84de6f50b85d19abbf2e2299729f711759be4530|0.97|2014-12-18 22:21:00|1.4057311447477159|4|7203603070|178|0.6225230078570788|0|52|29|-80.497332|3|35.667941|REMAINING BAKING SUPPLIES|0.0|1|HT PURE CORN STRCH|6866a4386ace8338ae5d257b0a2761ad443fa407|2.6513195023021012|0.6209993146566879|00072036030702|BAKING SUPPLIES|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.04711|d1885de7d80c53b70823f068066adf05005b3dad|2.69|2015-02-05 17:15:00|80.648225123995502|0|1450000253|129|35.076324003421938|0|30|1272|-80.758228|50|34.95459|BAG VEG STEAM|1.35|5|BE STEAMFRESH PREM BROCC FLRTS|696d084228372a53def6770c09e8923e281da0bb|2.0186192474650415|35.078006462436761|00014500011831|VEGETABLES-FROZEN|FROZEN|-80.64817|80.64822221554607|182|1
35.103409|d30c55c6841492fb26069e32e825637cafaf1953|0.99|2015-01-23 20:05:00|1.4132775322775095|3|7397010202|88|0.6126700657242101|0|58|55|-80.992182|8|35.103409|REGULAR|0.0|23|DR BROWNS ROOT BEER SODA|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00073970102067|CARBONATED BEVERAGES|BEVERAGE|-80.992182|1.413580244274486|88|1
35.103409|7476ba077fbc184ad651f64475dbd15eb560e2c7|7.35|2015-02-15 11:18:00|1.4132775322775095|3|4470002268|88|0.6126700657242101|0|58|358|-80.992182|100|35.103409|REGULAR BACON|3.68|19|OSCAR MAYER SLICED BACON|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00044700019887|BACON|CASE READY MEATS|-80.992182|1.413580244274486|88|1
35.103409|bb5d327f5c95a4f0b76bc811a820822a07a13ac3|8.58|2014-11-28 12:57:00|1.4132775322775095|3|4400003037|88|0.6126700657242101|0|58|90|-80.992182|13|35.103409|SNACK CRACKERS|2.15|1|WHEAT THINS RANCH|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00044000030421|CRACKERS|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|1a6a382469bba64649fad136eaf4169c72e0aabf|4.39|2015-01-29 20:48:00|1.4132775322775095|3|4400003037|88|0.6126700657242101|0|58|90|-80.992182|13|35.103409|SNACK CRACKERS|2.2|1|WHEAT THINS RANCH|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00044000030421|CRACKERS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|95c8a873b0a5f1e705fbe70e458d8a6e48f4a2fc|2.65|2014-12-07 20:58:00|1.4132775322775095|3|5150000094|88|0.6126700657242101|0|58|126|-80.992182|19|35.103409|PRESERVES/MARMALADE|0.0|1|SMUCKER STRAWBERRY PRESERVES|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00051500000953|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|79715d0f6087843a69e78b4c1ad376cbd3a8a19c|1.29|2015-02-07 21:28:00|1.4132775322775095|3|4920005675|88|0.6126700657242101|0|58|224|-80.992182|35|35.103409|SUGAR-BROWN|0.3|1|DOMINO DARK BROWN SUGAR-BX|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00049200056004|SUGAR/SUBSTITUTES|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|6825c79125876c32583737136007c3d601de4032|10.08|2015-01-09 19:14:00|1.4132775322775095|3|20895300000|88|0.6126700657242101|0|58|977|-80.992182|201|35.103409|FRESH HT CHICKEN|6.06|2|HT FRESH BNLS CHICKEN BREAST|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00208953000003|POULTRY|MEAT|-80.992182|1.413580244274486|88|1
35.103409|57e3ca07d4e18b0af6ee9dc85ff8116fd4f6b9a8|4.69|2014-12-24 12:25:00|1.4132775322775095|3|79452220065|88|0.6126700657242101|0|58|235|-80.992182|37|35.103409|GREEN TEA|1.19|1|TAZO BERRYBLOSSOM WHITE TEA|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00794522212019|TEA|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|13ab58d9df0aeeff52a3b75f79c893ab52a05ef5|4.8|2014-11-19 14:01:00|1.4132775322775095|3|2400001738|88|0.6126700657242101|0|58|257|-80.992182|39|35.103409|TOMATOES|0.2|1|DEL MONTE TOMATO CHILI STYLE|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00024000012672|VEGETABLES-CAN/JAR|G1 GROCERY|-80.992182|1.413580244274486|88|4
35.103409|9c8796b90936bcc3c244bb2e11f6185ae91b7c38|4.49|2014-09-15 00:38:00|1.4132775322775095|3|2620016236|88|0.6126700657242101|0|58|215|-80.992182|31|35.103409|JERKY SNACKS|0.0|1|SLIM JIM ORIGINAL 15 CT|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00026200162362|SNACKS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|f549820975e5b84e39bc506792737487be901b15|3.15|2015-02-09 00:06:00|80.992192682720116|3|7265500105|88|35.105739325068221|0|56|1278|-81.027334|48|34.977331|SINGLE SERVE NUTRITIONAL|0.65|5|HC CAFE STEAMER SWTSPC ORN CHK|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|35.113093007298254|00072655001091|FROZEN MEALS|FROZEN|-80.992182|80.99218618486077|149|1
35.103409|ae6793884d621308b3bd77f980c68587346a9682|3.25|2015-01-18 15:10:00|1.4132775322775095|3|7203656080|88|0.6126700657242101|0|58|318|-80.992182|52|35.103409|SHREDDED/GRATED CHEESE|1.58|3|HT SHREDDED MOZZ/PROVLONE|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00072036705174|CHEESE|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|773cbb9738dc53c0072f5fcbd61f4e8cc7a8b0f0|3.0|2015-02-05 17:37:00|1.4132775322775095|3|7203632016|88|0.6126700657242101|0|58|195|-80.992182|30|35.103409|SALAD & COOKING OIL|0.0|1|HT VEGETABLE OIL|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00072036320223|SHORTENING/OIL|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|5205783636a9e093a53ebe491c3897dc2364f943|14.98|2014-10-25 21:26:00|1.4132775322775095|3|8500000748|88|0.6126700657242101|0|58|9983|-80.992182|889|35.103409|NFS-SPARKLING|0.0|13|CB-ANDRE EXTRA DRY|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00085000007488|SPARKLING|WINE|-80.992182|1.413580244274486|88|2
35.103409|9a93b08d6229206dd174929bbd71210949fec036|3.59|2014-09-16 23:23:00|80.992192682720116|3|7203695890|88|35.105739325068221|0|56|1654|-81.027334|381|34.977331|DESSERT CAKES|0.0|14|GRANDE FINALE CAKE SLICE|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|35.113093007298254|00072036958907|CAKES|BAKERY|-80.992182|80.99218618486077|149|1
35.103409|30929de313eea544e9df415caf8e8d6876bc7cb8|3.49|2015-02-11 22:34:00|1.4132775322775095|3|2840023981|88|0.6126700657242101|0|58|203|-80.992182|31|35.103409|CHEESE SNACKS|1.75|1|CHEETOS JUMBO PUFFS|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00028400239875|SNACKS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|06580e4c1343694a66aa255944dea5c2c2686418|3.49|2014-12-31 20:51:00|1.4132775322775095|3|7797508161|88|0.6126700657242101|0|58|204|-80.992182|31|35.103409|TORTILLA CHIPS|1.75|1|SNYDERS YLLW CRN TORTILLA CHP|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00077975081624|SNACKS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|6cf330a0b524532079c8741b46283c6588105cf9|1.1|2015-02-06 17:24:00|1.4132775322775095|3|5000000124|88|0.6126700657242101|0|58|154|-80.992182|24|35.103409|NFS-CAT FOOD WET|0.0|1|FANCY FEAST SEAFOOD FEAST|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00050000429349|PET FOOD/SUPPLIES|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|b391cc23a5a5da23fbf9b968401a479fc4dbbaa2|2.59|2015-02-04 17:37:00|1.4132775322775095|3|7203608135|88|0.6126700657242101|0|58|82|-80.992182|11|35.103409|VINEGAR|0.0|1|HT VINEGAR WHITE DISTILLED 128|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00072036081353|CONDIMENTS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|01be2e0fd58fa27e51e86b10b6954152c4f6486b|1.27|2015-02-01 10:18:00|1.4132775322775095|3|7203613030|88|0.6126700657242101|0|58|101|-80.992182|15|35.103409|FLOUR-ALL PURPOSE|0.0|1|HARRIS TEETER ALL PRPOSE FLOUR|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00072036130303|FLOUR|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|8bff63b7dc136e897bbe7e53cc528c37ec62f5ff|2.27|2014-11-27 11:46:00|1.4132775322775095|3|7203611029|88|0.6126700657242101|0|58|55|-80.992182|8|35.103409|REGULAR|0.0|23|HT ROOT BEER 12PK|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00072036110701|CARBONATED BEVERAGES|BEVERAGE|-80.992182|1.413580244274486|88|1
35.103409|95d9e5c7bacfaf6eb6d4fbf7ec1ccc83c8305335|20.7|2015-02-13 18:41:00|1.4132775322775095|3|4460030438|88|0.6126700657242101|0|58|730|-80.992182|24|35.103409|NFS-CAT LITTER|5.18|1|FRESH STEP EXTRM SCOOPABLE LIT|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00044600306223|PET FOOD/SUPPLIES|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|6cdf236fe6acf0f3923e5bf3bf206b7085359841|9.99|2014-09-21 01:03:00|80.992192682720116|3|7203661033|88|35.105739325068221|0|56|666|-81.027334|145|34.977331|PACKAGED COOKED|0.0|12|HT COOKED SHRIMP RING 10OZ|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|35.113093007298254|00072036610331|SHRIMP|SEAFOOD|-80.992182|80.99218618486077|149|1
35.103409|e44d3194e6d5454c87825cbd0ebeb01f48d44924|0.64|2015-01-25 18:27:00|1.4132775322775095|3||88|0.6126700657242101|0|58|542|-80.992182|64|35.103409|FRESH VEGETABLES REMAIN|0.0|4|COO SNOW PEAS, BULK|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00204092000003|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|1
35.103409|58fec6d046dccced926d4d916598870f71d05fa3|3.39|2015-01-25 11:24:00|1.4132775322775095|3|2100002782|88|0.6126700657242101|0|58|182|-80.992182|28|35.103409|MAYO|0.0|1|KRAFT SQZ MAYO CHIPOTLE|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00021000027828|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|58930adea3e91cded3c2d1da05191b30eab20a45|0.99|2015-02-03 20:52:00|1.4132775322775095|3|1780014597|88|0.6126700657242101|0|58|154|-80.992182|24|35.103409|NFS-CAT FOOD WET|0.0|1|ONE BRAISED CUTS TUNA N GRAVY|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00017800146098|PET FOOD/SUPPLIES|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|54446d9597eaaccfdbac25ae34b09a915c4f931c|4.65|2014-10-25 00:34:00|1.4132775322775095|3|7218063473|88|0.6126700657242101|0|58|254|-80.992182|892|35.103409|PREMIUM PIZZA|0.0|5|RED BARON PEPPERONI|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00072180634733|FROZEN PIZZA|FROZEN|-80.992182|1.413580244274486|88|1
35.103409|b04b8926259b893d6215a84b6ea6693010e1bb43|2.49|2015-02-12 17:26:00|1.4132775322775095|3|20488400000|88|0.6126700657242101|0|58|544|-80.992182|64|35.103409|FRESH PRODUCE FRSH HERBS|0.0|4|BUNCH THYME|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00033383801179|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|1
35.103409|f97493e3b1802a0bab641307ce110901114a278c|4.29|2014-09-24 19:51:00|1.4132775322775095|3|7203695667|88|0.6126700657242101|0|58|1693|-80.992182|385|35.103409|CROISSANTS|0.0|14|MINI BUTTER CROISSANTS|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00072036956675|SWEET GOODS|BAKERY|-80.992182|1.413580244274486|88|1
35.103409|261c4ffe4035975d861987c4e8db78bc3da86a76|2.19|2015-01-28 17:55:00|1.4132775322775095|3|4300028543|88|0.6126700657242101|0|58|28|-80.992182|26|35.103409|STUFFING PRODUCTS|0.0|1|STOVE TOP STUFFING CHICKEN|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00043000285213|PREPARED FOODS-DRY MIXES|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|ce2cf1a2ded7742730d1bfe90effe18aa7644ce3|8.99|2014-11-18 21:11:00|1.4132775322775095|3|8600300502|88|0.6126700657242101|0|58|9917|-80.992182|891|35.103409|NFS-OTHER WINE|0.0|13|REX GOLIATH PINOT NOIR 1.5L|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00086003005020|WINE REMAINING|WINE|-80.992182|1.413580244274486|88|1
35.103409|441a329893426c23a4d678cf818cf6124f4c1767|9.99|2014-12-26 23:01:00|1.4132775322775095|3|8600300502|88|0.6126700657242101|0|58|9917|-80.992182|891|35.103409|NFS-OTHER WINE|0.0|13|REX GOLIATH PINOT NOIR 1.5L|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00086003005020|WINE REMAINING|WINE|-80.992182|1.413580244274486|88|1
35.103409|2a7e8dddcacafdafb219fb1aa0ca55f1f21f464c|2.29|2014-11-13 22:49:00|1.4132775322775095|3|7800023046|88|0.6126700657242101|0|58|55|-80.992182|8|35.103409|REGULAR|1.29|23|CANADA DRY CBRY G/ALE 2LTR|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00078000156461|CARBONATED BEVERAGES|BEVERAGE|-80.992182|1.413580244274486|88|1
35.103409|b7b8597ec194d7ad5b2cace263a6460249e785ae|12.99|2014-09-21 21:10:00|1.4132775322775095|3|7199009516|88|0.6126700657242101|0|58|458|-80.992182|82|35.103409|CRAFT BEER|0.0|16|BLUE MOON BELGIAN 12PK|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00071990095161|DOMESTIC BEER|BEER|-80.992182|1.413580244274486|88|1
35.103409|d699aa4a641efaa5f52a2f472104222d3a44ceb6|3.99|2014-12-08 19:13:00|1.4132775322775095|3|89504500027|88|0.6126700657242101|0|58|3177|-80.992182|1010|35.103409|MAKE UP REMOVER|0.0|17|EYE & MU REMVR TOWELETTES-REF|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00895045000272|NAIL CARE|HBC|-80.992182|1.413580244274486|88|1
35.103409|6c068cf5623d8957c0ce6be59cc1cd02a7b13e54|5.99|2014-09-11 16:53:00|1.4132775322775095|3|8143403123|88|0.6126700657242101|0|58|9934|-80.992182|885|35.103409|NFS POP CHARDONNAY|0.0|13|CB-REX GOLIATH CHARDONNAY|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00081434031235|POPULAR (4-$7.99)|WINE|-80.992182|1.413580244274486|88|1
35.103409|36a37a9353900e249c5fa0bf1c5451c478617d88|7.79|2015-01-13 21:57:00|1.4132775322775095|3|5400036413|88|0.6126700657242101|0|58|427|-80.992182|72|35.103409|NFS-TOILET TISSUE|0.0|1|SCOTT BATH SOFT 12 RL|6f703643b45c6c3522e05c5fcec8fb7f9d7befae|0.16102000845921496|0.61177642288969325|00054000364136|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.06858|b282105c5ca796fff865edc222ba2249dfed2776|4.29|2014-10-09 15:41:00|1.4091206135396188|3|2840006399|273|0.612062184999033|0|47|204|-80.7007|31|35.06858|TORTILLA CHIPS|0.29|1|TOSTITOS BITES|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00028400064057|SNACKS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|44a690aebaa456759e22387d9067bd3acc1086b3|11.98|2014-10-30 14:20:00|1.4091206135396188|3|7403008182|273|0.612062184999033|0|47|2017|-80.7007|505|35.06858|STRETCHED CURD CHEESE|2.99|6|SORRENTO FRESH MOZZARELLA|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00074030081827|SPECIALTY CHEESE|DELI|-80.7007|1.4084929236641879|273|2
35.06858|b2531ae30fee1b6de2fae8c9d1a1cd4bef33e447|6.78|2015-02-10 18:07:00|1.4091206135396188|3|7247010043|273|0.612062184999033|0|47|1641|-80.7007|377|35.06858|PACKAGED DONUTS|0.0|14|KK GLAZED MINI PIES-CHERRY 6PK|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00072470100436|DONUTS|BAKERY|-80.7007|1.4084929236641879|273|2
35.06858|32dd12b0dad5677f5f21fe4e66dee9310b0b899d|3.29|2015-01-25 13:10:00|1.4091206135396188|3|7225091171|273|0.612062184999033|0|47|1033|-80.7007|163|35.06858|HAMBURGER|0.0|7|NATOWN WHITEWHEAT HAMS|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00072250911719|BUNS/ROLLS|COMMERCIAL BAKERY|-80.7007|1.4084929236641879|273|1
35.06858|f0d368707883a9769d37afec6901071d48f48a91|5.99|2014-10-06 16:31:00|1.4091206135396188|3|7203688103|273|0.612062184999033|0|47|562|-80.7007|64|35.06858|FRESH CUT FRUIT|0.0|4|HT WATERMELON CHUNKS 32OZ|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00072036881038|FRESH PRODUCE|PRODUCE|-80.7007|1.4084929236641879|273|1
35.06858|aa18aa037b410e9ea223feaaae1be0c46aa0c14d|19.99|2014-12-16 12:57:00|80.700712769248256|3|7203695593|273|35.092106347882151|0|42|1653|-80.80146|381|35.17739|CELEBRATION CAKES|0.0|14|1/4 DL CHOC CK W WH BUTTRCRM|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|35.088667338853092|00072036955937|CAKES|BAKERY|-80.7007|80.700719457594474|208|1
35.06858|65338efa2b8421fc83dc96f5f829802fecb57595|5.99|2015-02-14 17:41:00|1.4091206135396188|3|7203688103|273|0.612062184999033|0|47|562|-80.7007|64|35.06858|FRESH CUT FRUIT|0.0|4|HT WATERMELON CHUNKS 32OZ|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00072036881038|FRESH PRODUCE|PRODUCE|-80.7007|1.4084929236641879|273|1
35.06858|3edef38c75c0171e38f179fa1ded8553d9874b4a|1.37|2014-12-03 18:29:00|1.4091206135396188|3|7203625014|273|0.612062184999033|0|47|145|-80.7007|22|35.06858|MILK-CANNED|0.0|1|HT SWEETENED CONDENSED MILK|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00072036250148|PACKAGED MILKS & MODIFIERS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|3e26f511d439f6452d950540e9d6f3af099295e4|6.69|2014-12-01 18:59:00|1.4091206135396188|3|7203618986|273|0.612062184999033|0|47|8433|-80.7007|1769|35.06858|ALKALINE AA|0.0|18|(FE)(JHK) HT AA BATTERIES|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00072036189868|BATTERY & FLASHLIGHT|GM|-80.7007|1.4084929236641879|273|1
35.06858|51c9f87d7dadd4d192072543e753afc83f094e41|4.98|2015-03-09 11:57:00|80.700712769248256|3|5040073942|273|35.092106347882151|0|42|1033|-80.80146|163|35.17739|HAMBURGER|0.0|7|BALL PARK WHITE HAMS 8PK PP|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|35.088667338853092|00050400739420|BUNS/ROLLS|COMMERCIAL BAKERY|-80.7007|80.700719457594474|208|2
35.06858|bd24a7e71ea0d1f992f3ef8c56f3f98bea1347b5|1.99|2014-10-10 16:31:00|80.700712769248256|3|3900004504|273|35.092106349736511|0|42|114|-80.709466|14|35.124987|PUMPKIN|0.0|1|LIBBY SOLID PACK PUMPKIN|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|35.088667338853092|00039000045049|DESSERTS/GELS/SYRUPS|G1 GROCERY|-80.7007|80.700715757861701|157|1
35.06858|f1ddc408054ecca39290136eae81ccd1f2a0326a|1.69|2014-12-02 16:43:00|1.4091206135396188|3|7203688003|273|0.612062184999033|0|47|527|-80.7007|64|35.06858|FRESH CARROTS|0.0|4|HT BABY CARROTS 1LB BAG|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00072036880031|FRESH PRODUCE|PRODUCE|-80.7007|1.4084929236641879|273|1
35.06858|3bde0592718bac2a5616d74013d193cc0aa92abf|26.76|2014-11-16 12:58:00|1.4091206135396188|3|20007200000|273|0.612062184999033|0|47|975|-80.7007|201|35.06858|POULTRY-FROZEN|10.1|2|16 X 20 H T PREMIUM TURKEY|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00200072000001|POULTRY|MEAT|-80.7007|1.4084929236641879|273|1
35.06858|671d0b48143dd93456f9e8bc8b65fb8e3914c455|3.29|2015-01-09 11:20:00|1.4091206135396188|3|2265530301|273|0.612062184999033|0|47|483|-80.7007|100|35.06858|TURKEY BACON|0.5|19|BBALL LOW SODIUM TURKEY BACON|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00022655300441|BACON|CASE READY MEATS|-80.7007|1.4084929236641879|273|1
35.06858|c9f386e574d201f195f0705d2ba13ad46426f043|3.29|2015-02-06 18:45:00|1.4091206135396188|3|2265530301|273|0.612062184999033|0|47|483|-80.7007|100|35.06858|TURKEY BACON|0.79|19|BUTTERBALL TURKEY BACON|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00022655303015|BACON|CASE READY MEATS|-80.7007|1.4084929236641879|273|1
35.06858|f2fbc1a6cbf53f27e11c9cb90b38ef907b10aec2|1.29|2015-02-20 12:33:00|1.4091206135396188|3|2880014315|273|0.612062184999033|0|47|242|-80.7007|39|35.06858|CANNED BEANS|0.29|1|HANOVER PEAS CHICK|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00028800159018|VEGETABLES-CAN/JAR|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|e2c89f522806f104bc3850fb2b151d738c8b4f95|1.79|2014-09-18 17:16:00|80.700712769248256|3|7339000393|273|35.092106349736511|0|42|48|-80.709466|7|35.124987|REGISTER GUM|0.0|1|MENTOS FRESH MINT GUM 15CT|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|35.088667338853092|00073390013936|CANDY|G1 GROCERY|-80.7007|80.700715757861701|157|1
35.06858|2e2ca735f7d5f60017e9620797d477d979b33e4c|2.49|2014-11-13 16:44:00|80.700712769248256|3|4133112001|273|35.092106353268306|0|42|1214|-80.64817|272|35.04711|AUTHENTIC HISPANIC|0.0|1|GOYA PEAS PIGEON|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|35.088667338853092|00041331120012|HISPANIC PREP. FOODS|G1 GROCERY|-80.7007|80.70070040694111|129|1
35.06858|4fa42b32633ee06b176faf7ebb7597572a4d408f|1.35|2014-10-13 17:24:00|1.4091206135396188|3|1530043023|273|0.612062184999033|0|47|238|-80.7007|38|35.06858|RICE FLAVORED|0.0|1|RICE A RONI RICE PILAF|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00015300430594|RICE GRAINS AND BEANS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|d31f2daf8e84d7ab29e8d0b77fe6ca22dbe09ac9|2.79|2015-02-13 21:16:00|1.4091206135396188|3|1800000501|273|0.612062184999033|0|47|328|-80.7007|54|35.06858|SWEET ROLLS-REFRIGERATED|0.0|3|PILLSBURY REDUCED FAT CINNAMON|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00018000005093|DOUGH PRODUCTS|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|9d47f263a64aac43486d7387791f7a946a4f986b|5.79|2015-02-24 18:06:00|1.4091206135396188|3|7247000603|273|0.612062184999033|0|47|1641|-80.7007|377|35.06858|PACKAGED DONUTS|0.0|14|K K 12 CT GLAZED DONUTS PP|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00072470006035|DONUTS|BAKERY|-80.7007|1.4084929236641879|273|1
35.06858|0ff5439e79f787c24126fa1e4e77e0adcb9e09bb|2.99|2015-02-07 12:43:00|1.4091206135396188|3|7433610102|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HIGHLAND CREST 2% REDUCE FAT|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00074336101021|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|bff9d48bbd2f23944de24f31164802cdf845ffdb|7.5|2014-09-13 21:32:00|80.700712769248256|3|7433610102|273|35.092106347340014|0|42|342|-80.699686|57|35.000049|FRESH MILK|0.0|3|HIGHLAND CREST 2% REDUCE FAT|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|35.088667338853092|00074336101021|MILK|DAIRY|-80.7007|80.700720412959697|249|2
35.06858|fe77569a242a50fe0bc0274d8d66a2af3c5a6d0a|2.69|2015-01-11 13:02:00|1.4091206135396188|3|7203698126|273|0.612062184999033|0|47|1132|-80.7007|55|35.06858|EGGS SUBSTITUTES|0.0|3|HARRIS TEETER LIQUID EGG WHITE|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00072036981264|EGGS FRESH|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|c9a8a7f7272bba21dbc651019bcfe75724770ffe|2.69|2015-01-15 15:39:00|1.4091206135396188|3|7225001739|273|0.612062184999033|0|47|1025|-80.7007|162|35.06858|WHITE|0.0|7|NATOWN WHITEWHEAT RTOP BRD|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00072250017398|SLICED BREAD|COMMERCIAL BAKERY|-80.7007|1.4084929236641879|273|1
35.06858|735fd4976d16f8ed36fe1462a3b04c6d8d1f1ae5|7.98|2014-12-23 15:58:00|80.700712769248256|3|7203663995|273|35.092106347882151|0|42|342|-80.80146|57|35.17739|FRESH MILK|0.0|3|HARRIS TEETER 1% MILK|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|35.088667338853092|00072036631275|MILK|DAIRY|-80.7007|80.700719457594474|208|2
35.06858|613ff579a8aafec6369c3b7620263e9d22c6bb6f|3.99|2014-09-18 17:48:00|1.4091206135396188|3|7203663995|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HARRIS TEETER 1% MILK|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00072036631275|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|2b5856bb1e9ea30869286f5c20f570cffc5e2b00|7.98|2014-10-17 18:35:00|1.4091206135396188|3|7203663995|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HARRIS TEETER 1% MILK|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00072036631275|MILK|DAIRY|-80.7007|1.4084929236641879|273|2
35.06858|d1e125b0b616bca41eb504eda973aba27d19989f|3.99|2014-10-15 20:55:00|1.4091206135396188|3|7203663995|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HARRIS TEETER 1% MILK|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00072036631275|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|eab20d8f03e7c0494730253526b7ff8733b3e25b|2.29|2014-09-19 19:53:00|1.4091206135396188|3|1800000260|273|0.612062184999033|0|47|325|-80.7007|54|35.06858|BISCUITS-REFRIGERATED|0.0|3|GRANDS BUTTERMILK BISCUITS|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00018000001828|DOUGH PRODUCTS|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|874f794f731154ffc72cc1aead0a606f148f3242|3.49|2014-11-12 19:42:00|1.4091206135396188|3|3800039118|273|0.612062184999033|0|47|81|-80.7007|9|35.06858|RTE CEREAL KIDS|0.99|1|KELLOGG FROOT LOOPS 12.2|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00038000391187|CEREAL|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|3ac2ca5218f2d876172131203d740d15ca19ed67|7.98|2015-02-16 14:56:00|1.4091206135396188|3|7430500116|273|0.612062184999033|0|47|82|-80.7007|11|35.06858|VINEGAR|0.0|1|BRAGG ORG VINEGAR APPLE CIDER|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00074305001161|CONDIMENTS|G1 GROCERY|-80.7007|1.4084929236641879|273|2
35.06858|4b5c15742dacaf2839c5f4b3179d42084457df94|4.85|2014-12-06 14:39:00|80.700712769248256|3|3450015136|273|35.092106347340014|0|42|312|-80.699686|51|35.000049|BUTTER|0.0|3|L O L UNSALTED BUTTER QUARTERS|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|35.088667338853092|00034500151504|BUTTER & MARGARINE|DAIRY|-80.7007|80.700720412959697|249|1
35.06858|85c04ee8bceb9fb61e591016f20afa64363b8619|2.79|2015-01-26 16:14:00|1.4091206135396188|3|1600043776|273|0.612062184999033|0|47|24|-80.7007|3|35.06858|FROSTING-READY-TO-SPREAD|0.0|1|BC HRSHY MLK CHOC FROSTING|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00016000437760|BAKING SUPPLIES|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|a444b435c607b0a7713992e072f6cbb5d7dd8bf8|1.99|2014-09-28 18:03:00|80.700712769248256|3|7203648011|273|35.092106347340014|0|42|274|-80.699686|44|35.000049|ICE|0.0|5|HT BAGGED ICE 10LB (456)|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|35.088667338853092|00000000004560|ICE|FROZEN|-80.7007|80.700720412959697|249|1
35.06858|678532e28b13ca197943f006164ebf843bf87e0e|1.99|2014-11-17 17:17:00|1.4091206135396188|3|7203648011|273|0.612062184999033|0|47|274|-80.7007|44|35.06858|ICE|0.0|5|HT BAGGED ICE 10LB (456)|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00000000004560|ICE|FROZEN|-80.7007|1.4084929236641879|273|1
35.06858|5625ee80d31c84c0fe0e0676dd098b97c41af28f|1.99|2014-11-08 16:12:00|1.4091206135396188|3|7203648011|273|0.612062184999033|0|47|274|-80.7007|44|35.06858|ICE|0.0|5|HT BAGGED ICE 10LB (456)|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00000000004560|ICE|FROZEN|-80.7007|1.4084929236641879|273|1
35.06858|6de3766a4986c8342db19894f4ef36c3e51786e9|3.99|2015-01-10 16:01:00|1.4091206135396188|3|7433610006|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HUNTER 1%  MILK  GALLON|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00074336100291|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|abd34cdcca43195901d5a5326d6cb83470bdb7ec|4.29|2015-01-16 16:15:00|1.4091206135396188|3|7203670353|273|0.612062184999033|0|47|442|-80.7007|76|35.06858|NFS-COOKING-STORAGE BAGS|0.79|1|YH RESEAL DBL ZIP STORAGE GAL|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00072036703545|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|09f1ed7802c4b97856c2fa5b88ca2555d263b091|2.5|2014-12-21 12:49:00|80.700712769248256|3|78142100610|273|35.092106349270338|0|42|1601|-80.739|371|35.141204|BRANDED BREAD|0.0|14|LA BREA FRENCH BAGUETTE|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|35.088667338853092|00781421006108|BREAD|BAKERY|-80.7007|80.700716764981351|171|1
35.06858|3f9d5e594cb71e52a6361b288d8b1ea6644137b1|3.29|2014-10-10 17:51:00|1.4091206135396188|3|71514150349|273|0.612062184999033|0|47|330|-80.7007|55|35.06858|EGGS|0.0|3|EGGLAND BEST GRADE A LARGE EGG|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00715141503494|EGGS FRESH|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|3d70328af4847a0419f607098ff53a25ab58ab60|7.29|2014-10-11 17:56:00|1.4091206135396188|3|1780013465|273|0.612062184999033|0|47|156|-80.7007|24|35.06858|NFS-DOG FOOD-DRY|0.8|1|BENEFUL INCREDIBITES|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00017800136402|PET FOOD/SUPPLIES|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|b0b2a264e3792d8dce49b27c2eaf4cf81b964b25|2.19|2014-11-28 16:43:00|1.4091206135396188|3|1200000230|273|0.612062184999033|0|47|55|-80.7007|8|35.06858|REGULAR|0.2|23|DR PEPPER 2 LITER|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00078000082463|CARBONATED BEVERAGES|BEVERAGE|-80.7007|1.4084929236641879|273|1
35.06858|909a7419b1110d33e659bfd56056b452ff6ac132|9.49|2014-12-11 17:23:00|1.4091206135396188|3|3680021544|273|0.612062184999033|0|47|4379|-80.7007|1210|35.06858|ACID BLOCKER-SWALLOW|0.0|17|TC OMEPRAZOLE ACID REDUCER|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|0.61242566243833529|00036800215443|STOMACH REMEDIES|HBC|-80.7007|1.4084929236641879|273|1
35.06858|bd29fa250655e76317aaef35ba3043a24d0e1e35|9.63|2015-01-29 16:38:00|80.700712769248256|3|20894800000|273|35.092106348840751|0|42|977|-80.816172|201|35.059823|FRESH HT CHICKEN|0.0|2|HT FRESH CUT-UP CHICKEN|74c2c4dd089708706b78b990793e5858455561ae|1.6256141968941031|35.088667338853092|00208948000001|POULTRY|MEAT|-80.7007|80.700717642194732|66|1
35.297134|ede70d473cf2f51e838a22b13e7a7ccd0c195cf2|1.99|2015-03-05 09:14:00|80.737901233649083|2|71146450634|258|35.346914866494124|0|46|79|-80.810056|273|35.219587|ASIAN SAUCES/SEASONINGS|1.0|1|BLUE DRAGON SC HNY TERIYAKI|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00711464506242|ASIAN PREP. FOODS|G1 GROCERY|-80.737839|80.737908221770127|401|1
35.297134|cc12a27f8c2b66188ca78c7fe1cf7f9e71200c2d|10.76|2014-12-31 07:11:00|80.737901233649083|2|70935100013|258|35.346914866494124|0|46|556|-80.810056|64|35.219587|PACKAGED VEGETABLES|0.0|4|APIO BROCCOLI FLORETS|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00709351000133|FRESH PRODUCE|PRODUCE|-80.737839|80.737908221770127|401|4
35.297134|bc3a397f5d3f813a87754190cf9ef25fe9475b84|6.58|2014-11-16 16:16:00|80.737901233649083|2|1204403891|258|35.34691489783858|0|46|3876|-80.66939|1070|35.28326|SOLID-MALE|0.8|17|OLD SPICE HI ENDURNC STCK ORIG|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00012044038888|DEODORANT|HBC|-80.737839|80.737849194022729|46|2
35.297134|d91bc3b1351b8a16ba94e6e65e754c7a3b0b32b2|1.39|2014-10-13 17:33:00|80.737901233649083|2|4920005675|258|35.34691489783858|0|46|224|-80.66939|35|35.28326|SUGAR-BROWN|0.4|1|DOMINO LT BRWN SUGAR-BOX|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00049200056752|SUGAR/SUBSTITUTES|G1 GROCERY|-80.737839|80.737849194022729|46|1
35.297134|5551d3d68f7c675a7bbf290c11cc2c5f16db4a07|2.89|2014-10-26 18:51:00|1.4094857484078087|2|7203697887|258|0.6160512048176361|0|26|61|-80.737839|9|35.297134|RTE CEREAL ADULT|0.92|1|HT CER BRAN FLAKES|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|0.61471665291522548|00072036060174|CEREAL|G1 GROCERY|-80.737839|1.409141121495086|258|1
35.297134|3c3b99150575db9136bd4f8e06b1acb618872d57|4.98|2014-12-17 08:39:00|80.737901233649083|2|3080000920|258|35.346914866494124|0|46|727|-80.810056|7|35.219587|SEASONAL CANDY-SINGLE FAC|0.98|1|I/O(C15)SPNGLR MINI CANES|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00030800009200|CANDY|G1 GROCERY|-80.737839|80.737908221770127|401|2
35.297134|662f94494d1c6c422940c0dd8648879fcf53c68a|22.3|2014-11-22 10:47:00|80.737901233649083|2|20092500000|258|35.34691489783858|0|46|974|-80.66939|201|35.28326|FRESH TURKEY|5.59|2|ALL NATURAL FRESH DUCK|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00200925000004|POULTRY|MEAT|-80.737839|80.737849194022729|46|1
35.297134|5ccdbc786eb8cc2cc468fbc6d61adaa2bfeda4c0|26.369999999999997|2015-02-18 18:25:00|1.4094857484078087|2|7274580677|258|0.6160512048176361|0|26|353|-80.737839|110|35.297134|FROZEN CASE MEAT|4.4|19|PERDUE SIMPLY SMART GF NUGGETS|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|0.61471665291522548|00072745805776|FROZEN CASE MEAT|CASE READY MEATS|-80.737839|1.409141121495086|258|3
35.297134|5f36ceb0ad56b2543c05fb8e27d213b5f13ec38c|2.65|2015-01-08 13:39:00|80.737901233649083|2|4119601000|258|35.34691489783858|0|46|1201|-80.66939|33|35.28326|RTS CANNED|2.65|1|PROG TRAD CHICKEN ROTINI|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00041196910582|SOUP|G1 GROCERY|-80.737839|80.737849194022729|46|1
35.297134|6f2e4d96e7345fb3ec5b11ca85c90f8edfcb8856|1.89|2015-02-12 08:14:00|80.737901233649083|2|4010000928|258|35.346914866494124|0|46|29|-80.810056|3|35.219587|REMAINING BAKING SUPPLIES|0.0|1|FLEISCHMAN YEAST PACKETS|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00040100009282|BAKING SUPPLIES|G1 GROCERY|-80.737839|80.737908221770127|401|1
35.297134|24bbde92297665747016bcc320849493a329ba5e|2.65|2015-01-07 19:06:00|1.4094857484078087|2|4119601000|258|0.6160512048176361|0|26|1201|-80.737839|33|35.297134|RTS CANNED|0.0|1|PROG TRAD CHICKEN ROTINI|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|0.61471665291522548|00041196910582|SOUP|G1 GROCERY|-80.737839|1.409141121495086|258|1
35.297134|55fe7b1151f9928d43fc917f2737496a6dc26f36|3.39|2014-10-16 10:56:00|80.737901233649083|2|4450034122|258|35.34691489783858|0|46|357|-80.66939|104|35.28326|SMOKED SAUSAGE ROPES|0.0|19|HILLSHIRE TURKEY SMOKED SAUSAG|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00044500341157|DINNER SAUSAGE|CASE READY MEATS|-80.737839|80.737849194022729|46|1
35.297134|59aea76d2fd9b9aee3522fa1a1f775967ec3e66d|2.0|2014-11-23 17:25:00|80.737901233649083|2|4300000953|258|35.34691489783858|0|46|272|-80.66939|307|35.28326|TOPPINGS FROZEN|1.01|5|COOL WHIP WHIPPED TOPPING|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00043000009536|DESSERTS FROZEN|FROZEN|-80.737839|80.737849194022729|46|1
35.297134|fb39caeb73290cef08c5c453ced4a06166a30a57|6.49|2015-01-18 16:08:00|80.737901233649083|2|85281048912|258|35.34691489783858|0|46|364|-80.66939|55|35.28326|ORGANIC AND CF EGGS|0.0|3|LOL CAGE FREE A LRG BRWN EGGS|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00852810489120|EGGS FRESH|DAIRY|-80.737839|80.737849194022729|46|2
35.297134|b822ad299b30c8024e6ac062218ac3154f2c5973|10.99|2014-11-25 08:27:00|80.737901233649083|2|85139000300|258|35.346914866494124|0|46|9957|-80.810056|886|35.219587|NFS-PREM-OTHER RED|0.0|13|EPPA SANGRIA RED|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00851390003009|PREMIUM ($8-$10.99)|WINE|-80.737839|80.737908221770127|401|1
35.297134|89e377b2d4f0d1a1c135f099f5e1b2da6612ded1|3.69|2015-02-12 16:43:00|80.737901233649083|2|7373100830|258|35.34691489783858|0|46|495|-80.66939|108|35.28326|NON REFRIGERATED|1.2|19|MISSION FAJITA TORTILLA 20 CT|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00073731008300|TORTILLAS|CASE READY MEATS|-80.737839|80.737849194022729|46|1
35.297134|c2d74441aa2021d2deae73e347f6681769fe91ae|2.19|2015-02-20 17:16:00|80.737901233649083|2|7910000367|258|35.346914866494124|0|46|154|-80.810056|24|35.219587|NFS-CAT FOOD WET|0.0|1|9LIVES LIVER & CHICKEN 4PK|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00079100003129|PET FOOD/SUPPLIES|G1 GROCERY|-80.737839|80.737908221770127|401|1
35.297134|9a7875c1ce76012e104fbd9ac3861168a9c23dbe|5.97|2014-10-18 16:43:00|1.4094857484078087|2|7910000367|258|0.6160512048176361|0|26|154|-80.737839|24|35.297134|NFS-CAT FOOD WET|0.98|1|9LIVES LIVER & CHICKEN 4PK|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|0.61471665291522548|00079100003129|PET FOOD/SUPPLIES|G1 GROCERY|-80.737839|1.409141121495086|258|3
35.297134|5343d8f266e941389a3ab19326ce102cfbb0499f|7.78|2015-03-02 13:13:00|80.737901233649083|2|7332100018|258|35.346914866494124|0|46|1277|-80.810056|279|35.219587|FROZEN SNACKS|0.0|5|SUPERPRETZEL SOFT PRETZELS|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00073321000189|FROZEN SANDWICH AND SNACKS|FROZEN|-80.737839|80.737908221770127|401|2
35.297134|56bf51b80e9171274b07d6d6d058be851d002ad2|15.99|2015-02-23 17:22:00|1.4094857484078087|2|7203696987|258|0.6160512048176361|0|26|751|-80.737839|87|35.297134|NFS-BOUQUETS|0.0|9|15.99 SUNFLOWER BQT|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|0.61471665291522548|00072036969873|FLORAL|FLORAL|-80.737839|1.409141121495086|258|1
35.297134|7fcdf2e2521a162c859d061d1a62ef6cd0bc8f75|2.99|2014-12-07 18:36:00|1.4094857484078087|2|9396600091|258|0.6160512048176361|0|26|345|-80.737839|57|35.297134|ORGANIC MILK|0.0|3|ORGANIC VALLEY WHOLE MILK|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|0.61471665291522548|00093966000917|MILK|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|af53eaeea1a08e29e381232eab6ed98a75ee2934|4.99|2015-02-04 17:58:00|1.4094857484078087|2|2100061526|258|0.6160512048176361|0|26|315|-80.737839|52|35.297134|CHEESE-PROCESSED-SLICED|1.0|3|KRAFT SINGLE WRAP CHS|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|0.61471665291522548|00021000615261|CHEESE|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|9299c4fec2c1a5051bccf156b118a9ab7cdbf4c3|3.29|2015-01-12 16:27:00|80.737901233649083|2|2265530301|258|35.34691489783858|0|46|483|-80.66939|100|35.28326|TURKEY BACON|0.5|19|BBALL LOW SODIUM TURKEY BACON|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00022655300441|BACON|CASE READY MEATS|-80.737839|80.737849194022729|46|1
35.297134|fd7d23ce743795f20013a71bba5f34778478fc84|5.98|2014-12-02 18:56:00|1.4094857484078087|2|20424200000|258|0.6160512048176361|0|26|512|-80.737839|64|35.297134|FRSH PROD FRSH FRUIT REM|0.0|4|CRANBERRIES 12 OZ|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|0.61471665291522548|00038900071769|FRESH PRODUCE|PRODUCE|-80.737839|1.409141121495086|258|2
35.297134|bc0bbd0ef75ae3c3ec87b6d37d6703af36de9540|3.94|2014-12-24 15:30:00|1.4094857484078087|2|7203614993|258|0.6160512048176361|0|26|105|-80.737839|16|35.297134|FRUIT CUPS AND GELS|0.0|1|HT 4PK FRT CUP MANDARIN|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|0.61471665291522548|00072036980564|FRUIT-CAN/JAR|G1 GROCERY|-80.737839|1.409141121495086|258|2
35.297134|8063f07b00584d1b6836742bdbc1641e2a810937|3.99|2015-03-02 09:01:00|80.737901233649083|2|4973309101|258|35.346914866494124|0|46|76|-80.810056|11|35.219587|MEAT SAUCES|0.0|1|CHOLULA HOT SC CHILI LIME|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00049733840118|CONDIMENTS|G1 GROCERY|-80.737839|80.737908221770127|401|1
35.297134|9c9797340dfc51e13f30095e22e6fa0d9adff2d6|3.99|2014-10-06 08:13:00|80.737901233649083|2|4973309101|258|35.346914866494124|0|46|76|-80.810056|11|35.219587|MEAT SAUCES|1.0|1|ECHOLULA CHIPOTLE SAUCE|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00049733830119|CONDIMENTS|G1 GROCERY|-80.737839|80.737908221770127|401|1
35.297134|4e20a48a0dd6d49fc7d5af447aa3ec2d5dbbb43e|5.3|2014-10-26 18:49:00|1.4094857484078087|2|5150000094|258|0.6160512048176361|0|26|126|-80.737839|19|35.297134|PRESERVES/MARMALADE|0.0|1|D SMUCKER BLUEBERRY PRESERVES|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|0.61471665291522548|00051500000793|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.737839|1.409141121495086|258|2
35.297134|dd910a3dd2e75c3545f2dbe5a3fc7c1f7be6018e|0.99|2014-10-23 18:31:00|1.4094857484078087|2|7203698291|258|0.6160512048176361|0|26|245|-80.737839|39|35.297134|VEGETABLES-CORE|0.39|1|HT CORN WK GOLDEN|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|0.61471665291522548|00072036411815|VEGETABLES-CAN/JAR|G1 GROCERY|-80.737839|1.409141121495086|258|1
35.297134|215a861b2abcd6dc0b5e75386572f893c23d90d8|2.85|2015-01-11 15:28:00|80.737901233649083|2|4133500053|258|35.34691489783858|0|46|184|-80.66939|28|35.28326|SALAD DRESSINGS-LIQUID|1.43|1|KENS DRS LT APPLE CIDER|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00041335356219|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.737839|80.737849194022729|46|1
35.297134|781f1a308e2b25b9820b985625beb9bc2ecbff1c|11.94|2014-11-25 08:27:00|80.737901233649083|2|3900004504|258|35.346914866494124|0|46|114|-80.810056|14|35.219587|PUMPKIN|0.2|1|LIBBY SOLID PACK PUMPKIN|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00039000045049|DESSERTS/GELS/SYRUPS|G1 GROCERY|-80.737839|80.737908221770127|401|6
35.297134|7e7c388c9d1614555fd0809f5c463e1f0c8a48a8|0.99|2014-09-15 19:47:00|80.737901233649083|2|7203698291|258|35.34691489783858|0|46|245|-80.66939|39|35.28326|VEGETABLES-CORE|0.22|1|HT GREEN BEANS CUT|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00072036982919|VEGETABLES-CAN/JAR|G1 GROCERY|-80.737839|80.737849194022729|46|1
35.297134|d01930c2d40e351fc2f56252f711cad8b540f531|14.99|2014-12-31 17:13:00|1.4094857484078087|2|84323700815|258|0.6160512048176361|0|26|670|-80.737839|146|35.297134|CRAB PACKAGED|0.0|12|CHICKEN OF THE SEA CLAW CRAB|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|0.61471665291522548|00843237008155|CRAB|SEAFOOD|-80.737839|1.409141121495086|258|1
35.297134|60a2d15d78099d9b23d6bf60979eff429994f8b7|4.49|2014-12-07 18:39:00|1.4094857484078087|2|7203695755|258|0.6160512048176361|0|26|1647|-80.737839|379|35.297134|PACKAGED MUFFINS|0.0|14|12CT MINI BLUEBERRY MUFFINS|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|0.61471665291522548|00072036957559|MUFFINS|BAKERY|-80.737839|1.409141121495086|258|1
35.297134|47fd293b45045ac4014cd88e13ceb95f6c7104a5|3.99|2014-12-02 18:55:00|1.4094857484078087|2|7203663995|258|0.6160512048176361|0|26|342|-80.737839|57|35.297134|FRESH MILK|1.52|3|HARRIS TEETER FF SKIM MILK|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|0.61471665291522548|00072036631282|MILK|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|7657d142b907476066d4b92e948678b90f40bdbd|2.49|2014-10-26 10:45:00|80.737901233649083|2||258|35.34691489783858|0|46|500|-80.66939|64|35.28326|FRESH APPLES|0.0|4|BRAEBURN APPLES|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00204103000008|FRESH PRODUCE|PRODUCE|-80.737839|80.737849194022729|46|1
35.297134|eb99aef9f69f4e88852a977379372dc67bef31ae|8.0|2014-10-23 09:11:00|80.737901233649083|2||258|35.346914866494124|0|46|511|-80.810056|64|35.219587|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00204770000004|FRESH PRODUCE|PRODUCE|-80.737839|80.737908221770127|401|4
35.297134|66c19bff15b534be2f3d42b953ed3ef2e24b14be|3.34|2014-12-28 11:12:00|80.737901233649083|2|7203657050|258|35.346914866494124|0|46|687|-80.810056|61|35.219587|BLENDED|0.0|3|HT VANILLA NONFAT YOGURT|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00072036570512|YOGURT|DAIRY|-80.737839|80.737908221770127|401|2
35.297134|2664feaf16fc5f91523486486727cf187c17be4f|2.99|2015-02-03 17:27:00|80.737901233649083|2|5100015339|258|35.346914866494124|0|46|137|-80.810056|20|35.219587|TOMATO & VEGETABLE JUICE|1.0|1|V8 VFUSION PINEAPPLE STRAWBRY|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00051000206442|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.737839|80.737908221770127|401|1
35.297134|2da23b4deb61029c4cd6f903e1b1df6846fe37d0|3.99|2015-01-28 07:33:00|80.737901233649083|2|4973309101|258|35.346914866494124|0|46|76|-80.810056|11|35.219587|MEAT SAUCES|0.0|1|ECHOLULA HOT SAUCE 5|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00049733091015|CONDIMENTS|G1 GROCERY|-80.737839|80.737908221770127|401|1
35.297134|4f3a04cd00bcf1027e1dfd8474082ee3fe312013|3.99|2015-02-11 08:58:00|80.737901233649083|2|4973309101|258|35.346914866494124|0|46|76|-80.810056|11|35.219587|MEAT SAUCES|0.0|1|ECHOLULA HOT SAUCE 5|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00049733091015|CONDIMENTS|G1 GROCERY|-80.737839|80.737908221770127|401|1
35.297134|7d4691209d5153e7144686732ed027987ec44f12|7.98|2014-10-09 08:42:00|80.737901233649083|2|4973309101|258|35.346914866494124|0|46|76|-80.810056|11|35.219587|MEAT SAUCES|2.0|1|ECHOLULA HOT SAUCE 5|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00049733091015|CONDIMENTS|G1 GROCERY|-80.737839|80.737908221770127|401|2
35.297134|b779a34a2d2b47df041b0e90ba39e4922b5252be|2.99|2014-10-10 08:23:00|80.737901233649083|2|4142074425|258|35.346914866494124|0|46|727|-80.810056|7|35.219587|SEASONAL CANDY-SINGLE FAC|0.3|1|I/O(H14)BF MINI BEAR FUN PACK|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00041420744259|CANDY|G1 GROCERY|-80.737839|80.737908221770127|401|1
35.297134|9811d048877613c456ac0145b70efbb6f2c2cb2f|3.98|2014-10-01 06:10:00|80.737901233649083|2|7203671215|258|35.346914866494124|0|46|225|-80.810056|35|35.219587|SUGAR-GRANULATED|0.0|1|HT GRANULATED SUGAR|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00072036712158|SUGAR/SUBSTITUTES|G1 GROCERY|-80.737839|80.737908221770127|401|2
35.297134|756e70308dc4a2a13ddf9507d01b0c06ac44381b|5.29|2014-09-15 19:47:00|80.737901233649083|2|7203698288|258|35.34691489783858|0|46|1262|-80.66939|57|35.28326|HALF N HALF WHIPPING CREAM|0.0|3|HT HEAVY CREAM|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00072036982889|MILK|DAIRY|-80.737839|80.737849194022729|46|1
35.297134|334f54db4032b8c2e619586366fbc9e029c7cb45|5.29|2014-09-16 09:37:00|80.737901233649083|2|7203698288|258|35.34691489558098|0|46|1262|-80.764523|57|35.341927|HALF N HALF WHIPPING CREAM|0.0|3|HT HEAVY CREAM|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00072036982889|MILK|DAIRY|-80.737839|80.737860013188453|220|1
35.297134|567f09d2bb629c2b2841b3eb575fd6898f0aac34|8.0|2015-01-28 07:36:00|80.737901233649083|2|85822200105|258|35.346914866494124|0|46|7209|-80.810056|1600|35.219587|BACK TO SCHOOL|6.0|18|I/OAPPLE COMPATIBLE CABLE|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00858222001059|SEASONAL MERCHANDISE|GM|-80.737839|80.737908221770127|401|1
35.297134|5572a341b6e309fa0521e127e1abd5d7dcaa1ce5|2.99|2015-01-13 09:02:00|80.737901233649083|2|3338322235|258|35.346914866494124|0|46|504|-80.810056|64|35.219587|FRESH BERRIES|0.0|4|BLUEBERRIES PINT|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00811654020036|FRESH PRODUCE|PRODUCE|-80.737839|80.737908221770127|401|1
35.297134|f2bc7ed610473fff527758c135ec410bf9d76bc1|4.24|2014-10-20 08:02:00|80.737901233649083|2||258|35.346914866494124|0|46|502|-80.810056|64|35.219587|FRESH BANANAS|0.0|4|BANANAS, YELLOW|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00204011000008|FRESH PRODUCE|PRODUCE|-80.737839|80.737908221770127|401|1
35.297134|fafc18fbf56215066006953f2c4ad933d02245ca|1.19|2014-09-16 09:38:00|80.737901233649083|2|7433686394|258|35.34691489558098|0|46|342|-80.764523|57|35.341927|FRESH MILK|0.2|3|HUNTER 2% MILK 14 OZ|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|35.349871187060224|00074336863950|MILK|DAIRY|-80.737839|80.737860013188453|220|1
35.297134|37fe25497c39ae63d379c98030ec1e68f2431e4e|6.68|2015-01-07 07:01:00|1.4094857484078087|2|7203657050|258|0.6160512048176361|0|26|687|-80.737839|61|35.297134|BLENDED|0.0|3|HT PLAIN NONFAT YOGURT|758e690e26c5db844ed611dfc012090b5178fe8d|3.4397398720937424|0.61471665291522548|00072036570505|YOGURT|DAIRY|-80.737839|1.409141121495086|258|4
34.95459|d8a5c7d2f14302ca2dc8c4c89f433664b7a46042|5.39|2015-02-12 17:48:00|1.4091206135396188|2|20596200000|182|0.6100726841846847|0|47|1821|-80.758228|410|34.95459|BH TURKEY|0.54|6|BOARS HEAD MAPLE HONEY TURKEY|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|0.61242566243833529|00205962000000|BH MEAT|DELI|-80.758228|1.4094969766762753|182|1
34.95459|4e7773284653d49a8fce2a5dbc274ae252c774bc|1.25|2014-12-27 13:27:00|80.758271881003409|2|4900005537|182|34.99821555170616|0|28|54|-80.847383|8|35.024464|DIET|0.25|23|COKE ZERO 1.25 LITER BOTTLE|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00049000055412|CARBONATED BEVERAGES|BEVERAGE|-80.758228|80.758245354037413|317|1
34.95459|dd5328f92d79065928490b0a5ed630a4f3d828e5|6.79|2014-11-25 16:53:00|1.4091206135396188|2|4900002890|182|0.6100726841846847|0|47|54|-80.758228|8|34.95459|DIET|1.8|23|FRESCA 12OZ 12PK FRIDGEPACK CN|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|0.61242566243833529|00049000031058|CARBONATED BEVERAGES|BEVERAGE|-80.758228|1.4094969766762753|182|1
34.95459|c1eb05f36d60650abd99823afa7dc30b403b108b|4.99|2015-03-07 18:12:00|80.758271881003409|2|7203695649|182|34.998215533527436|0|28|1699|-80.770346|387|35.052812|EVERYDAY (COOKIES)|1.5|14|HT CHOCO, CHOCO FROSTED COOKIE|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00072036956514|COOKIES|BAKERY|-80.758228|80.758279609797313|40|1
34.95459|1ac4cf44be6e1c449420916f16e8239546fd4a4c|7.75|2014-11-26 14:27:00|80.758271881003409|2|1258760034|182|34.998215508227183|0|28|443|-80.7007|76|35.06858|NFS-GARBAGE BAGS|0.76|1|GLAD TALL KTCH HAW ALOHA DRWST|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00012587786260|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.758228|80.758305145660316|273|1
34.95459|d90cde2f41b05f89f85b1f54a12bac4ea35139fa|3.99|2014-12-02 22:23:00|80.758271881003409|2|7203663995|182|34.99821554558163|0|28|342|-80.848528|57|35.053394|FRESH MILK|1.52|3|HARRIS TEETER 1% MILK|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00072036631275|MILK|DAIRY|-80.758228|80.758261122092662|11|1
34.95459|0e7d21fdfc47acd9f5cfe6fa4006ee7657be8f8c|2.59|2014-11-08 19:41:00|80.758271881003409|2|7203663996|182|34.998215511928066|0|28|342|-80.824767|57|35.116751|FRESH MILK|0.0|3|HARRIS TEETER 2%   MILK|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00072036639998|MILK|DAIRY|-80.758228|80.758301962859974|294|1
34.95459|88498f65b48e190c60981169da0e3496c2aaf6a5|3.99|2014-10-11 22:39:00|80.758271881003409|2|7203663995|182|34.99821555170616|0|28|342|-80.847383|57|35.024464|FRESH MILK|2.02|3|HARRIS TEETER 1% MILK|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00072036631275|MILK|DAIRY|-80.758228|80.758245354037413|317|1
34.95459|8c9c082031123226f94cd72310f6fd660c77126d|3.59|2014-11-11 18:01:00|1.4091206135396188|2|7203695890|182|0.6100726841846847|0|47|1654|-80.758228|381|34.95459|DESSERT CAKES|0.0|14|GRANDE FINALE CAKE SLICE|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|0.61242566243833529|00072036958907|CAKES|BAKERY|-80.758228|1.4094969766762753|182|1
34.95459|764277e438d5cf66a6fe20b260f15219bf6b2d99|2.5|2014-10-18 16:25:00|80.758271881003409|2|7203698670|182|34.998215533527436|0|28|99|-80.770346|32|35.052812|LIQUID TEA|0.0|1|HT DT GRN TEA W/HONEY&GINSENG|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00072036986719|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.758228|80.758279609797313|40|1
34.95459|ba41e25c3e41e1fda9c673f8084f20d0eaac7a9c|1.29|2015-01-27 17:21:00|80.758271881003409|2|7565600119|182|34.998215542116455|0|28|6407|-80.699686|1556|35.000049|BALLOONS|0.0|18|BALLOONS 20 ROUND|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00075656001190|TOYS|GM|-80.758228|80.758267336860058|249|1
34.95459|655e73c7b8806a769135f184e156771175f801c8|5.99|2014-11-03 12:55:00|80.758271881003409|2|7766113749|182|34.998215542116455|0|28|577|-80.699686|136|35.000049|OTHER MERCH FR MSC JUICE|0.0|4|LITEHOUSE HONEY CRISP CIDER|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00077661137499|OTHER MERCHANDISE|PRODUCE|-80.758228|80.758267336860058|249|1
34.95459|6d073cab2b3265fded297511c906de8b5d41beba|1.94|2014-11-20 17:37:00|1.4091206135396188|2|7203688002|182|0.6100726841846847|0|47|527|-80.758228|64|34.95459|FRESH CARROTS|0.0|4|HT WHOLE CARROTS 2LB BAG|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|0.61242566243833529|00072036880024|FRESH PRODUCE|PRODUCE|-80.758228|1.4094969766762753|182|2
34.95459|b3bed9026eff29780abd18e7f37056a8c4dd3eb4|2.58|2014-09-26 11:52:00|80.758271881003409|2|8379152001|182|34.99821554558163|0|28|1981|-80.848528|480|35.053394|CHIPS|0.0|6|DIRTY POTATO CHIP BBQ|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00083791520049|DRY GOODS|DELI|-80.758228|80.758261122092662|11|2
34.95459|0088b6818cd940fd8b2bbbc4421f409d6081168b|6.79|2014-12-04 13:33:00|1.4091206135396188|2|7800008216|182|0.6100726841846847|0|47|55|-80.758228|8|34.95459|REGULAR|1.8|23|DR PEPPER TEN   12PK CANS|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|0.61242566243833529|00078000103168|CARBONATED BEVERAGES|BEVERAGE|-80.758228|1.4094969766762753|182|1
34.95459|6c8979819060007c61e6e2a4bee405dec3b33e91|3.49|2015-01-19 15:14:00|1.4091206135396188|2|8912522000|182|0.6100726841846847|0|47|151|-80.758228|23|34.95459|DSD PASTA CORE|0.0|1|ANCIENT HRVST ORG QUIN ROTELL|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|0.61242566243833529|00089125260001|PASTA|G1 GROCERY|-80.758228|1.4094969766762753|182|1
34.95459|83098d3d54917e9877bd78457c469634a04e59b6|5.99|2015-02-20 16:37:00|1.4091206135396188|2|8981908394|182|0.6100726841846847|0|47|9945|-80.758228|885|34.95459|NFS POP OTHER WHITE|0.0|13|BERINGER CHENIN BLANC|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|0.61242566243833529|00089819083947|POPULAR (4-$7.99)|WINE|-80.758228|1.4094969766762753|182|1
34.95459|15459bf5ef5ad38f159be0479bdae57a6da3dd4e|5.09|2014-12-12 13:12:00|80.758271881003409|2|20543600000|182|34.99821555170616|0|28|1832|-80.847383|415|35.024464|BH SLICING CHEESE|0.0|6|BOARS HEAD MONTEREY JACK CHSE|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00205436000000|SLICING CHEESE|DELI|-80.758228|80.758245354037413|317|1
34.95459|409a3a0459dcd66b15c67557ee843ec03b6795e5|6.58|2014-11-18 18:05:00|80.758271881003409|2|61144334026|182|34.998215542116455|0|28|214|-80.699686|33|35.000049|BROTH|1.0|1|KITCHEN BASICS STOCK CHICKEN|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00611443340013|SOUP|G1 GROCERY|-80.758228|80.758267336860058|249|2
34.95459|24fd5a8449cbbf52cb1e0e74cd78ca813410f7c0|4.94|2015-02-03 17:52:00|1.4091206135396188|2|20541300000|182|0.6100726841846847|0|47|1832|-80.758228|415|34.95459|BH SLICING CHEESE|0.0|6|BOARS HEAD WHITE AMER CHEESE|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|0.61242566243833529|00205413000009|SLICING CHEESE|DELI|-80.758228|1.4094969766762753|182|1
34.95459|2aa03ecc25c69d1df9d57380ef67a8ba852c9d40|8.98|2015-01-05 09:14:00|80.758271881003409|2|7203636053|182|34.99821554558163|0|28|31|-80.848528|4|35.053394|NON CARBONATED WATER|3.98|1|(U)HT SPRING WATER .5 LTR 24PK|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00072036360533|BOTTLED WATER|G1 GROCERY|-80.758228|80.758261122092662|11|2
34.95459|40b6a8e2838f1e8fd65bc0c58f59cc4e50075b3e|1.99|2014-10-07 13:37:00|80.758271881003409|2|7203688083|182|34.99821555170616|0|28|526|-80.847383|64|35.024464|FRESH MUSHROOMS|0.2|4|HT WHITE MUSHROOMS, 8 OZ WHOLE|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00072036880833|FRESH PRODUCE|PRODUCE|-80.758228|80.758245354037413|317|1
34.95459|d13e6e4ad92416c8620b67adf66a6eae4f29007d|2.97|2015-01-27 17:12:00|80.758271881003409|2|7203632014|182|34.998215542116455|0|28|194|-80.699686|30|35.000049|OLIVE OIL|0.0|1|HT EXTRA VIRGIN OLIVE OIL|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00072036320148|SHORTENING/OIL|G1 GROCERY|-80.758228|80.758267336860058|249|1
34.95459|1562818395f118d3e905a224cba4d5e3150b43e3|6.99|2014-12-31 14:57:00|80.758271881003409|2|4900002890|182|34.99821554762525|0|28|54|-80.837892|8|34.937113|DIET|2.0|23|COKE ZERO 12 OZ FRIDGEPACK CN|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00049000042559|CARBONATED BEVERAGES|BEVERAGE|-80.758228|80.758256835672356|372|1
34.95459|ed1fef200b3f9dd027c5c70770016fda11caa19f|8.99|2014-09-23 16:46:00|80.758271881003409|2|8130859207|182|34.99821555170616|0|28|9947|-80.847383|886|35.024464|NFS-PREM-CHARDONNAY|0.0|13|CB-CUPCAKE CHARDONNAY|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00081308592077|PREMIUM ($8-$10.99)|WINE|-80.758228|80.758245354037413|317|1
34.95459|8e474df2651415e17261d4de4237109cbe4e6691|3.55|2014-11-12 17:12:00|80.758271881003409|2|7433610102|182|34.99821555170616|0|28|342|-80.847383|57|35.024464|FRESH MILK|0.0|3|HIGHLAND CREST WHOLE MILK|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00074336879203|MILK|DAIRY|-80.758228|80.758245354037413|317|1
34.95459|b92731abe85431633e2df6fd35807d3dc20642aa|2.17|2014-09-14 15:43:00|1.4091206135396188|2|7433610204|182|0.6100726841846847|0|47|331|-80.758228|52|34.95459|NATURAL SLICED|0.0|3|HC MILD CHEDDAR SLICES|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|0.61242566243833529|00074336102042|CHEESE|DAIRY|-80.758228|1.4094969766762753|182|1
34.95459|116ac39cc1307d3b61fc2e8c6bcd030dc1ed5d4a|2.99|2015-02-25 18:43:00|80.758271881003409|2|7433610102|182|34.99821554762525|0|28|342|-80.837892|57|34.937113|FRESH MILK|0.0|3|HIGHLAND CREST 2% REDUCE FAT|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00074336101021|MILK|DAIRY|-80.758228|80.758256835672356|372|1
34.95459|8bb56930b925a5fdd2061643bcaad56bd5475140|1.29|2014-12-24 14:30:00|80.758271881003409|2|4920005675|182|34.998215542116455|0|28|224|-80.699686|35|35.000049|SUGAR-BROWN|0.0|1|DOMINO LT BRWN SUGAR-BOX|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00049200056752|SUGAR/SUBSTITUTES|G1 GROCERY|-80.758228|80.758267336860058|249|1
34.95459|114f9c6517dbf15bdf983949d236e3b54aef14d8|7.99|2014-10-24 16:50:00|1.4091206135396188|2|1820013986|182|0.6100726841846847|0|47|458|-80.758228|82|34.95459|CRAFT BEER|0.0|16|SHOCK TOP ALE 6PK|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|0.61242566243833529|00018200139864|DOMESTIC BEER|BEER|-80.758228|1.4094969766762753|182|1
34.95459|3b07a3fdee42bde95910b873a19827cb6ad6a847|1.49|2014-11-08 09:47:00|80.758271881003409|2|2840002819|182|34.998215520491044|0|28|206|-80.85753|31|35.116638|FRONT END SNACKS|0.0|1|RUFFLES CHED SOUR CREAM|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00028400028158|SNACKS|G1 GROCERY|-80.758228|80.758294012939444|204|1
34.95459|fa8b806c02e281eb24b4731681955c9606e7a0c6|0.85|2014-12-04 16:08:00|80.758271881003409|2|7203636026|182|34.99821553880691|0|28|55|-80.816172|8|35.059823|REGULAR|0.35|23|HT CLUB SODA|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00072036360274|CARBONATED BEVERAGES|BEVERAGE|-80.758228|80.758272468861847|66|1
34.95459|f8493ff77b08b4dc7849885ad55e4c50dad5e3ed|3.49|2014-10-16 12:04:00|80.758271881003409|2|7017715419|182|34.9982155449852|0|28|233|-80.8062|37|35.037115|BLACK TEA|0.5|1|TWININGS TEA BLK VARIETY PACK|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00070177154035|TEA|G1 GROCERY|-80.758228|80.758262272172516|27|1
34.95459|9dab7ebf7d11ce57e64ea93900b61c7243535cc6|1.98|2014-12-02 17:10:00|80.758271881003409|2|20584100000|182|34.99821555170616|0|28|1804|-80.847383|400|35.024464|FFM SALAMI|0.0|6|GENOA SALAMI|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00205841000008|FFM MEAT|DELI|-80.758228|80.758245354037413|317|1
34.95459|e99215dfe90d21fcb9bce7700d46ecd19925cf48|10.5|2014-12-10 21:16:00|80.758271881003409|2|20496000000|182|34.99821555170616|0|28|755|-80.847383|87|35.024464|NFS-BALLOONS|0.0|9|*BALLOONS|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00204960000005|FLORAL|FLORAL|-80.758228|80.758245354037413|317|3
34.95459|596143f93770be01db0800cfac0a875128c328b2|10.99|2015-01-12 07:25:00|80.758271881003409|2|7017787949|182|34.998215542868358|0|28|1247|-80.760919|37|35.024332|SINGLES PODS CUPS TEA|2.0|1|TWININGS TEA KCUP CHAI LATTE|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00070177879495|TEA|G1 GROCERY|-80.758228|80.758266074609352|343|1
34.95459|8abc3107bf1d72ef4015389d51396438e17cb09e|12.99|2015-02-06 18:06:00|80.758271881003409|2|1820015981|182|34.998215542116455|0|28|458|-80.699686|82|35.000049|CRAFT BEER|0.0|16|SHOCK TOP 12PK BOTTLES|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00018200159817|DOMESTIC BEER|BEER|-80.758228|80.758267336860058|249|1
34.95459|8dcf065f14460d4cc0abcad9a6f1608be5370f2d|2.69|2014-12-22 10:28:00|80.758271881003409|2|7203618197|182|34.99821555170616|0|28|6674|-80.847383|1564|35.024464|MAILING SUPPLIES TAPE|0.0|18|(FE)HT 2X1000 CLR MAILING TP|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00072036181978|SCHOOL & OFFICE SUPPLY|GM|-80.758228|80.758245354037413|317|1
34.95459|b63559890ea42571edf17b6d6eed37a1a9a9c0da|2.29|2015-01-08 21:38:00|80.758271881003409|2|3680031151|182|34.99821554868852|0|28|4502|-80.992182|1210|35.103409|LAXATIVE-STIMULANT|0.0|17|TC LAXATIVE ENEMA TWIN PK|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00036800311510|STOMACH REMEDIES|HBC|-80.758228|80.758254330947935|88|1
34.95459|53cea3b07ff1fd6b2b2096cd6fad1b3fd758c678|12.0|2015-02-10 16:45:00|80.758271881003409|2|84115200732|182|34.998215542116455|0|28|1165|-80.699686|87|35.000049|NFS-FRESH CONSUMER BUNCH|0.0|9|BUNCH- 3/$12 DAISY BUNCHES|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00841152007321|FLORAL|FLORAL|-80.758228|80.758267336860058|249|3
34.95459|39834fd97569359b9484c90b0aa472d3a9b083a8|1.39|2014-12-17 13:46:00|80.758271881003409|2|8265750067|182|34.99821554558163|0|28|31|-80.848528|4|35.053394|NON CARBONATED WATER|0.39|1|DEER PARK WATER 1LT|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00082657500676|BOTTLED WATER|G1 GROCERY|-80.758228|80.758261122092662|11|1
34.95459|1280662da87501826c3b123677ced5504f66773c|5.38|2015-01-05 09:15:00|80.758271881003409|2|3663202720|182|34.99821554558163|0|28|687|-80.848528|61|35.053394|BLENDED|0.69|3|DANNON RASP GOJI/ BLUE ACAI|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00036632021878|YOGURT|DAIRY|-80.758228|80.758261122092662|11|2
34.95459|768f99a4a6250907b9d0b0378e84f20512c555c6|7.65|2014-12-15 17:39:00|80.758271881003409|2|76211120604|182|34.99821555170616|0|28|35|-80.847383|10|35.024464|PREMIUM WHOLE BEAN|0.0|1|STARBUCKS SUMATRA WHL BEAN|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00762111622907|COFFEE|G1 GROCERY|-80.758228|80.758245354037413|317|1
34.95459|f9664c3cafdcacc01d206a87e70362372eb3c807|7.99|2014-10-11 22:46:00|80.758271881003409|2|89627000010|182|34.99821555170616|0|28|458|-80.847383|82|35.024464|CRAFT BEER|0.0|16|BIG BOSS HELL'S BELLE 6PK|75e7baf78fac4320cb7caa6574ab3500f81461ce|3.0144204310898743|34.992988447249964|00896270000105|DOMESTIC BEER|BEER|-80.758228|80.758245354037413|317|1
35.141204|abcb463d5f5f50183e89bb9f902f0d3e2bc8063c|7.99|2015-03-01 15:46:00|80.739023103730261|3|3077109653|171|35.170833847164609|0|16|499|-80.80146|110|35.17739|MEATBALLS|1.0|19|ALFRESCO MEATBALL ITALIAN|762b1b33f0fae7ebe2081ff643352dcc0922c57d|2.0473508945345538|35.169056414731678|00030771096544|FROZEN CASE MEAT|CASE READY MEATS|-80.739|80.739003394444566|208|1
35.141204|3517c91fd25c48ec8b80ae63c6017590351c5645|3.49|2015-02-14 15:26:00|80.739023103730261|3|7373100419|171|35.170833842304802|0|16|495|-80.732725|108|35.082768|NON REFRIGERATED|0.0|19|MISSION FLOUR TORTILLAS 8 CT|762b1b33f0fae7ebe2081ff643352dcc0922c57d|2.0473508945345538|35.169056414731678|00073731004197|TORTILLAS|CASE READY MEATS|-80.739|80.739021032245986|147|1
35.141204|d74c18682ceccf5f9e1606d86df0cec72e79d89e|9.99|2015-01-13 17:14:00|1.4091206135396188|3|7570615102|171|0.6133297129150015|0|47|254|-80.739|892|35.141204|PREMIUM PIZZA|0.0|5|PALERMOS  SS SPICY CLUCKER|762b1b33f0fae7ebe2081ff643352dcc0922c57d|2.0473508945345538|0.61242566243833529|00075706151059|FROZEN PIZZA|FROZEN|-80.739|1.4091613847677018|171|1
35.141204|83c7deabad9d44bc693aaa42640cb45db40fd1b8|2.01|2015-02-04 17:37:00|1.4091206135396188|3|7203637030|171|0.6133297129150015|0|47|212|-80.739|33|35.141204|CONDENSED SOUP|0.0|1|HT SP CHICKEN NOODLE|762b1b33f0fae7ebe2081ff643352dcc0922c57d|2.0473508945345538|0.61242566243833529|00072036370334|SOUP|G1 GROCERY|-80.739|1.4091613847677018|171|3
35.141204|c6fb8c27685d60641ebb82193ad32f406685acc3|7.99|2014-09-16 17:05:00|1.4091206135396188|3|1820017993|171|0.6133297129150015|0|47|458|-80.739|82|35.141204|CRAFT BEER|0.0|16|SHOCK TOP SEASONAL 6PK|762b1b33f0fae7ebe2081ff643352dcc0922c57d|2.0473508945345538|0.61242566243833529|00018200179938|DOMESTIC BEER|BEER|-80.739|1.4091613847677018|171|1
35.141204|dd53f51d182651c851edf24648a3b9382eaadd46|2.29|2014-09-24 17:28:00|1.4091206135396188|3|31254662920|171|0.6133297129150015|0|47|4207|-80.739|1200|35.141204|COUGH DROP-ADULT|0.0|17|HALLS DEF VIT. C WMLN-63158|762b1b33f0fae7ebe2081ff643352dcc0922c57d|2.0473508945345538|0.61242566243833529|00312546631588|COUGH/COLD/SINUS|HBC|-80.739|1.4091613847677018|171|1
35.141204|92e8d33499c92b96e1b3b787d84bc4f756a237d8|26.3|2015-03-08 11:26:00|80.739023103730261|3|20496000000|171|35.170833847164609|0|16|755|-80.80146|87|35.17739|NFS-BALLOONS|0.0|9|*BALLOONS|762b1b33f0fae7ebe2081ff643352dcc0922c57d|2.0473508945345538|35.169056414731678|00204960000005|FLORAL|FLORAL|-80.739|80.739003394444566|208|1
35.141204|6df5397fca7d878bcde3a87043dbb6de987f1bc3|0.77|2014-10-06 17:21:00|1.4091206135396188|3||171|0.6133297129150015|0|47|522|-80.739|64|35.141204|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|762b1b33f0fae7ebe2081ff643352dcc0922c57d|2.0473508945345538|0.61242566243833529|00204664000004|FRESH PRODUCE|PRODUCE|-80.739|1.4091613847677018|171|1
35.141204|55b7672e707b0da280ce1dbbc5238506e246877f|19.99|2014-10-02 16:58:00|1.4091206135396188|3|8210073846|171|0.6133297129150015|0|47|9924|-80.739|882|35.141204|NFS-PREMIUM BOX|0.0|13|BLACK BOX MALBEC 3L|762b1b33f0fae7ebe2081ff643352dcc0922c57d|2.0473508945345538|0.61242566243833529|00082100738465|PREMIUM BOX|WINE|-80.739|1.4091613847677018|171|1
35.141204|d74ebc477fb08ca6431ec4fe81a940290a61a3fb|29.98|2015-01-16 12:35:00|1.4091206135396188|3|7199031600|171|0.6133297129150015|0|47|455|-80.739|82|35.141204|DOMESTIC PREMIUM 12PK&>|0.0|16|COORS LIGHT 24PK 12OZ CAN|762b1b33f0fae7ebe2081ff643352dcc0922c57d|2.0473508945345538|0.61242566243833529|00071990316006|DOMESTIC BEER|BEER|-80.739|1.4091613847677018|171|2
35.141204|242a3dd70d87b133dcdab85b77456e8419bfa17b|29.98|2015-01-06 17:00:00|1.4091206135396188|3|7199031600|171|0.6133297129150015|0|47|455|-80.739|82|35.141204|DOMESTIC PREMIUM 12PK&>|0.0|16|COORS LIGHT 24PK 12OZ CAN|762b1b33f0fae7ebe2081ff643352dcc0922c57d|2.0473508945345538|0.61242566243833529|00071990316006|DOMESTIC BEER|BEER|-80.739|1.4091613847677018|171|2
35.141204|e42c7a1b25efb4c19a9f621f272b3140f262106c|5.0|2015-01-10 11:31:00|80.739023103730261|3|4138753020|171|35.170833847276391|0|16|120|-80.709466|15|35.124987|COATINGS & BREADERS|1.42|1|4C PANKO BREAD CRUMBS|762b1b33f0fae7ebe2081ff643352dcc0922c57d|2.0473508945345538|35.169056414731678|00041387530209|FLOUR|G1 GROCERY|-80.739|80.739001269626044|157|2
35.141204|de81c572451536b3b1c54902211ceeed3765cd1a|3.49|2014-09-15 16:52:00|1.4091206135396188|3|4610000012|171|0.6133297129150015|0|47|318|-80.739|52|35.141204|SHREDDED/GRATED CHEESE|0.0|3|SARGENTO OTB 4 CHSE MEX FINE C|762b1b33f0fae7ebe2081ff643352dcc0922c57d|2.0473508945345538|0.61242566243833529|00046100000922|CHEESE|DAIRY|-80.739|1.4091613847677018|171|1
35.141204|6156c89ddf1a085c706e4a29e343629c519c6b0a|3.89|2014-09-18 13:07:00|80.739023103730261|3|4400002827|171|35.170833834599989|0|16|1251|-80.771677|12|35.066546|WHOLESOME COOKIES|0.89|1|BELVITA BREAKFAST APPLE CINN|762b1b33f0fae7ebe2081ff643352dcc0922c57d|2.0473508945345538|35.169056414731678|00044000028251|COOKIES|G1 GROCERY|-80.739|80.739033547083153|45|1
35.141204|988741869fa156e8b46dddaf0fe6bc991e45ffee|12.99|2015-01-29 17:10:00|1.4091206135396188|3|5400041821|171|0.6133297129150015|0|47|426|-80.739|72|35.141204|NFS-PAPER TOWELS|0.0|1|SCOTT NAT TOWEL TUBE FREE 12MR|762b1b33f0fae7ebe2081ff643352dcc0922c57d|2.0473508945345538|0.61242566243833529|00054000418211|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.739|1.4091613847677018|171|1
35.141204|6dced3abcea4682e77337a51b3f05c7a3c64cda0|3.79|2014-12-16 17:29:00|1.4091206135396188|3|7203688014|171|0.6133297129150015|0|47|581|-80.739|136|35.141204|FRESH SALSA|0.0|4|HT FRESH MEDIUM SALSA|762b1b33f0fae7ebe2081ff643352dcc0922c57d|2.0473508945345538|0.61242566243833529|00072036880222|OTHER MERCHANDISE|PRODUCE|-80.739|1.4091613847677018|171|1
35.141204|b8e79c04e490a92dfce4d1200b51607488e36116|3.69|2015-01-05 12:01:00|80.739023103730261|3|4400001570|171|35.170833834599989|0|16|1256|-80.771677|13|35.066546|WHOLESOME CRACKERS|0.69|1|RITZ TOASTED CHIPS CHEDDAR|762b1b33f0fae7ebe2081ff643352dcc0922c57d|2.0473508945345538|35.169056414731678|00044000015701|CRACKERS|G1 GROCERY|-80.739|80.739033547083153|45|1
35.141204|595406202c1e6fc489ba2596f858588aab9f5985|3.49|2014-11-15 14:42:00|1.4091206135396188|3|4400001473|171|0.6133297129150015|0|47|1248|-80.739|12|35.141204|SANDWICH COOKIES|0.49|1|WHITE FUDGE OREO|762b1b33f0fae7ebe2081ff643352dcc0922c57d|2.0473508945345538|0.61242566243833529|00044000014735|COOKIES|G1 GROCERY|-80.739|1.4091613847677018|171|1
35.141204|90c9fe332e752f7de077233848be1adba81f87d7|4.99|2014-10-14 07:18:00|80.739023103730261|3|7336070341|171|35.170833842304802|0|16|30|-80.732725|4|35.082768|CARBONATED WATER|0.0|1|LACROIX WTR CRAN RSP 12PK|762b1b33f0fae7ebe2081ff643352dcc0922c57d|2.0473508945345538|35.169056414731678|00073360323416|BOTTLED WATER|G1 GROCERY|-80.739|80.739021032245986|147|1
35.141204|1f24b0c87dd01c02704efe429ccd970a4fa50cee|3.39|2014-09-19 16:23:00|80.739023103730261|3|4920004550|171|35.1708338406441|0|16|225|-80.78468|35|35.096737|SUGAR-GRANULATED|0.0|1|DOMINO GRANULATED SUGAR 4 LB|762b1b33f0fae7ebe2081ff643352dcc0922c57d|2.0473508945345538|35.169056414731678|00049200045503|SUGAR/SUBSTITUTES|G1 GROCERY|-80.739|80.739024281293382|30|1
35.141204|08a7cba2d45c86678bec67128ba62915b1c6e771|4.49|2014-09-13 16:03:00|80.739023103730261|3|4812127707|171|35.170833847276391|0|16|1036|-80.709466|164|35.124987|BREAKFAST BAGELS|0.0|7|THOMAS PUMPKIN BAGELS 6CT PP|762b1b33f0fae7ebe2081ff643352dcc0922c57d|2.0473508945345538|35.169056414731678|00048121226220|BREAKFAST|COMMERCIAL BAKERY|-80.739|80.739001269626044|157|1
35.006282|1681993a991718703018380ab0e8fa7a701c6174|12.59|2014-11-10 15:02:00|1.4091206135396188|4|20598600000|60|0.6109748797816256|0|47|1800|-80.562829|400|35.006282|FFM BEEF|2.1|6|HT ROAST  BEEF|7a9fe7b0685b663a067825eca6e51e9f5eeda85f|0.4474017081721333|0.61242566243833529|00205986000000|FFM MEAT|DELI|-80.562829|1.4060866207711706|60|1
35.006282|a020841f036b23b4321b546b4d4704088d2f587d|7.98|2015-01-07 14:57:00|80.562862110758871|4|1630016564|60|35.012756925386626|0|21|335|-80.64817|56|35.04711|ORANGE JUICE-REGRIGERATED|0.0|3|FL NAT W/PULP ORANGE JUICE|7a9fe7b0685b663a067825eca6e51e9f5eeda85f|0.4474017081721333|35.054042368968126|00016300165653|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.562829|80.562829308840179|129|2
35.006282|e7a057b5199bc2e994c8592f301587f5be710843|5.99|2014-11-21 11:33:00|80.562862110758871|4|5450010174|60|35.012756925386626|0|21|485|-80.64817|101|35.04711|PREMIUM WIENERS|0.0|19|BALL PARK LEAN ANGUS FRANK|7a9fe7b0685b663a067825eca6e51e9f5eeda85f|0.4474017081721333|35.054042368968126|00054500193397|WIENERS|CASE READY MEATS|-80.562829|80.562829308840179|129|1
35.006282|2de7406f8f1c0070458e02a4cedb25f1223a6c2d|2.69|2015-02-17 18:36:00|80.562862110758871|4|7225001739|60|35.012756925386626|0|21|1025|-80.64817|162|35.04711|WHITE|0.5|7|NATOWN WHITEWHEAT RTOP BRD|7a9fe7b0685b663a067825eca6e51e9f5eeda85f|0.4474017081721333|35.054042368968126|00072250017398|SLICED BREAD|COMMERCIAL BAKERY|-80.562829|80.562829308840179|129|1
35.006282|d09d0a5daddbbafd0c1565224879b44f248ba66a|2.69|2015-02-03 09:58:00|80.562862110758871|4|7225001739|60|35.012756925386626|0|21|1025|-80.64817|162|35.04711|WHITE|0.0|7|NATOWN WHITEWHEAT RTOP BRD|7a9fe7b0685b663a067825eca6e51e9f5eeda85f|0.4474017081721333|35.054042368968126|00072250017398|SLICED BREAD|COMMERCIAL BAKERY|-80.562829|80.562829308840179|129|1
35.006282|6d888718d13702a51e80d03ab40d9fdb0fb49e89|2.69|2015-01-14 17:57:00|80.562862110758871|4|7225001739|60|35.012756925386626|0|21|1025|-80.64817|162|35.04711|WHITE|0.0|7|NATOWN WHITEWHEAT RTOP BRD|7a9fe7b0685b663a067825eca6e51e9f5eeda85f|0.4474017081721333|35.054042368968126|00072250017398|SLICED BREAD|COMMERCIAL BAKERY|-80.562829|80.562829308840179|129|1
35.006282|d27ac2c6de5e2b71c5de940e0a7ed7c7d3bddec3|2.69|2014-12-11 16:08:00|1.4091206135396188|4|7225001739|60|0.6109748797816256|0|47|1025|-80.562829|162|35.006282|WHITE|0.5|7|NATOWN WHITEWHEAT RTOP BRD|7a9fe7b0685b663a067825eca6e51e9f5eeda85f|0.4474017081721333|0.61242566243833529|00072250017398|SLICED BREAD|COMMERCIAL BAKERY|-80.562829|1.4060866207711706|60|1
35.006282|3d9e07af5b1ca5cd2173e1701d43c88835ac3ec8|2.69|2014-12-02 11:53:00|80.562862110758871|4|7225001739|60|35.012756925386626|0|21|1025|-80.64817|162|35.04711|WHITE|0.0|7|NATOWN WHITEWHEAT RTOP BRD|7a9fe7b0685b663a067825eca6e51e9f5eeda85f|0.4474017081721333|35.054042368968126|00072250017398|SLICED BREAD|COMMERCIAL BAKERY|-80.562829|80.562829308840179|129|1
35.006282|3418d818094fa4e54207ef46814e7f6ffff35f2f|2.69|2014-10-15 14:39:00|1.4091206135396188|4|7225001739|60|0.6109748797816256|0|47|1025|-80.562829|162|35.006282|WHITE|0.5|7|NATOWN WHITEWHEAT RTOP BRD|7a9fe7b0685b663a067825eca6e51e9f5eeda85f|0.4474017081721333|0.61242566243833529|00072250017398|SLICED BREAD|COMMERCIAL BAKERY|-80.562829|1.4060866207711706|60|1
35.006282|2b3415b6529e96fdb2209feddd952f80b23cfdef|2.69|2015-03-02 10:51:00|1.4091206135396188|4|7225001739|60|0.6109748797816256|0|47|1025|-80.562829|162|35.006282|WHITE|0.5|7|NATOWN WHITEWHEAT RTOP BRD|7a9fe7b0685b663a067825eca6e51e9f5eeda85f|0.4474017081721333|0.61242566243833529|00072250017398|SLICED BREAD|COMMERCIAL BAKERY|-80.562829|1.4060866207711706|60|1
35.006282|56f36554d3f27f636627daa19fe7eb478b99773b|2.69|2015-03-09 16:35:00|80.562862110758871|4|7225001739|60|35.012756925386626|0|21|1025|-80.64817|162|35.04711|WHITE|0.0|7|NATOWN WHITEWHEAT RTOP BRD|7a9fe7b0685b663a067825eca6e51e9f5eeda85f|0.4474017081721333|35.054042368968126|00072250017398|SLICED BREAD|COMMERCIAL BAKERY|-80.562829|80.562829308840179|129|1
35.006282|b8b2ded81375957b7c8a0419e069aaed923c39a3|2.69|2014-12-22 19:15:00|80.562862110758871|4|7225001739|60|35.012756925386626|0|21|1025|-80.64817|162|35.04711|WHITE|1.35|7|NATOWN WHITEWHEAT RTOP BRD|7a9fe7b0685b663a067825eca6e51e9f5eeda85f|0.4474017081721333|35.054042368968126|00072250017398|SLICED BREAD|COMMERCIAL BAKERY|-80.562829|80.562829308840179|129|1
35.006282|e507bc6638873a93d96d6baa369900f6d6ad63d8|14.99|2014-10-03 19:16:00|80.562862110758871|4|1820053218|60|35.012756925379158|0|21|455|-80.78468|82|35.096737|DOMESTIC PREMIUM 12PK&>|0.0|16|BUD LIGHT 18PK 12OZ CAN|7a9fe7b0685b663a067825eca6e51e9f5eeda85f|0.4474017081721333|35.054042368968126|00018200532184|DOMESTIC BEER|BEER|-80.562829|80.562829489316272|30|1
35.006282|5d3a43bbc7fd55b9f68686e942a3d41af0f85b65|11.43|2014-10-27 14:34:00|80.562862110758871|4|20596200000|60|35.012756925386626|0|21|1821|-80.64817|410|35.04711|BH TURKEY|2.08|6|BOARS HEAD MAPLE HONEY TURKEY|7a9fe7b0685b663a067825eca6e51e9f5eeda85f|0.4474017081721333|35.054042368968126|00205962000000|BH MEAT|DELI|-80.562829|80.562829308840179|129|1
35.006282|84fb0b80fe113f0f6eec5cd232011f05a73a1b33|2.79|2015-01-12 13:29:00|80.562862110758871|4|7203698374|60|35.01275692538907|0|21|423|-80.732725|72|35.082768|NFS-DISPOSE PLATES/BOWLS|0.0|1|YH ULTRA DESIGNER PLATES|7a9fe7b0685b663a067825eca6e51e9f5eeda85f|0.4474017081721333|35.054042368968126|00072036983725|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.562829|80.562829219313898|147|1
35.006282|257130e72670dc1f27d5a155c9cb919f8d90445d|15.99|2015-02-14 15:55:00|80.562862110758871|4|20310500000|60|35.012756925386626|0|21|1153|-80.64817|87|35.04711|NFS-FRESH CUT ARRANGE|0.0|9|*BUDVASE|7a9fe7b0685b663a067825eca6e51e9f5eeda85f|0.4474017081721333|35.054042368968126|00203105000009|FLORAL|FLORAL|-80.562829|80.562829308840179|129|1
35.006282|ee08c7b490fbc9388032a3464a4659d20bff8b98|2.25|2015-01-10 12:28:00|80.562862110758871|4|7203663215|60|35.01275692538907|0|21|330|-80.732725|55|35.082768|EGGS|0.0|3|HT GRADE A    JUMBO WHITE EGGS|7a9fe7b0685b663a067825eca6e51e9f5eeda85f|0.4474017081721333|35.054042368968126|00072036632159|EGGS FRESH|DAIRY|-80.562829|80.562829219313898|147|1
35.585842|df9435e28be166925d3aa8a9d18b31fca6a8c886|4.99|2015-01-06 13:31:00|1.4102725052409182|3|1200001425|99|0.6210901099944839|1|1|54|-80.875654|8|35.585842|DIET|1.0|23|DT PEPSI 8 PK 12 OZ PET BOTTLE|80ff9063f6c3081131625fb62e311ca30814a57a|2.0992101274652777|0.61833652052202714|00012000014307|CARBONATED BEVERAGES|BEVERAGE|-80.875654|1.411546447003722|99|1
35.585842|c6ad7f5b42e108a3a9e01696a15ecfb92f5cd026|5.49|2015-01-27 11:43:00|1.4102725052409182|3|1200001425|99|0.6210901099944839|1|1|54|-80.875654|8|35.585842|DIET|0.5|23|DT PEPSI 8 PK 12 OZ PET BOTTLE|80ff9063f6c3081131625fb62e311ca30814a57a|2.0992101274652777|0.61833652052202714|00012000014307|CARBONATED BEVERAGES|BEVERAGE|-80.875654|1.411546447003722|99|1
35.585842|978e030eead039ab9a330764336e3c767b169819|4.99|2014-10-21 14:43:00|1.4102725052409182|3|1200001425|99|0.6210901099944839|1|1|54|-80.875654|8|35.585842|DIET|1.0|23|DT PEPSI 8 PK 12 OZ PET BOTTLE|80ff9063f6c3081131625fb62e311ca30814a57a|2.0992101274652777|0.61833652052202714|00012000014307|CARBONATED BEVERAGES|BEVERAGE|-80.875654|1.411546447003722|99|1
35.585842|a04df4b524717b33d9d57de4c93567eac9b52ed3|4.99|2014-11-11 14:45:00|1.4102725052409182|3|1200001425|99|0.6210901099944839|1|1|54|-80.875654|8|35.585842|DIET|1.0|23|DT PEPSI 8 PK 12 OZ PET BOTTLE|80ff9063f6c3081131625fb62e311ca30814a57a|2.0992101274652777|0.61833652052202714|00012000014307|CARBONATED BEVERAGES|BEVERAGE|-80.875654|1.411546447003722|99|1
35.585842|f014d03ad7866491093ce4e038fa3940de900a2e|4.69|2014-10-27 16:36:00|1.4102725052409182|3|7203695754|99|0.6210901099944839|0|1|1603|-80.875654|371|35.585842|PRIVATE LABEL BREAD|0.0|14|BAND OF BAKERS ROASTED GARLIC|80ff9063f6c3081131625fb62e311ca30814a57a|2.0992101274652777|0.61833652052202714|00072036957542|BREAD|BAKERY|-80.875654|1.411546447003722|99|1
35.585842|21e7a75629188dcc189dbf57b3dda0e109bac54e|3.69|2015-02-04 10:43:00|1.4102725052409182|3|4300095051|99|0.6210901099944839|1|1|209|-80.875654|20|35.585842|POWDERED SOFT DRINKS|0.0|1|CRYSTAL LIGHT RASPBERRY ICE 12|80ff9063f6c3081131625fb62e311ca30814a57a|2.0992101274652777|0.61833652052202714|00043000950685|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.875654|1.411546447003722|99|1
35.585842|84d08e804716f70f3fd7b650cecd5f0a81f5e72e|3.58|2015-02-11 14:02:00|1.4102725052409182|3|3940001614|99|0.6210901099944839|1|1|243|-80.875654|39|35.585842|BAKED BEANS|0.0|1|BUSH BKD BEAN VEGETARIAN 28|80ff9063f6c3081131625fb62e311ca30814a57a|2.0992101274652777|0.61833652052202714|00039400016359|VEGETABLES-CAN/JAR|G1 GROCERY|-80.875654|1.411546447003722|99|2
35.585842|99f6af58255f77dc7399ac88cb47fc4135c0ffd4|5.58|2014-11-25 14:56:00|1.4102725052409182|3|1800000501|99|0.6210901099944839|1|1|328|-80.875654|54|35.585842|SWEET ROLLS-REFRIGERATED|1.58|3|PILLSBURY CINNAMON ROLLS|80ff9063f6c3081131625fb62e311ca30814a57a|2.0992101274652777|0.61833652052202714|00018000005017|DOUGH PRODUCTS|DAIRY|-80.875654|1.411546447003722|99|2
35.585842|b74d0deb40900ff103e05a3a4a6d4c1622e5e648|8.7|2014-09-12 19:40:00|1.4102725052409182|3|4400002747|99|0.6210901099944839|0|1|91|-80.875654|13|35.585842|SPRAYED BUTTER CRACKERS|2.17|1|RITZ CRACKERS|80ff9063f6c3081131625fb62e311ca30814a57a|2.0992101274652777|0.61833652052202714|00044000031114|CRACKERS|G1 GROCERY|-80.875654|1.411546447003722|99|2
35.585842|955fae2cb9e04b26de0e004099709bef5200ed4b|2.34|2014-09-29 13:55:00|1.4102725052409182|3|20039000000|99|0.6210901099944839|1|1|1801|-80.875654|400|35.585842|FFM TURKEY|0.0|6|HONEY SMOKED TURKEY BREAST|80ff9063f6c3081131625fb62e311ca30814a57a|2.0992101274652777|0.61833652052202714|00200397000007|FFM MEAT|DELI|-80.875654|1.411546447003722|99|1
35.478031|d5827b2680f3ce625cecf33136f6bfe8ce0250b8|2.59|2014-11-05 17:40:00|80.8939826282094|2|7203663996|179|35.49452270106449|0|2|342|-80.8955|57|35.4437|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|35.490689277687849|00072036631299|MILK|DAIRY|-80.893784|80.893791368780597|272|1
35.478031|0919945c430ace11478564d4acf5b6409876523f|2.59|2014-11-16 10:43:00|80.8939826282094|2|7203663996|179|35.494522699524069|0|2|342|-80.86175|57|35.40953|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|35.490689277687849|00072036631299|MILK|DAIRY|-80.893784|80.893795442534781|209|1
35.478031|6f665f978cac49a1d0187ea6cd410cc1c4763910|2.0|2015-02-01 13:43:00|1.4102725052409182|2|7203605067|179|0.6192084530746164|0|1|60|-80.893784|9|35.478031|HOT CEREAL|0.0|1|HT OATS 18 OLD FASHIONED|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|0.61833652052202714|00072036050670|CEREAL|G1 GROCERY|-80.893784|1.4118628751971085|179|1
35.478031|691041783dac799167d7ae3010b39775a9990ee5|1.97|2014-12-18 18:31:00|1.4102725052409182|2|7203613031|179|0.6192084530746164|0|1|716|-80.893784|15|35.478031|SELF-RISING|0.0|1|HARRIS TEETER S/RISING FLOUR|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|0.61833652052202714|00072036130310|FLOUR|G1 GROCERY|-80.893784|1.4118628751971085|179|1
35.478031|531a2d094a651d5b8ae667f9b984a3a3add01b3c|1.98|2014-11-25 20:34:00|1.4102725052409182|2|7203698291|179|0.6192084530746164|0|1|245|-80.893784|39|35.478031|VEGETABLES-CORE|0.44|1|HT CORN WK GOLDEN NS|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|0.61833652052202714|00072036411822|VEGETABLES-CAN/JAR|G1 GROCERY|-80.893784|1.4118628751971085|179|2
35.478031|1e9df1b82e5958406f6cc7092c17d88691b59b86|1.39|2014-10-31 15:34:00|1.4102725052409182|2|7152401767|179|0.6192084530746164|0|1|1214|-80.893784|272|35.478031|AUTHENTIC HISPANIC|0.0|1|LA PREF BLACK BEANS W/S|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|0.61833652052202714|00071524017676|HISPANIC PREP. FOODS|G1 GROCERY|-80.893784|1.4118628751971085|179|1
35.478031|3eddd03bb490caf5433f2e2934114183935f42af|5.49|2014-12-04 19:42:00|1.4102725052409182|2|7352585596|179|0.6192084530746164|0|1|7431|-80.893784|1600|35.478031|CHRISTMAS GIFT BOXES|1.99|18|TREAT BOX CMAS 6CT|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|0.61833652052202714|00073525855967|SEASONAL MERCHANDISE|GM|-80.893784|1.4118628751971085|179|1
35.478031|3278f7a059dea5dfc485322d50dfc196ff766bdd|20.37|2015-01-24 10:52:00|1.4102725052409182|2|7800001180|179|0.6192084530746164|0|1|55|-80.893784|8|35.478031|REGULAR|3.4|23|CHEERWINE 12PK CANS|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|0.61833652052202714|00070925000102|CARBONATED BEVERAGES|BEVERAGE|-80.893784|1.4118628751971085|179|3
35.478031|f9a79a174357583cdee3314c4ebe762d26a7608f|1.69|2014-09-28 10:05:00|1.4102725052409182|2|7203688003|179|0.6192084530746164|0|1|527|-80.893784|64|35.478031|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|0.61833652052202714|00072036880031|FRESH PRODUCE|PRODUCE|-80.893784|1.4118628751971085|179|1
35.478031|28194f9964333ee88a052a80ad08d66193d636bd|2.79|2014-09-19 16:00:00|1.4102725052409182|2|7203688211|179|0.6192084530746164|0|1|555|-80.893784|64|35.478031|PACKAGED SALADS|0.0|4|HT PREMIUM ROMAINE|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|0.61833652052202714|00072036882110|FRESH PRODUCE|PRODUCE|-80.893784|1.4118628751971085|179|1
35.478031|891611bf1cebfa9f439ebf2a3d69e912a33b4bc0|1.69|2014-09-13 15:31:00|1.4102725052409182|2|7203688003|179|0.6192084530746164|0|1|527|-80.893784|64|35.478031|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|0.61833652052202714|00072036880031|FRESH PRODUCE|PRODUCE|-80.893784|1.4118628751971085|179|1
35.478031|2e9e406196a81d0ad666ebf3c25447defe86a6ea|1.69|2014-09-21 10:19:00|1.4102725052409182|2|7203688003|179|0.6192084530746164|0|1|527|-80.893784|64|35.478031|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|0.61833652052202714|00072036880031|FRESH PRODUCE|PRODUCE|-80.893784|1.4118628751971085|179|1
35.478031|baaa30411b67889b7481f76c10555e1fda854d35|1.69|2014-11-03 17:28:00|1.4102725052409182|2|7203688003|179|0.6192084530746164|0|1|527|-80.893784|64|35.478031|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|0.61833652052202714|00072036880031|FRESH PRODUCE|PRODUCE|-80.893784|1.4118628751971085|179|1
35.478031|55acc2976790a2c53c78a73d067ed73c61ac1956|3.79|2014-12-22 15:20:00|80.8939826282094|2|2100062503|179|35.49452270106449|0|2|318|-80.8955|52|35.4437|SHREDDED/GRATED CHEESE|1.29|3|KRAFT SHREDDED FIVE CHEESE|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|35.490689277687849|00021000607082|CHEESE|DAIRY|-80.893784|80.893791368780597|272|1
35.478031|7cea27ea8dfea0032ac164ce4e061782484d96a9|2.49|2014-09-22 19:07:00|1.4102725052409182|2|4150108320|179|0.6192084530746164|0|1|77|-80.893784|272|35.478031|HISP SAUCES/SEASONINGS|0.82|1|ORTEGA SKILLET SC FAJITA|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|0.61833652052202714|00041501083215|HISPANIC PREP. FOODS|G1 GROCERY|-80.893784|1.4118628751971085|179|1
35.478031|9f7f07aa05fef51cf0d047126b77c2b9dffd9cf4|4.29|2015-01-15 17:24:00|1.4102725052409182|2|2840015636|179|0.6192084530746164|0|1|204|-80.893784|31|35.478031|TORTILLA CHIPS|0.0|1|DORTIOS NACHO CHEESE|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|0.61833652052202714|00028400156363|SNACKS|G1 GROCERY|-80.893784|1.4118628751971085|179|1
35.478031|ce69029f1f9ecea8d99c76ce7aac02e4f361240c|9.47|2014-09-30 17:25:00|1.4102725052409182|2|20744800000|179|0.6192084530746164|0|1|1945|-80.893784|465|35.478031|SUPERFLAG CHEF CASE|0.0|6|COCONUT CHICKEN|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|0.61833652052202714|00207448000009|COLD PREPARED FOODS|DELI|-80.893784|1.4118628751971085|179|1
35.478031|b6ee7768809aeef3c070df14e808a9d5315ee90b|3.98|2014-12-20 12:49:00|80.8939826282094|2|64420900438|179|35.494522701825836|0|2|24|-80.861571|3|35.444615|FROSTING-READY-TO-SPREAD|1.0|1|DH CHOCOLATE FROSTING|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|35.490689277687849|00644209004461|BAKING SUPPLIES|G1 GROCERY|-80.893784|80.893788052598069|340|2
35.478031|ed009a54ca93e4b08ba6d30fa2a7674eef68a4f6|11.15|2014-12-11 18:18:00|1.4102725052409182|2|2550000367|179|0.6192084530746164|0|1|66|-80.893784|10|35.478031|GROUND CAN|0.0|1|FOLGERS CLASSIC ROAS CONTAINER|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|0.61833652052202714|00025500003672|COFFEE|G1 GROCERY|-80.893784|1.4118628751971085|179|1
35.478031|aaca4d52da3b896154d68d7b9015a318a03ec2b2|5.99|2014-10-04 16:56:00|1.4102725052409182|2|3545777001|179|0.6192084530746164|0|1|1611|-80.893784|371|35.478031|PITA'S AND FLAT BREADS|3.0|14|MAMA MARYS THIN CRUST 12 IN|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|0.61833652052202714|00035457770084|BREAD|BAKERY|-80.893784|1.4118628751971085|179|1
35.478031|40e46ec54c24521be1988da3b1e26449881d6ee7|9.99|2015-02-13 15:16:00|1.4102725052409182|2|7203678030|179|0.6192084530746164|0|1|458|-80.893784|82|35.478031|CRAFT BEER|0.0|16|HT CREATE YOUR OWN SAMPLER|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|0.61833652052202714|00072036780300|DOMESTIC BEER|BEER|-80.893784|1.4118628751971085|179|1
35.478031|57853451510da57f8ccea0ce8b5277f680e9d88f|3.49|2015-01-23 14:55:00|80.8939826282094|2|7203688133|179|35.49452270106449|0|2|556|-80.8955|64|35.4437|PACKAGED VEGETABLES|0.0|4|HT FAJITA MIX|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|35.490689277687849|00072036881335|FRESH PRODUCE|PRODUCE|-80.893784|80.893791368780597|272|1
35.478031|09d2e1811cf23c1debabfaa4bcdd348475666c51|13.29|2014-12-08 16:58:00|80.8939826282094|2|3700013882|179|35.49452270106449|0|2|389|-80.8955|66|35.4437|NFS-LAUNDRY DETERGENTS|0.0|1|TIDE HE ORIGINAL|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|35.490689277687849|00037000875888|DETERGENTS|G1 GROCERY|-80.893784|80.893791368780597|272|1
35.478031|c857469a270d8082d4c4a2adc1d346af83386a0d|2.65|2014-09-16 17:48:00|80.8939826282094|2|4530000549|179|35.49452270106449|0|2|125|-80.8955|19|35.4437|PEANUT BUTTER|0.0|1|PETER PAN RF CRNHY PBUTTR|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|35.490689277687849|00045300005393|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.893784|80.893791368780597|272|1
35.478031|1dd7d7da2f0e813d5ba7697960ab734b64aac720|8.99|2015-02-17 16:46:00|80.8939826282094|2|4900003165|179|35.49452270106449|0|2|31|-80.8955|4|35.4437|NON CARBONATED WATER|4.0|1|DASANI .5 LITER 24 PK|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|35.490689277687849|00049000031652|BOTTLED WATER|G1 GROCERY|-80.893784|80.893791368780597|272|1
35.478031|e4f6bb90a90061f6d260c3c395b4c9e96477b84f|3.29|2015-01-20 17:29:00|1.4102725052409182|2|7265546007|179|0.6192084530746164|0|1|1278|-80.893784|48|35.478031|SINGLE SERVE NUTRITIONAL|0.0|5|HC RSTD CHK & POTATO BAKE|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|0.61833652052202714|00072655460034|FROZEN MEALS|FROZEN|-80.893784|1.4118628751971085|179|1
35.478031|5b58214025e889c61cd35cefc6e908df82aa056d|4.49|2014-12-23 12:01:00|80.8939826282094|2|4000031532|179|35.49452270106449|0|2|727|-80.8955|7|35.4437|SEASONAL CANDY-SINGLE FAC|1.49|1|I/O(C14)M&M PLAIN CHRISTMAS|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|35.490689277687849|00040000315322|CANDY|G1 GROCERY|-80.893784|80.893791368780597|272|1
35.478031|6eac57d45a0d71019591c5b52954e44f1bcc6655|3.89|2015-01-12 17:25:00|80.8939826282094|2|7684010015|179|35.494522701825836|0|2|275|-80.861571|45|35.444615|SUPER PREMIUM ICE CREAM|0.0|5|BEN & JERRY FRO YO FDGE BRW|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|35.490689277687849|00076840100569|ICE CREAM|FROZEN|-80.893784|80.893788052598069|340|1
35.478031|fdf558cf858e24cc4a617040494aefb25edb66d1|19.99|2014-10-08 17:52:00|1.4102725052409182|2|4933100230|179|0.6192084530746164|0|1|9976|-80.893784|888|35.478031|NFS-U/PREM-PINOT NOIR|0.0|13|LA CREMA PINOT NOIR|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|0.61833652052202714|00049331002307|ULTRA PREMIUM ($15-$19.99)|WINE|-80.893784|1.4118628751971085|179|1
35.478031|ae88dd1286e2d3465dbb6438a85dc7c376d7328e|6.15|2014-12-01 19:22:00|80.8939826282094|2|20596500000|179|35.494522701825836|0|2|1821|-80.861571|410|35.444615|BH TURKEY|0.0|6|BH OVENGOLD TURKEY - SKINLESS|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|35.490689277687849|00205965000007|BH MEAT|DELI|-80.893784|80.893788052598069|340|1
35.478031|5c373082e7f3b313cbda6823df3c3b60ce017e49|9.98|2015-02-08 16:51:00|80.8939826282094|2|2310027789|179|35.49452270106449|0|2|155|-80.8955|24|35.4437|NFS-DOG TREATS|1.49|1|PEDIGREE DENTASTIX MINI|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|35.490689277687849|00023100277899|PET FOOD/SUPPLIES|G1 GROCERY|-80.893784|80.893791368780597|272|2
35.478031|b4b54a2235b36e7e347577698a4a0a8e6ec66964|16.95|2014-12-22 14:48:00|80.8939826282094|2|76211103168|179|35.49452270106449|0|2|1598|-80.8955|369|35.4437|NFS MERCHANDISE|6.78|22|GOLD GREEN DOT TMBLR HLDY14|836a90942a88a85deb7b738a28894bd0a155ff17|1.1395367929427804|35.490689277687849|00762111031686|NFS STARBUCKS|COFFEE SHOP|-80.893784|80.893791368780597|272|1
35.03469|1c3e663d46787c4c08511265ffb249fd814cc862|8.98|2014-10-22 23:07:00|80.970590786568081|4|61344000003|82|35.077267856220722|0|55|1211|-80.992182|272|35.103409|HISP SALSA/DIPS|0.0|1|CLINTS SALSA MEDIUM|864e22778cd9359b63eae206b0faed24a2797cdf|2.942027603840212|35.077427448337218|00613440000013|HISPANIC PREP. FOODS|G1 GROCERY|-80.97058|80.970612116190694|88|2
35.053394|21ee7273df22a93cc71b69a58049e470c8c4d750|7.07|2015-02-01 13:38:00|80.848351720559364|4|20496000000|11|35.099982697217257|0|25|755|-80.994596|87|35.061685|NFS-BALLOONS|0.0|9|*BALLOONS|8a6f71939c916cd94ae913fb13d7f9e0014d4009|3.2191669972596455|35.082633588753836|00204960000005|FLORAL|FLORAL|-80.848528|80.848560580979537|475|1
35.053394|621ce1e0b9b936798524a4994ca7b113b9bcb678|14.99|2014-11-25 14:12:00|80.848351720559364|4|7314321373|11|35.099982697217257|0|25|7407|-80.994596|1600|35.061685|CHRISTMAS PARTY GOODS/DECOR|5.0|18|I/O DECK THE HALL GLS CUT BRD|8a6f71939c916cd94ae913fb13d7f9e0014d4009|3.2191669972596455|35.082633588753836|00073143213736|SEASONAL MERCHANDISE|GM|-80.848528|80.848560580979537|475|1
35.053394|e306ceec124789193f7b3fcb08c772fb62460543|7.99|2014-12-19 16:30:00|80.848351720559364|4|4145810534|11|35.099982691917425|0|25|265|-80.97058|307|35.03469|FROZEN PIES|3.0|5|EDWARDS CHOC CREAM W/HERSHEY'S|8a6f71939c916cd94ae913fb13d7f9e0014d4009|3.2191669972596455|35.082633588753836|00041458105565|DESSERTS FROZEN|FROZEN|-80.848528|80.84857041278471|82|1
35.053394|56bfaf8b18dbb0399c3b4602d0359444f51d3496|1.69|2014-10-29 13:53:00|80.848351720559364|4|4900000044|11|35.099982673300509|0|25|54|-80.837892|8|34.937113|DIET|0.0|23|CB DIET DR PEPPER 20OZ NR|8a6f71939c916cd94ae913fb13d7f9e0014d4009|3.2191669972596455|35.082633588753836|00078000083408|CARBONATED BEVERAGES|BEVERAGE|-80.848528|80.848594248562506|372|1
35.053394|75f59b5dc0978d2365f2c2b6b18fbc786e6b67a2|2.55|2014-12-24 13:01:00|80.848351720559364|4|7203663996|11|35.099982691917425|0|25|342|-80.97058|57|35.03469|FRESH MILK|0.0|3|HARRIS TEETER WHOLE MILK|8a6f71939c916cd94ae913fb13d7f9e0014d4009|3.2191669972596455|35.082633588753836|00072036639967|MILK|DAIRY|-80.848528|80.84857041278471|82|1
35.053394|f567fabfc335dfed95f3c697e843fd36ba48949a|5.29|2014-10-30 17:11:00|80.848351720559364|4|5150024177|11|35.099982673300509|0|25|125|-80.837892|19|34.937113|PEANUT BUTTER|1.3|1|JIF CREAMY PEANUT BUTTER|8a6f71939c916cd94ae913fb13d7f9e0014d4009|3.2191669972596455|35.082633588753836|00051500241776|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.848528|80.848594248562506|372|1
35.053394|7bb763e6fb3a9015891415e798d01d900e57c5d1|1.69|2014-12-10 12:11:00|80.848351720559364|4|1200000129|11|35.099982673300509|0|25|54|-80.837892|8|34.937113|DIET|0.0|23|CB DIET PEPSI 20 OZ NR|8a6f71939c916cd94ae913fb13d7f9e0014d4009|3.2191669972596455|35.082633588753836|00012000001307|CARBONATED BEVERAGES|BEVERAGE|-80.848528|80.848594248562506|372|1
35.053394|ddb848637156391328211d21b49331292f10ad2e|1.69|2014-12-04 14:47:00|80.848351720559364|4|1200000129|11|35.099982673300509|0|25|54|-80.837892|8|34.937113|DIET|0.0|23|CB DIET PEPSI 20 OZ NR|8a6f71939c916cd94ae913fb13d7f9e0014d4009|3.2191669972596455|35.082633588753836|00012000001307|CARBONATED BEVERAGES|BEVERAGE|-80.848528|80.848594248562506|372|1
35.053394|86bef3a877cf59af0212adf5e44984d9aca76c86|1.69|2014-11-11 11:15:00|80.848351720559364|4|1200000129|11|35.099982673300509|0|25|54|-80.837892|8|34.937113|DIET|0.0|23|CB DIET PEPSI 20 OZ NR|8a6f71939c916cd94ae913fb13d7f9e0014d4009|3.2191669972596455|35.082633588753836|00012000001307|CARBONATED BEVERAGES|BEVERAGE|-80.848528|80.848594248562506|372|1
35.053394|8e9a2b7a2bdc23589171f7af9398d6a0e6151f79|10.17|2014-10-22 10:13:00|80.848351720559364|4|3800031829|11|35.099982673300509|0|25|74|-80.837892|9|34.937113|RTE CEREAL ALL FAMILY|1.7|1|KELL MIN WHEATS BITE SIZE|8a6f71939c916cd94ae913fb13d7f9e0014d4009|3.2191669972596455|35.082633588753836|00038000318290|CEREAL|G1 GROCERY|-80.848528|80.848594248562506|372|3
35.053394|f6811cd1cfda491fa422de429767c659d945b8c3|1.89|2015-02-01 08:31:00|80.848351720559364|4|2700038811|11|35.099982697217257|0|25|257|-80.994596|39|35.061685|TOMATOES|0.0|1|HUNTS TOMATO PASTE 12 OZ.|8a6f71939c916cd94ae913fb13d7f9e0014d4009|3.2191669972596455|35.082633588753836|00027000388112|VEGETABLES-CAN/JAR|G1 GROCERY|-80.848528|80.848560580979537|475|1
35.053394|36550576718270c2d483c15d01c58803e49ff5a4|1.29|2014-12-19 16:32:00|80.848351720559364|4|2200000899|11|35.099982691917425|0|25|48|-80.97058|7|35.03469|REGISTER GUM|0.0|1|EXTRA SPEARMINT|8a6f71939c916cd94ae913fb13d7f9e0014d4009|3.2191669972596455|35.082633588753836|00022000008992|CANDY|G1 GROCERY|-80.848528|80.84857041278471|82|1
35.006282|52e240efe9f099fc091954328c2413a1eef919b8|53.0|2015-01-07 15:56:00|1.4091206135396188|4|20895300000|60|0.6109748797816256|0|47|977|-80.562829|201|35.006282|FRESH HT CHICKEN|6.63|2|HT FRESH BNLS CHICKEN BREAST|905a9b0dccd7f02494c034badeea23eb0b80d8a2|15.168720624842049|0.61242566243833529|00208953000003|POULTRY|MEAT|-80.562829|1.4060866207711706|60|5
35.17739|33f54cd31805b0a02e0e45589aca06435cc8b103|5.99|2015-01-08 17:52:00|80.801203185414451|1|7203688215|208|35.191861823669299|0|24|500|-80.826724|64|35.195689|FRESH APPLES|0.0|4|HT GALA APPLE 5LB|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036882158|FRESH PRODUCE|PRODUCE|-80.80146|80.801461344519637|412|1
35.17739|cbd3a693721c97882b5678c74303103eae699825|2.49|2014-12-21 14:32:00|80.801203185414451|1|7203688130|208|35.191861822752038|0|24|556|-80.825175|64|35.152722|PACKAGED VEGETABLES|0.0|4|HT DICED GREEN PEPPERS|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036881311|FRESH PRODUCE|PRODUCE|-80.80146|80.801466446147188|160|1
35.17739|aa8142b4f7295e5e1cc8526df986afdda2cd126f|20.76|2015-02-04 12:43:00|80.801203185414451|1|7203698020|208|35.191861823657021|0|24|1243|-80.844274|21|35.204336|MIXED NUTS CASHEWS|2.59|1|HT CASHEW HALVES LT SALTED|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036980212|NUTS|G1 GROCERY|-80.80146|80.801461529555027|61|4
35.17739|1359dcbbe25a6e459167bdf24f779e2dacb5d6c3|3.99|2015-01-26 09:43:00|80.801203185414451|1|7203695558|208|35.191861822752038|0|24|2010|-80.825175|500|35.152722|FFM PICKLES|0.0|6|F.F KOSHR DILL SANDWICH SLICE|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036957948|PICKLES|DELI|-80.80146|80.801466446147188|160|1
35.17739|dd5ae791f3b029fbe39af925d51e9c2a6dacbcfb|10.38|2014-11-10 12:29:00|80.801203185414451|1|7203698020|208|35.191861823657021|0|24|1243|-80.844274|21|35.204336|MIXED NUTS CASHEWS|0.0|1|HT CASHEW HALVES LT SALTED|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036980212|NUTS|G1 GROCERY|-80.80146|80.801461529555027|61|2
35.17739|6b9d6a4497e3c023e25137674531fb40a4becbfe|3.49|2014-11-21 10:18:00|80.801203185414451|1|7203698205|208|35.191861823669299|0|24|1250|-80.826724|12|35.195689|SPECIALTY COOKIES|0.49|1|HTT LEMON COOKIE STRAWS|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036982049|COOKIES|G1 GROCERY|-80.80146|80.801461344519637|412|1
35.17739|9af21bbbf82a12787ece9aec03197a6c46277366|10.38|2014-09-22 12:04:00|80.801203185414451|1|7203698020|208|35.191861823657021|0|24|1243|-80.844274|21|35.204336|MIXED NUTS CASHEWS|1.2|1|HT CASHEW HALVES LT SALTED|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036980212|NUTS|G1 GROCERY|-80.80146|80.801461529555027|61|2
35.17739|deb68c43ffde317174d9459af8f5d2c23570ada6|20.76|2015-01-13 11:54:00|80.801203185414451|1|7203698020|208|35.191861823657021|0|24|1243|-80.844274|21|35.204336|MIXED NUTS CASHEWS|2.59|1|HT CASHEW HALVES LT SALTED|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036980212|NUTS|G1 GROCERY|-80.80146|80.801461529555027|61|4
35.17739|1ff0f3300f334e3ec0698d25e5a8d7dd95081af8|5.98|2014-10-06 10:51:00|1.4094857484078087|1|7203697784|208|0.613961277758128|0|26|2020|-80.80146|505|35.17739|CHEESE SPECIALTIES|0.0|6|HT FETA CHEESE CRMBLD|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00072036977847|SPECIALTY CHEESE|DELI|-80.80146|1.4102515174184975|208|2
35.17739|cd36bcfc4dbea14c33185a394594da1b1d2b7d01|4.99|2015-01-12 10:26:00|1.4094857484078087|1|71575620002|208|0.613961277758128|0|26|504|-80.80146|64|35.17739|FRESH BERRIES|2.5|4|STRAWBERRIES 1LB CLAM|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00769197404021|FRESH PRODUCE|PRODUCE|-80.80146|1.4102515174184975|208|1
35.17739|9f72dc8c862569cd0276c18a7d1d54255aaef013|3.9|2014-12-04 10:48:00|1.4094857484078087|1|1450001098|208|0.613961277758128|0|26|1272|-80.80146|50|35.17739|BAG VEG STEAM|0.0|5|BE STEAMFRESH L GRN WHT RICE|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00014500012753|VEGETABLES-FROZEN|FROZEN|-80.80146|1.4102515174184975|208|2
35.17739|92fb2d9f223c2b7bc5adcf626c32312001c46fc3|3.75|2015-01-15 16:14:00|80.801203185414451|1|4139000107|208|35.191861823669299|0|24|79|-80.826724|273|35.195689|ASIAN SAUCES/SEASONINGS|0.0|1|KIKKOMAN SOY SAUCE LT 15|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00041390001079|ASIAN PREP. FOODS|G1 GROCERY|-80.80146|80.801461344519637|412|1
35.17739|adf34087dc297262a9486151e73662d201894d40|7.79|2015-02-09 14:46:00|1.4094857484078087|1|4116709433|208|0.613961277758128|0|26|4035|-80.80146|1080|35.17739|ORAL RINSE-FLOURIDE|0.0|17|ACT MINT RINSE|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00041167094334|ORAL HYGIENE|HBC|-80.80146|1.4102515174184975|208|1
35.17739|dfa3f6beab12abbe94bbd5411a6a89cde4ca79d1|4.49|2014-09-26 12:33:00|80.801203185414451|1|88491201426|208|35.191861822752038|0|24|74|-80.825175|9|35.152722|RTE CEREAL ALL FAMILY|0.0|1|POST HNY BUNCHES FAM HNY RSTD|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00884912014269|CEREAL|G1 GROCERY|-80.80146|80.801466446147188|160|1
35.17739|fd26772e36157ff2b91d9eb0eb974aa06b02e3ed|7.99|2015-01-20 11:41:00|1.4094857484078087|1|1251145124|208|0.613961277758128|0|26|228|-80.80146|36|35.17739|TABLE SYRUP|0.0|1|WHLSM ORGANIC PANCAKE SYRUP.|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00012511451240|TABLE SYRUPS|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|6f369314c4690af70f8b768fe6b90abc90f2389e|4.49|2015-02-25 16:38:00|80.801203185414451|1|88491201426|208|35.191861823657021|0|24|74|-80.844274|9|35.204336|RTE CEREAL ALL FAMILY|0.0|1|POST HNY BUNCHES FAM HNY RSTD|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00884912014269|CEREAL|G1 GROCERY|-80.80146|80.801461529555027|61|1
35.17739|0f1540125e32b19b1e70544eac38db4782d38a37|4.49|2014-09-10 13:54:00|1.4094857484078087|1|88491201426|208|0.613961277758128|0|26|74|-80.80146|9|35.17739|RTE CEREAL ALL FAMILY|0.0|1|POST HNY BUNCHES FAM HNY RSTD|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00884912014269|CEREAL|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|542a2da32c2e7a28c6ba7e10fa95a44ea056fc5f|4.49|2015-03-04 16:52:00|80.801203185414451|1|87989000001|208|35.191861823669299|0|24|1982|-80.826724|480|35.195689|DRY GOODS CRACKERS|0.0|6|ORIGINAL MULTI-SEED CRACKERS|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00879890000014|DRY GOODS|DELI|-80.80146|80.801461344519637|412|1
35.17739|c28a581ffa64fa8a5b2acabcad6fed8423a0123b|4.49|2014-10-22 15:03:00|1.4094857484078087|1|88491201426|208|0.613961277758128|0|26|74|-80.80146|9|35.17739|RTE CEREAL ALL FAMILY|0.0|1|POST HNY BUNCHES FAM HNY RSTD|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00884912014269|CEREAL|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|e8e69934418c31b933baa479db444fcdd5a15a0a|4.49|2014-10-12 14:07:00|80.801203185414451|1|88491201426|208|35.191861822752038|0|24|74|-80.825175|9|35.152722|RTE CEREAL ALL FAMILY|0.0|1|POST HNY BUNCHES FAM HNY RSTD|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00884912014269|CEREAL|G1 GROCERY|-80.80146|80.801466446147188|160|1
35.17739|7b0f73a8072f442e3252157bd7755c0a9facee87|9.99|2014-09-21 16:32:00|1.4094857484078087|1|74052210023|208|0.613961277758128|0|26|458|-80.80146|82|35.17739|CRAFT BEER|0.0|16|BELL'S AMBER ALE 6PK|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00740522100238|DOMESTIC BEER|BEER|-80.80146|1.4102515174184975|208|1
35.17739|7fb6c609147c31f7c9ae7f1fd7501f48d4b22bf8|15.87|2015-01-27 12:23:00|1.4094857484078087|1|71210200100|208|0.613961277758128|0|26|69|-80.80146|26|35.17739|CANNED GRAVY|0.0|1|MORE THAN GOURMET DEMI GLACE|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00712102001006|PREPARED FOODS-DRY MIXES|G1 GROCERY|-80.80146|1.4102515174184975|208|3
35.17739|c4413765f041559b87caffe28058caa2a4da8338|9.99|2015-01-02 17:29:00|80.801203185414451|1|74052210023|208|35.191861823669299|0|24|458|-80.826724|82|35.195689|CRAFT BEER|0.0|16|BELL'S AMBER ALE 6PK|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00740522100238|DOMESTIC BEER|BEER|-80.80146|80.801461344519637|412|1
35.17739|965e3bec754ce1dd86721197fbfcc6c2ac876a2a|2.99|2014-09-15 14:57:00|80.801203185414451|1|20443000000|208|35.191861822752038|0|24|510|-80.825175|64|35.152722|FRESH PINEAPPLE|0.0|4|GOLD PINEAPPLES|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00643126072003|FRESH PRODUCE|PRODUCE|-80.80146|80.801466446147188|160|1
35.17739|e816f8e77aaf7df5ea51c816fd9d851fe94addb0|3.25|2015-01-04 14:45:00|1.4094857484078087|1|7203656080|208|0.613961277758128|0|26|318|-80.80146|52|35.17739|SHREDDED/GRATED CHEESE|0.0|3|HT FANCY SHRED MILD CHED CHES|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00072036560810|CHEESE|DAIRY|-80.80146|1.4102515174184975|208|1
35.17739|8cc416e1e5e8049f9a210b640aa160f235189f22|11.94|2014-11-30 16:47:00|1.4094857484078087|1|7203676359|208|0.613961277758128|0|26|345|-80.80146|57|35.17739|ORGANIC MILK|0.0|3|HTO ORGANIC 1% MILK GAL|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00072036763617|MILK|DAIRY|-80.80146|1.4102515174184975|208|2
35.17739|087933cbe475eb260ea49f40aab85f937ef69259|9.58|2014-09-19 16:35:00|80.801203185414451|1|7203676457|208|35.191861823669299|0|24|312|-80.826724|51|35.195689|BUTTER|0.0|3|HTO ORGANIC BUTTER SALTED|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036763419|BUTTER & MARGARINE|DAIRY|-80.80146|80.801461344519637|412|2
35.17739|cb96cf5ba9549b193853abccf03561fe74841137|3.25|2014-11-02 15:41:00|80.801203185414451|1|7203656080|208|35.191861823669299|0|24|318|-80.826724|52|35.195689|SHREDDED/GRATED CHEESE|0.0|3|HT FANCY SHRED MILD CHED CHES|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036560810|CHEESE|DAIRY|-80.80146|80.801461344519637|412|1
35.17739|4d80f450c6056a3472ff80e81f150cff0f387126|9.75|2014-12-29 17:27:00|80.801203185414451|1|7203656080|208|35.191861823669299|0|24|318|-80.826724|52|35.195689|SHREDDED/GRATED CHEESE|0.0|3|HT FANCY SHRED MILD CHED CHES|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036560810|CHEESE|DAIRY|-80.80146|80.801461344519637|412|3
35.17739|23b7041abc614e62955a6f00582620e0476e7779|3.25|2015-02-19 10:22:00|80.801203185414451|1|7203656080|208|35.191861822752038|0|24|318|-80.825175|52|35.152722|SHREDDED/GRATED CHEESE|0.0|3|HT SHRED SHARP CHED CHEESE 2%|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036590466|CHEESE|DAIRY|-80.80146|80.801466446147188|160|1
35.17739|cb44d3819b49a868d4ee6c2db7ddb9bb788179d1|3.25|2015-02-03 11:48:00|80.801203185414451|1|7203656080|208|35.191861823669299|0|24|318|-80.826724|52|35.195689|SHREDDED/GRATED CHEESE|0.0|3|HT SHRED SHARP CHED CHEESE 2%|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036590466|CHEESE|DAIRY|-80.80146|80.801461344519637|412|1
35.17739|99ac11954a08c8b584b10c2548007d4527d5f311|2.69|2014-10-20 10:06:00|80.801203185414451|1|7203688023|208|35.191861822752038|0|24|555|-80.825175|64|35.152722|PACKAGED SALADS|0.0|4|HT CURLY SPINACH,PKG|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036880239|FRESH PRODUCE|PRODUCE|-80.80146|80.801466446147188|160|1
35.17739|085ef2dc973886e41e185c19eb98b9b226e44293|5.49|2015-01-24 14:38:00|1.4094857484078087|1|4900000548|208|0.613961277758128|0|26|55|-80.80146|8|35.17739|REGULAR|0.5|23|SPRITE 12OZ PET8PK FRIDGEPK|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00049000006124|CARBONATED BEVERAGES|BEVERAGE|-80.80146|1.4102515174184975|208|1
35.17739|c3cdae56023c75f31328f2351bade9f01fe712c4|1.15|2014-09-21 14:34:00|80.801203185414451|1|4920005675|208|35.191861823669299|0|24|224|-80.826724|35|35.195689|SUGAR-BROWN|0.0|1|DOMINO LT BRWN SUGAR-BOX|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00049200056752|SUGAR/SUBSTITUTES|G1 GROCERY|-80.80146|80.801461344519637|412|1
35.17739|c9eb27c06b6dcba38129db989b400b2a20230806|1.49|2015-01-06 16:04:00|1.4094857484078087|1|2840002819|208|0.613961277758128|0|26|206|-80.80146|31|35.17739|FRONT END SNACKS|0.0|1|LAYS BBQ|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00028400025904|SNACKS|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|3ede8baae5285ee4818824721ec441bbd2e7543b|1.5|2014-12-09 13:11:00|1.4094857484078087|1|7203670990|208|0.613961277758128|0|26|22|-80.80146|28|35.17739|CROUTONS|0.5|1|HT CROUTONS SEASONED|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00072036709905|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|ef6ea92a9f295ce6719712e4e55abdabcaea847c|5.23|2014-10-16 08:38:00|80.801203185414451|1||208|35.191861822752038|0|24|500|-80.825175|64|35.152722|FRESH APPLES|1.97|4|HONEY CRISP APPLE|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00233283000003|FRESH PRODUCE|PRODUCE|-80.80146|80.801466446147188|160|1
35.17739|82a7edafb05ac78c299fab60d45141ece9a26eb4|2.17|2014-12-17 15:32:00|80.801203185414451|1|7203631017|208|35.191861822752038|0|24|1245|-80.825175|34|35.152722|SINGLE SPICES|0.0|1|E  HT CHILI POWDER|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036310170|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.80146|80.801466446147188|160|1
35.17739|7ae022ea0064a615035025dc3887449842261c57|1.7999999999999998|2015-02-01 15:43:00|1.4094857484078087|1|7047000100|208|0.613961277758128|0|26|687|-80.80146|61|35.17739|BLENDED|0.0|3|YOPLAIT STRAWBERRY CUSTARD|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00070470001005|YOGURT|DAIRY|-80.80146|1.4102515174184975|208|3
35.17739|c37a6d5c0e1a7c0b4c1de7dee4533b014291160f|5.19|2015-01-03 19:42:00|80.801203185414451|1|1204401560|208|35.191861823669299|0|24|3816|-80.826724|1070|35.195689|INVISIBLE-MALE|1.2|17|O.S. FRESH COLL AP/DEO DENALI|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00012044015612|DEODORANT|HBC|-80.80146|80.801461344519637|412|1
35.17739|27b58439cefa456f99b3fe890f38abbc776d8175|2.99|2014-10-27 17:39:00|80.801203185414451|1|7203695121|208|35.191861823306901|0|24|1629|-80.85013|373|35.175855|TAKE & BAKE ROLLS|0.0|14|TAKE & BAKE WHEAT PETIT PN RL|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036951212|ROLLS|BAKERY|-80.80146|80.801464184541501|218|1
35.17739|6cf732203301c45924e99fdefdec148d21f0d686|5.69|2015-03-02 12:15:00|80.801203185414451|1|7203633086|208|35.191861823657021|0|24|1148|-80.844274|21|35.204336|ALMONDS|1.21|1|HT ROASTED ALMONDS LIGHT SALT|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036979537|NUTS|G1 GROCERY|-80.80146|80.801461529555027|61|1
35.17739|3fec72d82f70bff0d4d9eeeefcd1e1fb7a99e604|2.99|2014-10-04 21:43:00|80.801203185414451|1|7203695678|208|35.191861823669299|0|24|1677|-80.826724|383|35.195689|INDIVIDUALS (PASTRY CASE)|0.0|14|FFM COCONUT CREAM PIE MINI|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036957658|PASTRY CASE|BAKERY|-80.80146|80.801461344519637|412|1
35.17739|3cad1783ea0d623eac3d9778b92e8743659018e1|8.98|2014-11-06 09:39:00|80.801203185414451|1|7203695755|208|35.191861822752038|0|24|1647|-80.825175|379|35.152722|PACKAGED MUFFINS|0.0|14|12CT MINI BLUEBERRY MUFFINS|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036957559|MUFFINS|BAKERY|-80.80146|80.801466446147188|160|2
35.17739|3cede6129faf7a0b18531efee9b794d46187d95d|4.89|2014-12-28 19:41:00|80.801203185414451|1|7365111709|208|35.191861822752038|0|24|160|-80.825175|25|35.152722|OLIVES|1.39|1|MARIO OLIVE MANZ 13.|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00073651117090|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.80146|80.801466446147188|160|1
35.17739|bb152c680d7486da23fc567e2e2a94e43a609a43|3.25|2015-03-01 19:35:00|1.4094857484078087|1|7203656080|208|0.613961277758128|0|26|318|-80.80146|52|35.17739|SHREDDED/GRATED CHEESE|0.0|3|HT FANCY SHRED MEXICAN CHS 2%|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00072036560827|CHEESE|DAIRY|-80.80146|1.4102515174184975|208|1
35.17739|c4f25e09e7ba77898ed8c0face7e21fe48b8e1d0|3.09|2014-10-13 18:17:00|80.801203185414451|1|7225002313|208|35.191861823669299|0|24|1033|-80.826724|163|35.195689|HAMBURGER|0.0|7|NATOWN 8PK BUTTER HAMS|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072250023139|BUNS/ROLLS|COMMERCIAL BAKERY|-80.80146|80.801461344519637|412|1
35.17739|5993fe7c7dd99e585ca28bfbe69d598aef86d811|11.58|2014-11-24 09:11:00|1.4094857484078087|1|20193000000|208|0.613961277758128|0|26|299|-80.80146|49|35.17739|ANGUS BEEF|0.0|2|ANGUS BEEF CHUCK TENDER ROAST|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00201930000003|BEEF|MEAT|-80.80146|1.4102515174184975|208|1
35.17739|9d96d84dbdb1089816a16290dd781e00766d9a95|9.87|2015-01-30 14:49:00|80.801203185414451|1|7203644036|208|35.191861823669299|0|24|273|-80.826724|43|35.195689|PREMIUM NOVELTIES|0.0|5|HT MINI ICE CREAM SANDWICH|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036460479|FROZEN NOVELTIES|FROZEN|-80.80146|80.801461344519637|412|3
35.17739|37acf80458bfce5c736a7f78daa52d4c3bb2421d|9.99|2014-09-29 17:01:00|80.801203185414451|1|7826407706|208|35.191861823306901|0|24|583|-80.85013|136|35.175855|NUTS|0.0|4|HT PINE NUTS TRAY, 6 OZ|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00078264077069|OTHER MERCHANDISE|PRODUCE|-80.80146|80.801464184541501|218|1
35.17739|7a50d2dfa644cc24db0432533ab806af604751ef|4.99|2014-09-28 18:44:00|80.801203185414451|1|7203695714|208|35.191861823306901|0|24|1647|-80.85013|379|35.175855|PACKAGED MUFFINS|1.02|14|JUMBO LEM POPPY MUFFIN 4 CT.|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036957184|MUFFINS|BAKERY|-80.80146|80.801464184541501|218|1
35.17739|eaf9ce14dbd6d654b3ac7ad59b43195784c0f1f1|4.99|2014-12-19 11:03:00|1.4094857484078087|1|7447034190|208|0.613961277758128|0|26|6785|-80.80146|1568|35.17739|MAGAZINES WEEKLY|0.0|18|US WEEKLY|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00074470341901|MAGAZINES|GM|-80.80146|1.4102515174184975|208|1
35.17739|ad9a5f2bae8d7c9e78a17787b084a6c4fa590f11|8.69|2014-10-20 13:19:00|80.801203185414451|1|7203653118|208|35.191861822752038|0|24|1243|-80.825175|21|35.152722|MIXED NUTS CASHEWS|2.7|1|HT CASHEWS HALVES|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036531186|NUTS|G1 GROCERY|-80.80146|80.801466446147188|160|1
35.17739|4768e9eacba1e524dee705b807ae87608c5eb289|4.98|2015-01-28 16:01:00|80.801203185414451|1||208|35.191861823669299|0|24|561|-80.826724|64|35.195689|FR PROD ORGANIC PRODUCE|0.49|4|ORG HASS AVOCADOS|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00294225000000|FRESH PRODUCE|PRODUCE|-80.80146|80.801461344519637|412|2
35.17739|83244cda3c98fc00173e33541413d7e531897021|39.98|2014-11-09 17:51:00|80.801203185414451|1|66957601926|208|35.191861823669299|0|24|9972|-80.826724|888|35.195689|NFS-U/PREM-CAB SAUVIGNON|0.0|13|DUCKHORN DECOY CAB SAUV|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00669576019269|ULTRA PREMIUM ($15-$19.99)|WINE|-80.80146|80.801461344519637|412|2
35.17739|b4ee3e29c71b27c079562005d208d7b3ee8caf3f|7.38|2015-02-23 17:12:00|80.801203185414451|1|61144334026|208|35.191861823306901|0|24|214|-80.85013|33|35.175855|BROTH|0.0|1|KITCHEN BASICS STOCK BEEF|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00611443340112|SOUP|G1 GROCERY|-80.80146|80.801464184541501|218|2
35.17739|087f116d54221fb9769781d797dc32d5d55e7cdf|17.99|2015-02-22 17:16:00|80.801203185414451|1|8841578405|208|35.191861823669299|0|24|9971|-80.826724|888|35.195689|NFS-U/PREM-CHARDONNAY|0.0|13|CB-SIMI CHARDONNAY|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00088415784050|ULTRA PREMIUM ($15-$19.99)|WINE|-80.80146|80.801461344519637|412|1
35.17739|760bb2f3e0d04942b3191634e93a687c382ed371|34.99|2014-09-17 16:49:00|1.4094857484078087|1|4667745185|208|0.613961277758128|0|26|6156|-80.80146|1546|35.17739|BULB-L.E.D. LIGHTING|0.0|18|PHLPS LED 8W BRIGHT WHITE|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00046677426118|LIGHT BULBS/ELECTRICAL|GM|-80.80146|1.4102515174184975|208|1
35.17739|3b974b32cbf61133375904dd248490d280c4a111|6.99|2014-11-10 14:31:00|1.4094857484078087|1|67043309410|208|0.613961277758128|0|26|1419|-80.80146|201|35.17739|SMART CHICKEN ORGANIC|0.0|2|SMART ORGANIC GROUND CHICKEN|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00670433094107|POULTRY|MEAT|-80.80146|1.4102515174184975|208|1
35.17739|045ce9ec24dbc24184f1d19c71c9a93431cfa2b9|6.99|2015-02-08 17:53:00|1.4094857484078087|1|67043309410|208|0.613961277758128|0|26|1419|-80.80146|201|35.17739|SMART CHICKEN ORGANIC|0.0|2|SMART ORGANIC GROUND CHICKEN|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00670433094107|POULTRY|MEAT|-80.80146|1.4102515174184975|208|1
35.17739|1f973c82f31b9a27ccef350f5fcf14b7c82238c8|1.65|2014-10-18 19:11:00|80.801203185414451|1|20892500000|208|35.191861823669299|0|24|658|-80.826724|137|35.195689|FRESH PORK SAUSAGE|0.0|2|PORK ITALIAN SWEET SAUSAGE|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00208925000000|PORK|MEAT|-80.80146|80.801461344519637|412|1
35.17739|0a7e21911d975d5c474a21d86b8541b86509bb3a|4.99|2015-01-30 18:10:00|1.4094857484078087|1|7800000119|208|0.613961277758128|0|26|55|-80.80146|8|35.17739|REGULAR|1.0|23|CANADA DRY CLUB SODA 10 OZ|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00078000001198|CARBONATED BEVERAGES|BEVERAGE|-80.80146|1.4102515174184975|208|1
35.17739|cf9c4b8f1272ab662405dca8d731eeef57f566f2|3.99|2014-09-27 19:58:00|80.801203185414451|1|7684010015|208|35.191861823669299|0|24|275|-80.826724|45|35.195689|SUPER PREMIUM ICE CREAM|0.0|5|BEN & JERRY RED VELVET CAKE|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00076840128358|ICE CREAM|FROZEN|-80.80146|80.801461344519637|412|1
35.17739|100a2aa9fc27b62d0c6a3eaee6a1c157af6a38e2|4.19|2014-12-02 12:05:00|1.4094857484078087|1|4812110208|208|0.613961277758128|0|26|1037|-80.80146|164|35.17739|ENGLISH MUFFINS|2.1|7|THOMAS ENG MUFFN ORIG 6 PK PP|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00048121102081|BREAKFAST|COMMERCIAL BAKERY|-80.80146|1.4102515174184975|208|1
35.17739|21c96c94d48f64f18c162001523344b771ded0e2|2.69|2014-09-23 13:45:00|80.801203185414451|1|5000032822|208|35.191861823669299|0|24|341|-80.826724|57|35.195689|CREAMERS|0.0|3|COFFEE-MATE HAZLENUT|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00050000328222|MILK|DAIRY|-80.80146|80.801461344519637|412|1
35.17739|a5d1ccc640b0420200cefa9cf5f6f9c556175a5c|5.97|2014-10-02 15:13:00|1.4094857484078087|1|7203676359|208|0.613961277758128|0|26|345|-80.80146|57|35.17739|ORGANIC MILK|0.0|3|HTO ORGANIC FF SKIM GAL|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00072036763624|MILK|DAIRY|-80.80146|1.4102515174184975|208|1
35.17739|15fe32662c133a28715c508b4ca2d9c586ced19a|4.29|2014-12-10 16:13:00|80.801203185414451|1|2840006399|208|35.191861823669299|0|24|204|-80.826724|31|35.195689|TORTILLA CHIPS|1.29|1|TOSTITOS BITES|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00028400064057|SNACKS|G1 GROCERY|-80.80146|80.801461344519637|412|1
35.17739|aed62cb4f5143894872f79b5565ba04155b059af|1.99|2014-12-24 10:51:00|80.801203185414451|1|88596708120|208|35.191861823669299|0|24|422|-80.826724|71|35.195689|NFS-REMAIN LAUNDRY SUPPL|0.0|1|NIAGARA STARCH|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00885967081206|LAUNDRY SUPPLIES|G1 GROCERY|-80.80146|80.801461344519637|412|1
35.17739|aab6ae6934d87af907604e6be678fcfed5779e0f|3.49|2014-11-12 10:16:00|1.4094857484078087|1|2840008294|208|0.613961277758128|0|26|201|-80.80146|31|35.17739|POTATO CHIPS|0.99|1|LAYS KETTLE SALT & VINEGAR|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00028400082921|SNACKS|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|c173047a14edb3c66d21835d696a8b926d999751|5.39|2015-03-07 10:11:00|80.801203185414451|1|7027200217|208|35.191861823669299|0|24|1132|-80.826724|55|35.195689|EGGS SUBSTITUTES|0.0|3|EGGBEATER CARTON 32|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00070272002170|EGGS FRESH|DAIRY|-80.80146|80.801461344519637|412|1
35.17739|32433f37b3af5042d0837427b7f86584ca2bb357|3.39|2015-01-16 19:15:00|80.801203185414451|1|61300873513|208|35.191861819785494|0|24|99|-80.824767|32|35.116751|LIQUID TEA|0.6|1|ARIZONA DIET PEACH TEA GALLON|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00613008719760|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.80146|80.801473042011608|294|1
35.17739|3677ea2ee88b6d5a5538d6f6ccd83a620b262869|4.69|2014-11-16 12:32:00|1.4094857484078087|1|7047046158|208|0.613961277758128|0|26|685|-80.80146|61|35.17739|GREEK|1.35|3|YOPLAIT GRK 100 MIX BERRY 4PK|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00070470455914|YOGURT|DAIRY|-80.80146|1.4102515174184975|208|1
35.17739|711c9a6d469cc83e4e178e311a2bc227800221e6|8.79|2015-02-17 15:55:00|1.4094857484078087|1|20597600000|208|0.613961277758128|0|26|1821|-80.80146|410|35.17739|BH TURKEY|0.0|6|BOARS HEAD GOLDEN CATERING TRK|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|0.61471665291522548|00205976000003|BH MEAT|DELI|-80.80146|1.4102515174184975|208|1
35.17739|47c8d6cacebd3b5ffa0d658ca0d2f775dfc3c25d|5.99|2014-10-28 10:05:00|80.801203185414451|1|7356100924|208|35.191861822752038|0|24|7632|-80.825175|1630|35.152722|HOUSE PLANT FOOD|0.0|18|M/GRO SHK N FEED ALL PURP PLNT|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00073561009249|INDOOR PLANT CARE|GM|-80.80146|80.801466446147188|160|1
35.17739|72891b1d246621428252e5076ae766cb328e31b7|2.49|2015-01-21 17:30:00|80.801203185414451|1|4156514116|208|35.191861819785494|0|24|1211|-80.824767|272|35.116751|HISP SALSA/DIPS|0.0|1|PACE REST SALSA MED|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00041565193882|HISPANIC PREP. FOODS|G1 GROCERY|-80.80146|80.801473042011608|294|1
35.17739|6df0583d74d0c96fd9438ba8b9d0a5458f1a00c6|1.99|2015-02-11 18:14:00|80.801203185414451|1|1130010497|208|35.191861819785494|0|24|727|-80.824767|7|35.116751|SEASONAL CANDY-SINGLE FAC|0.74|1|I/O(V15)BRACH SM CONV HEARTS|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00011300104978|CANDY|G1 GROCERY|-80.80146|80.801473042011608|294|1
35.17739|c10c3a871829606144a6482d053fa7e82cb0b6e9|4.81|2014-10-30 09:12:00|80.801203185414451|1||208|35.191861819785494|0|24|502|-80.824767|64|35.116751|FRESH BANANAS|0.0|4|BANANAS, YELLOW|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00204011000008|FRESH PRODUCE|PRODUCE|-80.80146|80.801473042011608|294|1
35.17739|d2f66d9310ef6ca8aeb78ed79233e6d1ba89e3e3|6.27|2014-09-11 14:51:00|80.801203185414451|1||208|35.191861823669299|0|24|502|-80.826724|64|35.195689|FRESH BANANAS|0.0|4|BANANAS, YELLOW|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00204011000008|FRESH PRODUCE|PRODUCE|-80.80146|80.801461344519637|412|2
35.17739|f481162d176f509808c8b4fafa385fdb353067e4|10.0|2015-02-20 20:09:00|80.801203185414451|1|20564800000|208|35.191861822752038|0|24|1945|-80.825175|465|35.152722|SUPERFLAG CHEF CASE|0.0|6|TWICE BAKED POTATOES W/HAM|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00205648000003|COLD PREPARED FOODS|DELI|-80.80146|80.801466446147188|160|1
35.17739|a3cfc12b7d1817cc4ba943859331634aa3a44723|22.99|2014-11-20 18:29:00|80.801203185414451|1|69874390750|208|35.191861823669299|0|24|9985|-80.826724|890|35.195689|NFS-LUX-CAB SAUVIGNON|0.0|13|ROTH ESTATE CABERNET|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00698743907504|LUXURY (OVER $20)|WINE|-80.80146|80.801461344519637|412|1
35.17739|d8f33eade59be6d0c72ed2f67f817838d93d0683|25.0|2014-12-23 12:51:00|80.801203185414451|1|1030093302|208|35.191861823657021|0|24|1243|-80.844274|21|35.204336|MIXED NUTS CASHEWS|1.76|1|EMERALD DELUXE MIXED NUTS|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00010300536222|NUTS|G1 GROCERY|-80.80146|80.801461529555027|61|4
35.17739|6b073065aae2c428fb586fe07afb7d2ee5bc1ff0|7.49|2014-10-28 09:51:00|80.801203185414451|1|3800077259|208|35.191861819785494|0|24|43|-80.824767|6|35.116751|INSTANT BREAKFAST-POWDERED|0.0|1|KELL TGO BRKFST SHK MILK CHOC|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00038000772573|BREAKFAST FOODS|G1 GROCERY|-80.80146|80.801473042011608|294|1
35.17739|f92cd2be79567e34995538d8d56a838c77db5032|9.98|2014-12-12 13:47:00|80.801203185414451|1|7203698017|208|35.191861823657021|0|24|1243|-80.844274|21|35.204336|MIXED NUTS CASHEWS|0.5|1|HT MIX NUTS LT SALT|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036980182|NUTS|G1 GROCERY|-80.80146|80.801461529555027|61|2
35.17739|589fc1c9670d7946ae763fdb61b151427c0ef851|9.19|2015-01-20 16:18:00|80.801203185414451|1|7910090244|208|35.191861822553221|0|24|155|-80.810056|24|35.219587|NFS-DOG TREATS|0.0|1|MILK-BONE FLAVOR SNACKS ECONO|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00079100822393|PET FOOD/SUPPLIES|G1 GROCERY|-80.80146|80.80146708290944|401|1
35.17739|f7cc89858306243e0c6c6a46f9ae08a0ad1bbe3c|4.59|2015-02-24 12:32:00|80.801203185414451|1|7203670570|208|35.191861823657021|0|24|1149|-80.844274|21|35.204336|PEANUTS|0.6|1|HT TRADER SALTED VIRGINIA PNT|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00072036705709|NUTS|G1 GROCERY|-80.80146|80.801461529555027|61|1
35.17739|d769d920c3a3f2d1b5e19e5399a20678547e5b82|25.96|2014-10-02 12:43:00|80.801203185414451|1|2900001669|208|35.191861823657021|0|24|1243|-80.844274|21|35.204336|MIXED NUTS CASHEWS|0.0|1|PLANTERS MIXED NUTS LT SALT|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00029000016699|NUTS|G1 GROCERY|-80.80146|80.801461529555027|61|4
35.17739|5212e0e9a446897c156ed4cbe5762798d2bcc81a|19.99|2014-09-25 17:45:00|80.801203185414451|1|1951822043|208|35.191861823669299|0|24|742|-80.826724|87|35.195689|"NFS-BLOOMING 4"""|0.0|9|"5"" PHAL. ORCHID IN CERAMIC"|924566a1487df9f3778654dd1c6f116aa0af2b5e|0.9999680702282295|35.194272495053255|00019518220435|FLORAL|FLORAL|-80.80146|80.801461344519637|412|1
35.024464|149cb54a438080216436d7460fdb367906c93487|3.39|2015-02-16 11:48:00|1.41290891556208|1|7203646021|317|0.6112922155462233|0|33|1463|-80.847383|42|35.024464|REGULAR FROZEN FRUIT|0.39|5|HT BERRY MEDLEY|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00072036460622|FROZEN FRUIT|FROZEN|-80.847383|1.4110530249708906|317|1
35.024464|03aa3a1366123d9bd40896e9792a8f2cfc23c8e7|3.99|2014-12-03 10:32:00|1.41290891556208|1|7127927100|317|0.6112922155462233|0|33|555|-80.847383|64|35.024464|PACKAGED SALADS|0.99|4|F.E. BABY SPINACH|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00071279271002|FRESH PRODUCE|PRODUCE|-80.847383|1.4110530249708906|317|1
35.024464|75bbe1805c878bf6ff5c0bf696de947b11716cc5|1.25|2015-03-05 10:43:00|1.41290891556208|1|7203624020|317|0.6112922155462233|1|33|149|-80.847383|23|35.024464|WHSE PASTA CORE|0.0|1|HT PASTA ORZO|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00072036240248|PASTA|G1 GROCERY|-80.847383|1.4110530249708906|317|1
35.024464|926faea66c5665ae9356e130837c886f9416bd77|4.29|2014-12-10 09:18:00|1.41290891556208|1|2898905534|317|0.6112922155462233|1|33|286|-80.847383|194|35.024464|MEATLESS|0.96|5|MSF MED VEGGIE BURGER|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00028989759849|MEATLESS-FROZEN|FROZEN|-80.847383|1.4110530249708906|317|1
35.024464|ebdc011ca7811ff4d88d13aac2e52cbdfa026046|4.39|2014-10-05 11:25:00|1.41290891556208|1|2898905534|317|0.6112922155462233|0|33|286|-80.847383|194|35.024464|MEATLESS|0.89|5|MSF MED VEGGIE BURGER|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00028989759849|MEATLESS-FROZEN|FROZEN|-80.847383|1.4110530249708906|317|1
35.024464|6cd54f02ed48ccac63282dada4ab044b3012a13d|4.25|2015-02-19 10:52:00|1.41290891556208|1|2898997310|317|0.6112922155462233|1|33|286|-80.847383|194|35.024464|MEATLESS|0.0|5|MSF  BRKFAST LINKS|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00028989971104|MEATLESS-FROZEN|FROZEN|-80.847383|1.4110530249708906|317|1
35.024464|dc8c1b98fede4a21e2a3fed9fd6d6be74150af44|1.25|2015-01-07 08:48:00|1.41290891556208|1|2400016286|317|0.6112922155462233|1|33|245|-80.847383|39|35.024464|VEGETABLES-CORE|0.25|1|DEL MONTE CORN WK NS|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00024000163053|VEGETABLES-CAN/JAR|G1 GROCERY|-80.847383|1.4110530249708906|317|1
35.024464|a984daba62621294b6957569beebaaeb2a41e50e|1.25|2014-12-06 09:52:00|80.811922674510953|1|2400016286|317|35.032960594179002|0|12|245|-80.8062|39|35.037115|VEGETABLES-CORE|0.25|1|DEL MONTE CORN WK NS|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|35.037868710371079|00024000163053|VEGETABLES-CAN/JAR|G1 GROCERY|-80.847383|80.847386296408544|27|1
35.024464|54aa88290b2ec261c6961d3a23c2f07298d2aebd|4.29|2014-12-26 11:29:00|1.41290891556208|1|2840016014|317|0.6112922155462233|0|33|201|-80.847383|31|35.024464|POTATO CHIPS|0.29|1|LAYS WAVY REGULAR|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00028400160209|SNACKS|G1 GROCERY|-80.847383|1.4110530249708906|317|1
35.024464|9ba697b96bbf1764ec0154dfd0c3ce96c5380cd6|2.79|2015-01-26 12:07:00|1.41290891556208|1|4144930022|317|0.6112922155462233|0|33|8|-80.847383|2|35.024464|BROWNIE MIXES|0.0|1|GHIRADELLI SYRUP BROWNIE|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00041449302546|BAKING MIXES|G1 GROCERY|-80.847383|1.4110530249708906|317|1
35.024464|d0fb2dcc6565658b2b082498f4aa2ca19d412bdb|2.89|2014-10-15 11:28:00|1.41290891556208|1|4400000055|317|0.6112922155462233|0|33|88|-80.847383|13|35.024464|FLAKED SODA CRACKERS|0.0|1|NABISCO PREMIUMS|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00044000000578|CRACKERS|G1 GROCERY|-80.847383|1.4110530249708906|317|1
35.024464|d0bafb0cc1988ef30ee6691416d81e0ad85a063a|5.58|2014-09-11 14:45:00|1.41290891556208|1|4144930022|317|0.6112922155462233|0|33|8|-80.847383|2|35.024464|BROWNIE MIXES|0.0|1|GHIRADELLI ULTIMATE FUDGE BRWN|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00041449302645|BAKING MIXES|G1 GROCERY|-80.847383|1.4110530249708906|317|2
35.024464|ad2be20d997e1b10eec4254c1d131f375e4943bf|4.99|2015-01-20 09:01:00|1.41290891556208|1|4082201114|317|0.6112922155462233|1|33|1878|-80.847383|435|35.024464|HUMMUS|2.5|6|HUMMUS W/ ROASTED PINE NUTS|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00040822011747|SALADS|DELI|-80.847383|1.4110530249708906|317|1
35.024464|1d80a19242a5921c6d90836c2503de810f799b80|1.29|2014-11-06 08:42:00|1.41290891556208|1|3940001810|317|0.6112922155462233|1|33|242|-80.847383|39|35.024464|CANNED BEANS|0.29|1|BUSH BEAN RS GRT NORTHERN|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00039400017790|VEGETABLES-CAN/JAR|G1 GROCERY|-80.847383|1.4110530249708906|317|1
35.024464|ba4ff4d4bda808aea303f9c44b862c916e9af3a7|19.96|2014-12-13 16:19:00|1.41290891556208|1|4082201114|317|0.6112922155462233|0|33|1878|-80.847383|435|35.024464|HUMMUS|0.0|6|ROASTED RED PEPPER HUMMUS|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00040822011549|SALADS|DELI|-80.847383|1.4110530249708906|317|4
35.024464|9b58bd37f3a14cc67d45d82418b279ab9b218e50|4.99|2014-09-18 19:53:00|1.41290891556208|1|4082201114|317|0.6112922155462233|0|33|1878|-80.847383|435|35.024464|HUMMUS|2.5|6|ROASTED RED PEPPER HUMMUS|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00040822011549|SALADS|DELI|-80.847383|1.4110530249708906|317|1
35.024464|d3b1cd6a562812e4cb37d084e842e0cd71656b9f|6.15|2014-10-25 08:08:00|1.41290891556208|1||317|0.6112922155462233|1|33|536|-80.847383|64|35.024464|FRESH SQUASH|2.55|4|BUTTERNUT SQUASH|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00204759000001|FRESH PRODUCE|PRODUCE|-80.847383|1.4110530249708906|317|1
35.024464|c7efd1dfe9b8a9dfd05303ba2e66cf55698202fa|4.19|2014-10-30 14:38:00|1.41290891556208|1||317|0.6112922155462233|0|33|536|-80.847383|64|35.024464|FRESH SQUASH|0.99|4|BUTTERNUT SQUASH|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00204759000001|FRESH PRODUCE|PRODUCE|-80.847383|1.4110530249708906|317|1
35.024464|00b5407ad8fccb819d87f4ba970a097a94c6c430|8.0|2015-01-24 12:42:00|1.41290891556208|1||317|0.6112922155462233|0|33|511|-80.847383|64|35.024464|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00204770000004|FRESH PRODUCE|PRODUCE|-80.847383|1.4110530249708906|317|4
35.024464|41946481cc0606a0e23158c6d011776ffad1b901|6.01|2014-12-20 12:38:00|1.41290891556208|1||317|0.6112922155462233|0|33|500|-80.847383|64|35.024464|FRESH APPLES|0.6|4|BRAEBURN APPLES|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00204103000008|FRESH PRODUCE|PRODUCE|-80.847383|1.4110530249708906|317|1
35.024464|f5e4cd77b1a1556b5a68110586769d1d8849e8e2|6.0|2014-12-15 16:44:00|1.41290891556208|1||317|0.6112922155462233|0|33|511|-80.847383|64|35.024464|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00204770000004|FRESH PRODUCE|PRODUCE|-80.847383|1.4110530249708906|317|3
35.024464|b66ca726b2731e95e22907920d099aa83a10ce58|6.0|2014-11-15 14:47:00|1.41290891556208|1||317|0.6112922155462233|0|33|511|-80.847383|64|35.024464|FRESH AVOCADOS|0.21|4|AVOCADOS, HASS XL 36CT|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00204770000004|FRESH PRODUCE|PRODUCE|-80.847383|1.4110530249708906|317|3
35.024464|1c395e8665244f8a45a126050c96192f5105a136|6.0|2014-12-24 14:50:00|1.41290891556208|1||317|0.6112922155462233|0|33|511|-80.847383|64|35.024464|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00204770000004|FRESH PRODUCE|PRODUCE|-80.847383|1.4110530249708906|317|3
35.024464|afa66609b4129240a423c8c99fade3154677824d|4.0|2014-09-30 10:33:00|1.41290891556208|1||317|0.6112922155462233|0|33|511|-80.847383|64|35.024464|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00204770000004|FRESH PRODUCE|PRODUCE|-80.847383|1.4110530249708906|317|2
35.024464|b5533e06eaddc5467b3f6f316449c88e0386c45d|4.0|2014-09-12 14:44:00|1.41290891556208|1||317|0.6112922155462233|0|33|511|-80.847383|64|35.024464|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00204770000004|FRESH PRODUCE|PRODUCE|-80.847383|1.4110530249708906|317|2
35.024464|771e13e627ce19400bfb8b38c7d04b5239c104af|2.0|2014-09-16 14:09:00|1.41290891556208|1||317|0.6112922155462233|0|33|511|-80.847383|64|35.024464|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00204770000004|FRESH PRODUCE|PRODUCE|-80.847383|1.4110530249708906|317|1
35.024464|b82c0cf69d3d19ff76af36c20b2b1d9a62759319|8.0|2015-02-04 09:00:00|1.41290891556208|1||317|0.6112922155462233|1|33|511|-80.847383|64|35.024464|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00204770000004|FRESH PRODUCE|PRODUCE|-80.847383|1.4110530249708906|317|4
35.024464|fbbb66260f0a2c3e9f2b16965f31fdfb799c079c|1.95|2015-02-02 15:11:00|1.41290891556208|1|64420941000|317|0.6112922155462233|0|33|10|-80.847383|2|35.024464|LAYER CAKE MIX|0.0|1|D HINES DEVIL FOOD CAKE MIX|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00644209410408|BAKING MIXES|G1 GROCERY|-80.847383|1.4110530249708906|317|1
35.024464|adcb2495fd2c8d6b469d51a41e25715ebd77252b|5.99|2014-12-22 21:05:00|1.41290891556208|1|7203676140|317|0.6112922155462233|0|33|239|-80.847383|38|35.024464|RICE-PACKAGED & BULK|1.0|1|HT TRADER RICE WILD BLEND|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00072036761446|RICE GRAINS AND BEANS|G1 GROCERY|-80.847383|1.4110530249708906|317|1
35.024464|2faca1db7813d12119b4f81651f30d79ff595ce7|1.98|2015-03-08 11:04:00|1.41290891556208|1|7203676439|317|0.6112922155462233|0|33|242|-80.847383|39|35.024464|CANNED BEANS|0.0|1|HTO BEAN BLACK|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00072036764416|VEGETABLES-CAN/JAR|G1 GROCERY|-80.847383|1.4110530249708906|317|2
35.024464|f5deafaee7f0396d52f8e1e32b7a3e56c0fdefad|2.79|2015-03-03 21:38:00|1.41290891556208|1|7203671028|317|0.6112922155462233|0|33|62|-80.847383|7|35.024464|SPECIALTY BAR/BOX CHOCOLATE|0.29|1|HT TRDRS CARM&S SALT MLK CHOC|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00072036710284|CANDY|G1 GROCERY|-80.847383|1.4110530249708906|317|1
35.024464|fda1ce737597e4b28558e3b4bd0e180a822be11c|3.89|2015-02-27 16:01:00|1.41290891556208|1|7184005080|317|0.6112922155462233|0|33|580|-80.847383|136|35.024464|OTHER MERCH DRESSINGS|0.89|4|MARIES CREAMY RANCH DRESSING|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00071840042819|OTHER MERCHANDISE|PRODUCE|-80.847383|1.4110530249708906|317|1
35.024464|d8d3d833588c6d7c18b4cab15602aca7fac9d31b|2.79|2015-03-02 18:00:00|1.41290891556208|1|3450015179|317|0.6112922155462233|0|33|312|-80.847383|51|35.024464|BUTTER|0.0|3|LOL HONEY BUTTER|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00034500151122|BUTTER & MARGARINE|DAIRY|-80.847383|1.4110530249708906|317|1
35.024464|629648512f9ead1503dd986655e5d1fdfd131390|5.69|2015-01-30 19:41:00|1.41290891556208|1|3680036723|317|0.6112922155462233|0|33|4236|-80.847383|1200|35.024464|DEX ADULT/CHILDREN|1.7|17|TC DAYTIME PE ORIGINAL LIQ|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00036800367326|COUGH/COLD/SINUS|HBC|-80.847383|1.4110530249708906|317|1
35.024464|d11812fa394216fe5a1439210ba91b31543dd3bf|4.49|2015-01-11 13:30:00|1.41290891556208|1||317|0.6112922155462233|0|33|557|-80.847383|64|35.024464|SPECIALTY-TROPICAL FRUIT|0.0|4|"HORNED MELON ""KIWANO"""|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00204302000007|FRESH PRODUCE|PRODUCE|-80.847383|1.4110530249708906|317|1
35.024464|1126e12fec7dd73b96e7af95e76697e61935c7e1|4.58|2015-02-14 10:51:00|1.41290891556208|1|20039000000|317|0.6112922155462233|0|33|1801|-80.847383|400|35.024464|FFM TURKEY|0.0|6|HONEY SMOKED TURKEY BREAST|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00200397000007|FFM MEAT|DELI|-80.847383|1.4110530249708906|317|1
35.024464|3c6fa0ccfcabb218afd4de1080ca62fbe0279766|1.29|2014-09-28 12:17:00|1.41290891556208|1||317|0.6112922155462233|0|33|505|-80.847383|64|35.024464|FRESH SOFT FRUIT|0.0|4|NECTARINES,TREE RIPE, XL|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00204378000000|FRESH PRODUCE|PRODUCE|-80.847383|1.4110530249708906|317|1
35.024464|d23c0ee61a70ff0406693461ef23cd396e2e7988|3.99|2015-01-18 17:58:00|1.41290891556208|1|7835470843|317|0.6112922155462233|0|33|317|-80.847383|52|35.024464|CHUNK AND BAR CHEESE|1.49|3|CABOT SERIOUSLY SHARP YELLOW|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00078354717288|CHEESE|DAIRY|-80.847383|1.4110530249708906|317|1
35.024464|919446b9a8f07e4488a6e4b6840efe239c9b990f|5.99|2014-12-22 12:51:00|1.41290891556208|1|7756725423|317|0.6112922155462233|0|33|252|-80.847383|45|35.024464|PREMIUM ICE CREAM|3.0|5|BREYERS CHOCOLATE I/C|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00077567254207|ICE CREAM|FROZEN|-80.847383|1.4110530249708906|317|1
35.024464|0d0c8bc8cdba92c3ce9744298ec0f57f040d9395|4.19|2014-10-11 14:33:00|1.41290891556208|1|4812127620|317|0.6112922155462233|0|33|1037|-80.847383|164|35.024464|ENGLISH MUFFINS|2.1|7|THOMAS 100% WHEAT ENG MUFN PP|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00048121184070|BREAKFAST|COMMERCIAL BAKERY|-80.847383|1.4110530249708906|317|1
35.024464|e697f77b7fe34b572850bbcc05ceb76a72e16a57|4.19|2014-09-10 09:32:00|80.811922674510953|1|4812127620|317|35.032960594179002|0|12|1037|-80.8062|164|35.037115|ENGLISH MUFFINS|2.1|7|THOMAS 100% WHEAT ENG MUFN PP|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|35.037868710371079|00048121184070|BREAKFAST|COMMERCIAL BAKERY|-80.847383|80.847386296408544|27|1
35.024464|1ab3ff07eec9b23780ab8ede2ef1215f6efe5307|12.79|2015-02-09 19:32:00|1.41290891556208|1|3700050963|317|0.6112922155462233|0|33|1513|-80.847383|66|35.024464|NFS-LAUNDRY DETERGENT PODS|0.0|1|TIDE PODS SPRING MEADOW 35CT|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00037000509639|DETERGENTS|G1 GROCERY|-80.847383|1.4110530249708906|317|1
35.024464|feb1163b7df99593a60301da454ea7afcff85f5b|1.0|2014-11-18 17:01:00|80.811922674510953|1|4000000435|317|35.032960594179002|0|12|47|-80.8062|7|35.037115|REGISTER BARS|0.2|1|(FE)M&M PLAIN CANDY|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|35.037868710371079|00040000000310|CANDY|G1 GROCERY|-80.847383|80.847386296408544|27|1
35.024464|fc2cfc0af4b1a42966c0da645893db101a477889|4.49|2015-01-19 10:32:00|1.41290891556208|1|70897191772|317|0.6112922155462233|0|33|1703|-80.847383|387|35.024464|SEASONAL COOKIES|1.0|14|VALENTINE PINK FRSTD SGR COOK|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00708971917722|COOKIES|BAKERY|-80.847383|1.4110530249708906|317|1
35.024464|8383801f4084446c69f936a8ed5a7791a71de955|3.79|2014-12-28 14:35:00|1.41290891556208|1|2500005542|317|0.6112922155462233|0|33|335|-80.847383|56|35.024464|ORANGE JUICE-REGRIGERATED|0.0|3|SIMPLY ORANGE ORIGINAL|948557ea59187c597ed841719f1f7710396ed85b|0.5870941688564538|0.61055446569467375|00025000055423|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.847383|1.4110530249708906|317|1
35.318911|1ffeef76a12ec18f0752fba5c6b06951fd3a6d3e|0.77|2015-03-05 19:12:00|80.77969194620016|4|7530000115|167|35.340551139241278|0|20|145|-80.764523|22|35.341927|MILK-CANNED|0.0|1|SUNSHINE EVAPORATED MILK|957afd9ade1056c0c280750541ec25e2733f252b|1.495281435645218|35.345012799095393|00075300001156|PACKAGED MILKS & MODIFIERS|G1 GROCERY|-80.780702|80.780710296270954|220|1
35.318911|c6c55186647c6ae540e22f5e69b6deea060d0938|2.27|2014-11-26 23:17:00|1.4094857484078087|4|3400056002|167|0.616431285168843|0|26|52|-80.780702|7|35.318911|PKG NON CHOC|0.0|1|TWIZZLERS STRAWBERRY TWISTS|957afd9ade1056c0c280750541ec25e2733f252b|1.495281435645218|0.61471665291522548|00034000560028|CANDY|G1 GROCERY|-80.780702|1.4098892219723687|167|1
35.116638|43c18c70a922747d7a3d195c532d1805d0d18417|19.96|2014-09-10 22:04:00|80.856688219393845|4|4260845977|204|35.144216891694164|0|15|139|-80.992182|20|35.103409|REMAINING SHELF STABLE JUICES|0.0|1|LAKEWOOD ORG SMT HLTH BLK CHRY|961cbc9a8216c74093b3a76a63427a95fea49aa4|1.905635344615347|35.134355925261694|00042608470748|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.85753|80.857555130813353|88|4
35.116638|1db528d4ac9225ee43d7d90b23c2cc3c4a606f3b|9.98|2014-09-10 06:34:00|80.856688219393845|4|4260845977|204|35.144216891694164|0|15|139|-80.992182|20|35.103409|REMAINING SHELF STABLE JUICES|0.0|1|LAKEWOOD ORG SMT HLTH BLK CHRY|961cbc9a8216c74093b3a76a63427a95fea49aa4|1.905635344615347|35.134355925261694|00042608470748|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.85753|80.857555130813353|88|2
35.585842|da994f419f8b302d6045488fe0ca8cf4cc6330c8|3.69|2015-01-10 10:24:00|1.4102725052409182|3|61144334026|99|0.6210901099944839|0|1|214|-80.875654|33|35.585842|BROTH|0.0|1|KITCHEN BASICS STOCK SEAFOOD|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00611443340310|SOUP|G1 GROCERY|-80.875654|1.411546447003722|99|1
35.585842|eacc998230d6a29beca5b0b31e8ceb3c9f04d288|5.19|2015-02-19 18:05:00|80.891462859624312|3|63561700001|99|35.633817747328614|0|45|162|-80.860108|25|35.500972|PICKLES|0.0|1|WICKLES PICKLES SWEET CHIPS|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|35.636605227883024|00635617000015|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.875654|80.87570173971686|268|1
35.585842|8cc3d4c78dadf9c127abef6f6feb7f8093a39989|1.23|2015-01-13 18:35:00|1.4102725052409182|3||99|0.6210901099944839|0|1|501|-80.875654|64|35.585842|FRESH PEARS|0.0|4|BARTLETT PEARS|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00204409000009|FRESH PRODUCE|PRODUCE|-80.875654|1.411546447003722|99|1
35.585842|9af2ba0c0fe4bcc52444d3b05804017629d8d576|6.87|2014-10-10 21:41:00|80.891462859624312|3|20165700000|99|35.633817747328614|0|45|297|-80.860108|49|35.500972|GROUND BEEF|0.77|2|HT GROUND BEEF CHUCK 80% LEAN|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|35.636605227883024|00201657000003|BEEF|MEAT|-80.875654|80.87570173971686|268|1
35.585842|df3f1f0c4731409ff67f167dd58a1a60957f5fbc|3.29|2014-09-14 17:34:00|1.4102725052409182|3|7203695076|99|0.6210901099944839|0|1|1609|-80.875654|371|35.585842|TAKE & BAKE BREAD|0.0|14|TAKE & BAKE SMALL WHEAT FRENCH|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00072036950765|BREAD|BAKERY|-80.875654|1.411546447003722|99|1
35.585842|e81909726278fc838e08b20850b92b77ba47be8e|3.99|2014-09-16 18:05:00|1.4102725052409182|3|3338300084|99|0.6210901099944839|0|1|500|-80.875654|64|35.585842|FRESH APPLES|0.0|4|GOLD DEL APPLE 3LB BAG|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00072036880277|FRESH PRODUCE|PRODUCE|-80.875654|1.411546447003722|99|1
35.585842|19fecfca618a5ca5f5bb8dfcfe2e09d92d52d291|3.29|2015-01-04 15:33:00|1.4102725052409182|3|7203695076|99|0.6210901099944839|0|1|1609|-80.875654|371|35.585842|TAKE & BAKE BREAD|1.3|14|TAKE & BAKE SMALL WHEAT FRENCH|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00072036950765|BREAD|BAKERY|-80.875654|1.411546447003722|99|1
35.585842|ba16d10a02f553e11556d3111132cb7b54f1d511|3.99|2014-12-24 13:45:00|1.4102725052409182|3|3338324028|99|0.6210901099944839|0|1|504|-80.875654|64|35.585842|FRESH BERRIES|2.32|4|BLACKBERRIES 5.6 OZ|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00761635202602|FRESH PRODUCE|PRODUCE|-80.875654|1.411546447003722|99|1
35.585842|30482976055d2fd1a5ea492ccc4fe4fcc6fad576|2.29|2014-10-19 18:22:00|80.891462859624312|3|7203695739|99|35.633817715990887|0|45|1976|-80.861571|475|35.444615|COLD PIZZA OTHER|0.0|6|WHITE PIZZA DOUGH BALLS|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|35.636605227883024|00072036957399|PIZZA|DELI|-80.875654|80.875736633553203|340|1
35.585842|6085b3171f2f62419850f0d0cb62c99363aad390|2.29|2014-11-16 13:21:00|1.4102725052409182|3|7203695739|99|0.6210901099944839|0|1|1976|-80.875654|475|35.585842|COLD PIZZA OTHER|0.0|6|WHITE PIZZA DOUGH BALLS|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00072036957399|PIZZA|DELI|-80.875654|1.411546447003722|99|1
35.585842|ceb1e010f1cc6d50c9d5a494b735612010c09eec|2.29|2015-02-22 17:34:00|1.4102725052409182|3|7203695739|99|0.6210901099944839|0|1|1976|-80.875654|475|35.585842|COLD PIZZA OTHER|0.0|6|WHITE PIZZA DOUGH BALLS|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00072036957399|PIZZA|DELI|-80.875654|1.411546447003722|99|1
35.585842|96168a73d4b3238dda37ffc512a6d8707e9e1cb2|0.97|2015-02-03 18:57:00|1.4102725052409182|3|7203671102|99|0.6210901099944839|0|1|1025|-80.875654|162|35.585842|WHITE|0.0|7|HT OLD FASHIONED BREAD|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00072036711021|SLICED BREAD|COMMERCIAL BAKERY|-80.875654|1.411546447003722|99|1
35.585842|31463d02fb45dedd7580e48993e6efcdd7e005da|3.29|2014-12-15 19:33:00|1.4102725052409182|3|7203695358|99|0.6210901099944839|0|1|1609|-80.875654|371|35.585842|TAKE & BAKE BREAD|0.0|14|TAKE & BAKE SMALL FRENCH BRD|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00072036953582|BREAD|BAKERY|-80.875654|1.411546447003722|99|1
35.585842|cbfead5dcd2ec05adbd33b78ac9b753bb4f0b81e|3.29|2014-09-17 19:15:00|1.4102725052409182|3|7203695358|99|0.6210901099944839|0|1|1609|-80.875654|371|35.585842|TAKE & BAKE BREAD|0.0|14|TAKE & BAKE SMALL FRENCH BRD|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00072036953582|BREAD|BAKERY|-80.875654|1.411546447003722|99|1
35.585842|d973342c774f322c6778a37c85f4e9000bff8cd1|2.99|2015-02-07 21:58:00|1.4102725052409182|3|3338322235|99|0.6210901099944839|0|1|504|-80.875654|64|35.585842|FRESH BERRIES|0.0|4|BLUEBERRIES PINT|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00033383222011|FRESH PRODUCE|PRODUCE|-80.875654|1.411546447003722|99|1
35.585842|1ba011dca7ee5ede8e89448e27ea7c5053a94e9d|3.79|2015-02-15 18:15:00|1.4102725052409182|3|7127927119|99|0.6210901099944839|0|1|555|-80.875654|64|35.585842|PACKAGED SALADS|0.0|4|F.E. SPINACH & ARUGULA|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00071279271194|FRESH PRODUCE|PRODUCE|-80.875654|1.411546447003722|99|1
35.585842|a8fb569efe180fad99fc64f01f858b134a07c655|3.79|2014-12-03 16:21:00|1.4102725052409182|3|7127927119|99|0.6210901099944839|0|1|555|-80.875654|64|35.585842|PACKAGED SALADS|0.0|4|F.E. SPINACH & ARUGULA|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00071279271194|FRESH PRODUCE|PRODUCE|-80.875654|1.411546447003722|99|1
35.585842|7fb70f4472aee5372e418455841f5ead95334353|3.79|2015-03-01 17:04:00|1.4102725052409182|3|4470000063|99|0.6210901099944839|0|1|359|-80.875654|101|35.585842|MEAT WIENERS|0.0|19|OSCAR MAYER SELECTS TURKEY FRK|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00044700007440|WIENERS|CASE READY MEATS|-80.875654|1.411546447003722|99|1
35.585842|c286ad7c456791ed96c258a4d6813531633d8a06|2.19|2014-10-23 18:03:00|1.4102725052409182|3|4900005010|99|0.6210901099944839|0|1|54|-80.875654|8|35.585842|DIET|0.2|23|DT CLASSIC 2 LITER|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00049000050110|CARBONATED BEVERAGES|BEVERAGE|-80.875654|1.411546447003722|99|1
35.585842|2a1f44cbdb318b7780f7ab848b276bd00362595b|4.29|2015-02-24 19:16:00|1.4102725052409182|3|76351451420|99|0.6210901099944839|0|1|330|-80.875654|55|35.585842|EGGS|1.29|3|DAVIDSON'S GRADE A LARGE WHITE|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00763514514202|EGGS FRESH|DAIRY|-80.875654|1.411546447003722|99|1
35.585842|958be2118bce04226a7c042eef6ae9310441b8f9|4.29|2014-12-06 18:23:00|1.4102725052409182|3|76351451420|99|0.6210901099944839|0|1|330|-80.875654|55|35.585842|EGGS|0.0|3|DAVIDSON'S GRADE A LARGE WHITE|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00763514514202|EGGS FRESH|DAIRY|-80.875654|1.411546447003722|99|1
35.585842|911e6fac9c6457bca53f4b23245f6955c965f33d|2.99|2015-03-02 18:52:00|1.4102725052409182|3|81204900640|99|0.6210901099944839|0|1|504|-80.875654|64|35.585842|FRESH BERRIES|0.0|4|BLUEBERRIES 6 OZ|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00891700002124|FRESH PRODUCE|PRODUCE|-80.875654|1.411546447003722|99|1
35.585842|b65aefdb46d735e0c5300bdb30fad0e3a56b963a|9.99|2014-11-12 18:21:00|1.4102725052409182|3|8500001660|99|0.6210901099944839|0|1|9962|-80.875654|887|35.585842|NFS-PREM-SAUV/FUME'BLANC|0.0|13|CB-STARBOROUGH SAUV BLANC|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00085000016602|SUPER PREMIUM ($11-$14.99)|WINE|-80.875654|1.411546447003722|99|1
35.585842|02c561cf91a91e1bd2f529aa0b8f0d2c49fb367e|5.99|2014-12-22 20:49:00|80.891462859624312|3|7778200787|99|35.633817715990887|0|45|355|-80.861571|104|35.444615|FRESH GRILLING SAUSAGE|0.0|19|JOHNSONVILLE HOT ITALIAN|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|35.636605227883024|00077782008135|DINNER SAUSAGE|CASE READY MEATS|-80.875654|80.875736633553203|340|1
35.585842|60cf11cf52279e3a30c0310548f91c4855bbfd92|8.99|2015-01-19 18:55:00|1.4102725052409182|3|2370002188|99|0.6210901099944839|0|1|291|-80.875654|48|35.585842|FROZEN POUTLRY|0.0|5|TYSON SOUTHWST CHK BRST STRIPS|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00023700016263|FROZEN MEALS|FROZEN|-80.875654|1.411546447003722|99|1
35.585842|2c582f6df955ebb8d4cc3da2bdccb86f5a27c86e|1.29|2014-09-26 14:25:00|1.4102725052409182|3||99|0.6210901099944839|0|1|527|-80.875654|64|35.585842|FRESH CARROTS|0.0|4|COO CARROTS, BUNCHED|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00204094000001|FRESH PRODUCE|PRODUCE|-80.875654|1.411546447003722|99|1
35.585842|a5fce4df94f610d2ffdb9fd4bde0f59374b49ea7|3.99|2015-01-23 18:36:00|1.4102725052409182|3|7203676057|99|0.6210901099944839|0|1|1220|-80.875654|275|35.585842|PASTA SC PREMIUM|1.49|1|HT TRADER SAUCE PUTTENESCA|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00072036760593|PASTA SAUCES|G1 GROCERY|-80.875654|1.411546447003722|99|1
35.585842|f46aa17f1c21e4e3dbc2d829a6a768a4f6dd4f14|3.79|2014-10-08 18:50:00|1.4102725052409182|3|8411410812|99|0.6210901099944839|0|1|201|-80.875654|31|35.585842|POTATO CHIPS|0.0|1|KETTLE BUFF  KRINKLE CUT CHIPS|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00084114113368|SNACKS|G1 GROCERY|-80.875654|1.411546447003722|99|1
35.585842|81b4fb5c19737d07f2c61def73332e5238b69c75|3.99|2014-12-23 17:25:00|1.4102725052409182|3|7203688128|99|0.6210901099944839|0|1|523|-80.875654|64|35.585842|FRESH POTATOES|0.0|4|HT RED CREAMER 24OZ BAG|9b6fde5665f4963dda6ada9411757d911fc95112|3.315009367933584|0.61833652052202714|00072036881281|FRESH PRODUCE|PRODUCE|-80.875654|1.411546447003722|99|1
35.000049|a207628b768f7ca75d7c70111bf5dee330ac1422|5.74|2014-09-13 17:53:00|1.4091206135396188|1|8130831863|249|0.6108660934093487|0|47|9935|-80.699686|885|35.000049|NFS POP CAB SAUV|0.0|13|OAK CREEK CABERNET|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00081308318639|POPULAR (4-$7.99)|WINE|-80.699686|1.4084752260255726|249|2
35.000049|1dad65443ec1b5529d8ace10f9f70a98d5eed941|2.87|2015-02-07 14:19:00|80.699698036522989|1|8130831863|249|35.019719901926806|0|18|9935|-80.758228|885|34.95459|NFS POP CAB SAUV|0.0|13|OAK CREEK CABERNET|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|35.030887098939942|00081308318639|POPULAR (4-$7.99)|WINE|-80.699686|80.699703741785839|182|1
35.000049|5c9e4434d498e741b1a81c4cae5ef69c45b8f8ae|8.61|2015-01-09 12:33:00|1.4091206135396188|1|8130831863|249|0.6108660934093487|0|47|9935|-80.699686|885|35.000049|NFS POP CAB SAUV|0.0|13|OAK CREEK CABERNET|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00081308318639|POPULAR (4-$7.99)|WINE|-80.699686|1.4084752260255726|249|3
35.000049|15cd038d3714cf31c8849a45e4749cc26d757721|8.61|2015-01-25 16:31:00|1.4091206135396188|1|8130831863|249|0.6108660934093487|0|47|9935|-80.699686|885|35.000049|NFS POP CAB SAUV|0.0|13|OAK CREEK CABERNET|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00081308318639|POPULAR (4-$7.99)|WINE|-80.699686|1.4084752260255726|249|3
35.000049|4ce6557237a2a67acb815b67ef5f712e064fcc98|2.87|2014-12-12 16:50:00|80.699698036522989|1|8130831863|249|35.019719901926806|0|18|9935|-80.758228|885|34.95459|NFS POP CAB SAUV|0.0|13|OAK CREEK CABERNET|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|35.030887098939942|00081308318639|POPULAR (4-$7.99)|WINE|-80.699686|80.699703741785839|182|1
35.000049|b727d8b51fee6bd9d79164d9f53499f32bb55a5f|2.87|2014-10-04 12:43:00|1.4091206135396188|1|8130831863|249|0.6108660934093487|0|47|9935|-80.699686|885|35.000049|NFS POP CAB SAUV|0.0|13|OAK CREEK CABERNET|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00081308318639|POPULAR (4-$7.99)|WINE|-80.699686|1.4084752260255726|249|1
35.000049|e5692eaee8c12120dd05d262c066f86876524729|8.61|2014-11-21 17:17:00|1.4091206135396188|1|8130831863|249|0.6108660934093487|0|47|9935|-80.699686|885|35.000049|NFS POP CAB SAUV|0.0|13|OAK CREEK CABERNET|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00081308318639|POPULAR (4-$7.99)|WINE|-80.699686|1.4084752260255726|249|3
35.000049|5b9011463cbc650fbce305edfac192289757ef11|5.74|2014-12-20 17:28:00|80.699698036522989|1|8130831863|249|35.019719901926806|0|18|9935|-80.758228|885|34.95459|NFS POP CAB SAUV|0.0|13|OAK CREEK CABERNET|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|35.030887098939942|00081308318639|POPULAR (4-$7.99)|WINE|-80.699686|80.699703741785839|182|2
35.000049|1871a8df85813b740a2d4ea2ed7c9b204dfce7a2|5.74|2015-02-20 10:58:00|80.699698036522989|1|8130831863|249|35.019719901926806|0|18|9935|-80.758228|885|34.95459|NFS POP CAB SAUV|0.0|13|OAK CREEK CABERNET|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|35.030887098939942|00081308318639|POPULAR (4-$7.99)|WINE|-80.699686|80.699703741785839|182|2
35.000049|1aa49a422e06a148e5f829ae6fb00b870b8963bd|3.59|2014-11-10 15:01:00|1.4091206135396188|1|7342000024|249|0.6108660934093487|0|47|322|-80.699686|53|35.000049|SOUR CREAM|0.59|3|DAISY SOUR CREAM|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00073420000240|CULTURES|DAIRY|-80.699686|1.4084752260255726|249|1
35.000049|acd403a1a86c95730fd131c321ddcfd6439e4a92|0.47|2014-11-14 11:26:00|1.4091206135396188|1|7248600220|249|0.6108660934093487|0|47|11|-80.699686|2|35.000049|MUFFIN MIXES|0.0|1|JIFFY CORN MUFFIN MIX|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00072486002205|BAKING MIXES|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|c92daaa47c0b8139d7ad8ff90631ab58a60ef412|3.59|2014-10-24 17:05:00|1.4091206135396188|1|7342000024|249|0.6108660934093487|0|47|322|-80.699686|53|35.000049|SOUR CREAM|0.0|3|DAISY SOUR CREAM|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00073420000240|CULTURES|DAIRY|-80.699686|1.4084752260255726|249|1
35.000049|d7569358cb8f28058571ea5267294edb1887b73c|1.99|2014-10-06 16:49:00|80.699698036522989|1|7203698370|249|35.019719901926806|0|18|205|-80.758228|31|34.95459|REMAINING SNACKS|0.49|1|HT SNACK MIX TRADITIONAL|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|35.030887098939942|00072036983701|SNACKS|G1 GROCERY|-80.699686|80.699703741785839|182|1
35.000049|26f82766a279adc62d5c4712513f76611e3b1ef5|1.99|2014-09-22 15:34:00|1.4091206135396188|1|7203698370|249|0.6108660934093487|0|47|205|-80.699686|31|35.000049|REMAINING SNACKS|0.49|1|HT SNACK MIX TRADITIONAL|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00072036983701|SNACKS|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|5dbc0892c39b9702875e836290475027c8a99989|3.69|2014-11-25 18:23:00|1.4091206135396188|1|1800028794|249|0.6108660934093487|0|47|1268|-80.699686|54|35.000049|BAGELS AND MUFFINS|1.19|3|PILLSBURY ALL READY PIE CRUST|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00018000287949|DOUGH PRODUCTS|DAIRY|-80.699686|1.4084752260255726|249|1
35.000049|3a6e1650ec34de6996afd4e187e1826cbbc46672|2.77|2014-12-14 16:26:00|1.4091206135396188|1|3338353030|249|0.6108660934093487|0|47|523|-80.699686|64|35.000049|FRESH POTATOES|0.0|4|RUSSET POTATO 8LB BAG|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00033383530307|FRESH PRODUCE|PRODUCE|-80.699686|1.4084752260255726|249|1
35.000049|1cc1caf5cd31dfeb8b72633c089b5f9243deb43e|6.58|2014-09-12 16:15:00|1.4091206135396188|1|7203670548|249|0.6108660934093487|0|47|318|-80.699686|52|35.000049|SHREDDED/GRATED CHEESE|0.0|3|HTT PARMESAN/ROMANO SHRED|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00072036705488|CHEESE|DAIRY|-80.699686|1.4084752260255726|249|2
35.000049|bb4cb72ce25ec158a570454785fcb2457b03ba9c|6.58|2015-01-31 16:11:00|80.699698036522989|1|7203670548|249|35.019719901926806|0|18|318|-80.758228|52|34.95459|SHREDDED/GRATED CHEESE|1.58|3|HTT PARMESAN/ROMANO SHRED|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|35.030887098939942|00072036705488|CHEESE|DAIRY|-80.699686|80.699703741785839|182|2
35.000049|b3b97cec91b3555ff702a3b02a913e5f59a259f3|3.29|2015-02-16 14:23:00|1.4091206135396188|1|7203670548|249|0.6108660934093487|0|47|318|-80.699686|52|35.000049|SHREDDED/GRATED CHEESE|0.0|3|HTT PARMESAN/ROMANO SHRED|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00072036705488|CHEESE|DAIRY|-80.699686|1.4084752260255726|249|1
35.000049|ece9a8d223937572e93faaa96bb8b5c237e2767a|3.29|2015-03-07 17:22:00|80.699698036522989|1|7203661037|249|35.019719901926806|0|18|840|-80.758228|102|34.95459|TUBS|0.29|19|HT SMOKED PASTRAMI|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|35.030887098939942|00072036610492|LUNCHMEATS|CASE READY MEATS|-80.699686|80.699703741785839|182|1
35.000049|b405dd9455f078f7a9b77687f14399326a14294d|3.39|2014-11-15 12:23:00|1.4091206135396188|1|7203661037|249|0.6108660934093487|0|47|840|-80.699686|102|35.000049|TUBS|0.0|19|HT SMOKED PASTRAMI|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00072036610492|LUNCHMEATS|CASE READY MEATS|-80.699686|1.4084752260255726|249|1
35.000049|9ec794376360c5562c838e3a51e3aa7494533e2b|5.29|2014-11-28 20:06:00|1.4091206135396188|1|5150024177|249|0.6108660934093487|0|47|125|-80.699686|19|35.000049|PEANUT BUTTER|1.3|1|JIF CREAMY PEANUT BUTTER|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00051500241776|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|7a64cc92ac5ff92a5a4998b6cf8bc6150ff68a1f|5.29|2014-12-24 13:53:00|80.699698036522989|1|5150024177|249|35.019719901926806|0|18|125|-80.758228|19|34.95459|PEANUT BUTTER|1.3|1|JIF CREAMY PEANUT BUTTER|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|35.030887098939942|00051500241776|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.699686|80.699703741785839|182|1
35.000049|31929e826d4f2d53e62828004e9331502b291244|3.69|2014-11-07 17:46:00|80.699698036522989|1|74840428793|249|35.019719907205243|0|18|138|-80.8062|38|35.037115|RICE MICROWAVE|0.0|1|SEEDS MW ORG INDIAN RICE BLND|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|35.030887098939942|00748404288128|RICE GRAINS AND BEANS|G1 GROCERY|-80.699686|80.6996882842856|27|1
35.000049|19ea2c653266afc0a20af31bac44c20e46736c27|5.03|2014-10-16 16:30:00|80.699698036522989|1||249|35.019719901926806|0|18|529|-80.758228|64|34.95459|FRESH ASPARAGUS|1.89|4|GREEN  ASPARAGUS|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|35.030887098939942|00204080000008|FRESH PRODUCE|PRODUCE|-80.699686|80.699703741785839|182|1
35.000049|2bbdf65e50f8fb36ae13e2562e0e1a0a6f5a73a5|2.8|2014-11-26 17:14:00|80.699698036522989|1||249|35.019719901926806|0|18|526|-80.758228|64|34.95459|FRESH MUSHROOMS|0.0|4|USA OYSTER MUSHROOM, BULK|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|35.030887098939942|00204649000005|FRESH PRODUCE|PRODUCE|-80.699686|80.699703741785839|182|1
35.000049|0f4c592409a4f988c63c16081b5e6f65f721a235|10.49|2014-09-27 19:39:00|80.699698036522989|1|20889500000|249|35.019719901926806|0|18|648|-80.758228|154|34.95459|FISH FLTS/STK FARM RAISD|0.96|12|FR TILAPIA FILLET|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|35.030887098939942|00208895000000|FISH FILLETS/STEAKS|SEAFOOD|-80.699686|80.699703741785839|182|1
35.000049|5077d95535c1615f06836dd12d450355e4db50c6|13.69|2014-11-29 13:49:00|1.4091206135396188|1|20889500000|249|0.6108660934093487|0|47|648|-80.699686|154|35.000049|FISH FLTS/STK FARM RAISD|0.0|12|FR TILAPIA FILLET|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00208895000000|FISH FILLETS/STEAKS|SEAFOOD|-80.699686|1.4084752260255726|249|1
35.000049|7ec383b33f6c9c28d13ad1f51e346df7c1d39596|2.58|2014-09-17 16:49:00|1.4091206135396188|1||249|0.6108660934093487|0|47|508|-80.699686|64|35.000049|FRESH GRAPEFRUIT|0.0|4|RED GRAPEFRUIT LRG|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00204282000004|FRESH PRODUCE|PRODUCE|-80.699686|1.4084752260255726|249|2
35.000049|60d06b17892fe1c4e347505afdde5a0ef9c735a5|2.58|2014-10-01 15:12:00|80.699698036522989|1||249|35.019719907205243|0|18|508|-80.8062|64|35.037115|FRESH GRAPEFRUIT|0.0|4|RED GRAPEFRUIT LRG|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|35.030887098939942|00204282000004|FRESH PRODUCE|PRODUCE|-80.699686|80.6996882842856|27|2
35.000049|812862a76210ac9fce2662adf574c7ca5d1ce4e5|2.5|2015-02-21 11:35:00|1.4091206135396188|1|7203624020|249|0.6108660934093487|0|47|149|-80.699686|23|35.000049|WHSE PASTA CORE|0.0|1|HT PASTA PENNE RIGATE|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00072036240200|PASTA|G1 GROCERY|-80.699686|1.4084752260255726|249|2
35.000049|12355a43f170b1f7c55fc097d42533b86ed2693e|29.99|2015-02-13 18:18:00|1.4091206135396188|1|7023666023|249|0.6108660934093487|0|47|751|-80.699686|87|35.000049|NFS-BOUQUETS|0.0|9|EXPRESSIONS OF LOVE BOUQUET|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00070236660231|FLORAL|FLORAL|-80.699686|1.4084752260255726|249|1
35.000049|d86b2e2be55bddfc5c8d288e59de19f807310b3b|3.49|2014-10-03 18:03:00|1.4091206135396188|1|7225100347|249|0.6108660934093487|0|47|240|-80.699686|38|35.000049|COUS/ALT GRAINS|0.99|1|NEAR EAST COUS PRLD BASIL HERB|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00072251003536|RICE GRAINS AND BEANS|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|c04b4c162d59d74bada4a4cc458bc4005a335592|3.49|2014-12-08 12:53:00|1.4091206135396188|1|7225100347|249|0.6108660934093487|0|47|240|-80.699686|38|35.000049|COUS/ALT GRAINS|0.5|1|NEAR EAST COUS PRLD BASIL HERB|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00072251003536|RICE GRAINS AND BEANS|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|66b654bb2eccc313a5bfaf1bfbbf427744d11f21|1.79|2014-09-19 13:26:00|1.4091206135396188|1|7203670626|249|0.6108660934093487|0|47|1213|-80.699686|272|35.000049|HISP DINNERS/SHELLS|0.0|1|HT TACO SHELLS 12CT YELLOW|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00072036706263|HISPANIC PREP. FOODS|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|ecd56b1417e9f02361a0e2fc69d05003a5b1be0c|5.74|2014-11-02 14:43:00|80.699698036522989|1|8130831763|249|35.019719901926806|0|18|9934|-80.758228|885|34.95459|NFS POP CHARDONNAY|0.0|13|CB-OAK CREEK CHARDONNAY|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|35.030887098939942|00081308317632|POPULAR (4-$7.99)|WINE|-80.699686|80.699703741785839|182|2
35.000049|d8d1921e4c1604d25629fe51b2c0cb2ff49744be|5.79|2014-10-20 13:15:00|1.4091206135396188|1|3700035751|249|0.6108660934093487|0|47|417|-80.699686|71|35.000049|NFS-FABRIC SOFTENERS|0.0|1|DOWNY LIQ FAB SOFT CLEAN BREEZ|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00037000357568|LAUNDRY SUPPLIES|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|3b1714ff5cba3caa78568805df5c21b4aeb494dd|6.99|2014-12-09 13:34:00|1.4091206135396188|1|8813044434|249|0.6108660934093487|0|47|99|-80.699686|32|35.000049|LIQUID TEA|1.0|1|NESTEA DIET LEMON .5L 12PK|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00088130444383|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|f4fd6e0de5a1930967e33dbd9724449f66c4a029|7.99|2015-02-18 12:22:00|1.4091206135396188|1|8813044434|249|0.6108660934093487|0|47|99|-80.699686|32|35.000049|LIQUID TEA|1.0|1|NESTEA DIET LEMON .5L 12PK|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00088130444383|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|4fa85305df0b2074c82f308bfb7d92119757656f|14.99|2014-12-07 14:35:00|1.4091206135396188|1|62901400609|249|0.6108660934093487|0|47|1703|-80.699686|387|35.000049|SEASONAL COOKIES|5.0|14|EZ BUILD GINGERBREAD HOUSE KIT|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00629014006091|COOKIES|BAKERY|-80.699686|1.4084752260255726|249|1
35.000049|1c132c15f2d64c4e52fc18c4929c83175fb7cdc4|5.0|2014-11-16 15:33:00|80.699698036522989|1|8500001581|249|35.019719901926806|0|18|9943|-80.758228|885|34.95459|NFS POP RIESLING|0.0|13|BAREFOOT RIESLING|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|35.030887098939942|00085000015810|POPULAR (4-$7.99)|WINE|-80.699686|80.699703741785839|182|1
35.000049|c840d91eee8eb575de003cce2d8ff2b045994ca7|2.53|2014-09-21 13:47:00|80.699698036522989|1||249|35.019719902136032|0|18|522|-80.64817|64|35.04711|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|35.030887098939942|00204664000004|FRESH PRODUCE|PRODUCE|-80.699686|80.699703392557453|129|1
35.000049|4f508c33bca3b6200e28441f435ccf5674335d7d|1.39|2015-01-31 18:04:00|80.699698036522989|1|2146632306|249|35.019719901926806|0|18|1730|-80.758228|392|34.95459|CANDLES|0.0|14|ASST GLITTER CANDLE|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|35.030887098939942|00021466323069|DECORATING|BAKERY|-80.699686|80.699703741785839|182|1
35.000049|b8e450ab62ec64d39ae99265421d481472502436|3.99|2014-09-10 11:39:00|1.4091206135396188|1|1862703000|249|0.6108660934093487|0|47|42|-80.699686|6|35.000049|GRANOLA/YOGURT BARS|1.0|1|KASHI BAR CRN PUMPKIN SPICE FX|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00018627030126|BREAKFAST FOODS|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|489c65dfd50378518eda93155ff3bcf23407538b|3.59|2015-02-20 12:12:00|1.4091206135396188|1|5250005009|249|0.6108660934093487|0|47|182|-80.699686|28|35.000049|MAYO|1.09|1|DUKES MAYO 18 SQZ|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00052500050092|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|0dc8172466c2e6d71a025c3eafd763d58799264e|12.19|2015-01-27 20:18:00|1.4091206135396188|1|1380023260|249|0.6108660934093487|0|47|1280|-80.699686|48|35.000049|MULTI SERVE MEALS|0.0|5|STOUFFER LASAGNA|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00013800232601|FROZEN MEALS|FROZEN|-80.699686|1.4084752260255726|249|1
35.000049|93fe0cfa7260ca65da2fa55dd594bb8238844d2a|5.49|2014-12-26 13:22:00|1.4091206135396188|1|7895150058|249|0.6108660934093487|0|47|533|-80.699686|64|35.000049|FRESH PEPPERS|0.0|4|STOPLIGHT PEPPER 3PK|9bd29fd87c4ecbdb1069d98b4050807ca8ddbd60|1.3592121904901102|0.61242566243833529|00078951500580|FRESH PRODUCE|PRODUCE|-80.699686|1.4084752260255726|249|1
35.323246|390983027d2e20105f9963df4c4103487f070f9e|1.89|2014-10-17 17:44:00|80.945255278477163|4|3800084496|166|35.373402977206297|0|13|201|-80.780702|31|35.318911|POTATO CHIPS|0.0|1|PRINGLES CHEDDAR CHEESE|9c230de0a62ca51c981b996f144d96fd366a007f|3.4657268524388103|35.37387923947206|00038000844980|SNACKS|G1 GROCERY|-80.945176|80.945219124913962|167|1
35.323246|acb64dcc4ed1d4c13e4ef8ff68673aea8d6463c2|3.49|2014-11-26 15:28:00|80.945255278477163|4|3800039118|166|35.373402977206297|0|13|81|-80.780702|9|35.318911|RTE CEREAL KIDS|0.0|1|KELLOGG FROOT LOOPS 12.2|9c230de0a62ca51c981b996f144d96fd366a007f|3.4657268524388103|35.37387923947206|00038000391187|CEREAL|G1 GROCERY|-80.945176|80.945219124913962|167|1
35.323246|b9d4e57262556437bccaee3db55fd6fc757de647|1.49|2014-12-23 15:53:00|80.945255278477163|4|1254668004|166|35.373402978292219|0|13|48|-80.737839|7|35.297134|REGISTER GUM|0.0|1|STRIDE SPEARMINT SINGLES|9c230de0a62ca51c981b996f144d96fd366a007f|3.4657268524388103|35.37387923947206|00012546680042|CANDY|G1 GROCERY|-80.945176|80.945217182742951|258|1
35.323246|a7f5d0dd31489503f5cf8d25d2dde4cde3d0b9d9|29.98|2015-01-20 17:19:00|80.945255278477163|4|75444108251|166|35.373402977206297|0|13|663|-80.780702|154|35.318911|FISH FILLETS/STEAKS PKGD|10.04|12|TILAPIA FILLETS|9c230de0a62ca51c981b996f144d96fd366a007f|3.4657268524388103|35.37387923947206|00754441082513|FISH FILLETS/STEAKS|SEAFOOD|-80.945176|80.945219124913962|167|2
35.323246|a7034bdcb1251fd6f2e8803e01f4ffe5f7aa2200|2.65|2015-01-09 14:28:00|80.945255278477163|4|8768400095|166|35.373402978292219|0|13|121|-80.737839|20|35.297134|ASEPTIC JUICES|0.65|1|CAPRI SUN GRAPE 10 PACK|9c230de0a62ca51c981b996f144d96fd366a007f|3.4657268524388103|35.37387923947206|00087684001035|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.945176|80.945217182742951|258|1
35.323246|afbfc352f56c6c6a6616cdc35e3dd032716e6a22|2.79|2014-12-22 16:22:00|80.945255278477163|4|2740010307|166|35.373402977206297|0|13|313|-80.780702|51|35.318911|MARGARINE|0.0|3|COUNTRY CROCK SPREAD BOWL|9c230de0a62ca51c981b996f144d96fd366a007f|3.4657268524388103|35.37387923947206|00027400103070|BUTTER & MARGARINE|DAIRY|-80.945176|80.945219124913962|167|1
35.323246|e1f061e5f35e5d98bd3dbefabede082d2bdc02e6|2.79|2015-01-27 17:25:00|80.945255278477163|4|2740010307|166|35.373402977206297|0|13|313|-80.780702|51|35.318911|MARGARINE|0.0|3|COUNTRY CROCK SPREAD BOWL|9c230de0a62ca51c981b996f144d96fd366a007f|3.4657268524388103|35.37387923947206|00027400103070|BUTTER & MARGARINE|DAIRY|-80.945176|80.945219124913962|167|1
35.323246|34ad586edbc9b9e578fd0b0702e0759ae8743db1|3.79|2014-11-03 17:05:00|80.945255278477163|4|2500005542|166|35.373402977206297|0|13|335|-80.780702|56|35.318911|ORANGE JUICE-REGRIGERATED|0.0|3|SIMPLY ORANGE WITH MANGO|9c230de0a62ca51c981b996f144d96fd366a007f|3.4657268524388103|35.37387923947206|00025000054372|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.945176|80.945219124913962|167|1
35.323246|87df1b0713546513282d14c850fba0ff95e9cfb8|7.58|2014-12-01 18:11:00|80.945255278477163|4|2500005542|166|35.373402977206297|0|13|335|-80.780702|56|35.318911|ORANGE JUICE-REGRIGERATED|1.58|3|SIMPLY ORANGE WITH MANGO|9c230de0a62ca51c981b996f144d96fd366a007f|3.4657268524388103|35.37387923947206|00025000054372|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.945176|80.945219124913962|167|2
35.323246|bcfb257e9c1f8b60b5a7768072825178b271e8e9|4.49|2015-02-25 17:09:00|80.945255278477163|4|7203636053|166|35.373402978292219|0|13|31|-80.737839|4|35.297134|NON CARBONATED WATER|1.15|1|(U)HT SPRING WATER .5 LTR 24PK|9c230de0a62ca51c981b996f144d96fd366a007f|3.4657268524388103|35.37387923947206|00072036360533|BOTTLED WATER|G1 GROCERY|-80.945176|80.945217182742951|258|1
35.323246|efeaff93a8ea26f9a155cabb1fa21183f8d260f3|2.49|2015-01-02 13:41:00|80.945255278477163|4|60504939530|166|35.373402978292219|0|13|509|-80.737839|64|35.297134|FRESH CITRUS-REMAINING|0.0|4|LEMONS, SMALL 1LB BAG|9c230de0a62ca51c981b996f144d96fd366a007f|3.4657268524388103|35.37387923947206|00605049395300|FRESH PRODUCE|PRODUCE|-80.945176|80.945217182742951|258|1
35.323246|b79abcadee614a9441528ad6e1b730939aeb4bd4|1.69|2014-10-29 07:39:00|80.945255278477163|4|4900000044|166|35.373402977206297|0|13|55|-80.780702|8|35.318911|REGULAR|0.0|23|CB COKE SINGLE 20 OZ.|9c230de0a62ca51c981b996f144d96fd366a007f|3.4657268524388103|35.37387923947206|00049000000443|CARBONATED BEVERAGES|BEVERAGE|-80.945176|80.945219124913962|167|1
35.323246|adcb977422efad6a3bf96b771e02f85c36a880fc|0.99|2015-02-17 15:22:00|80.945255278477163|4||166|35.373402977206297|0|13|535|-80.780702|64|35.318911|FRESH GREENS|0.0|4|COO KALE, BULK|9c230de0a62ca51c981b996f144d96fd366a007f|3.4657268524388103|35.37387923947206|00204627000003|FRESH PRODUCE|PRODUCE|-80.945176|80.945219124913962|167|1
35.297134|d99497535c5102304f63a36c2dba6836b4c4da56|1.69|2015-01-03 17:11:00|80.737901233649083|1|4600082011|258|35.353744434231245|0|46|1212|-80.70901|272|35.17335|HISP BEANS/PEPPERS|0.0|1|OEP BEANS REFRIED FAT FREE|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|35.349871187060224|00046000820118|HISPANIC PREP. FOODS|G1 GROCERY|-80.737839|80.737919313662005|174|1
35.297134|a648740959460898b1a7279d2a7c40e40a79fb57|3.49|2015-01-18 17:45:00|1.4094857484078087|1|3800039118|258|0.6160512048176361|0|26|81|-80.737839|9|35.297134|RTE CEREAL KIDS|0.0|1|KELLOGG FROOT LOOPS 12.2|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00038000391187|CEREAL|G1 GROCERY|-80.737839|1.409141121495086|258|1
35.297134|9589cd79e7a514f6403a55b16545dc5d97bc9422|2.99|2014-10-27 20:12:00|1.4094857484078087|1|3620021922|258|0.6160512048176361|0|26|1219|-80.737839|275|35.297134|PASTA SC CORE|0.0|1|BERTOLLI SC CARBONA BACON|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00036200381052|PASTA SAUCES|G1 GROCERY|-80.737839|1.409141121495086|258|1
35.297134|0257d943ad843517f1f71146f8ff339bae90b4bd|2.99|2014-10-17 18:53:00|1.4094857484078087|1|81204900640|258|0.6160512048176361|0|26|504|-80.737839|64|35.297134|FRESH BERRIES|0.0|4|BLUEBERRIES 6 OZ|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00033383220222|FRESH PRODUCE|PRODUCE|-80.737839|1.409141121495086|258|1
35.297134|735710cb9f10f13cba565a0b568fb7e4f8d136d8|2.99|2014-11-22 16:42:00|1.4094857484078087|1|3620021922|258|0.6160512048176361|0|26|1219|-80.737839|275|35.297134|PASTA SC CORE|0.0|1|BERTOLLI SC CARBONA BACON|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00036200381052|PASTA SAUCES|G1 GROCERY|-80.737839|1.409141121495086|258|1
35.297134|f46d3537668dddc17c38a32b470b686409fe3b65|2.99|2015-02-15 18:54:00|1.4094857484078087|1||258|0.6160512048176361|0|26|504|-80.737839|64|35.297134|FRESH BERRIES|0.0|4|BLUEBERRIES PINT|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00033383222356|FRESH PRODUCE|PRODUCE|-80.737839|1.409141121495086|258|1
35.297134|fcb30fbedc48ca45771dca515c8e927f9fbbc0d5|3.99|2015-01-31 14:56:00|1.4094857484078087|1|7203671361|258|0.6160512048176361|0|26|317|-80.737839|52|35.297134|CHUNK AND BAR CHEESE|0.49|3|HT TRDR SHARP CHED CRACKER CUT|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00072036713612|CHEESE|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|67100b63b2ec19c72d4d184de28dc54658551bf7|3.38|2014-12-04 12:47:00|1.4094857484078087|1|7203688003|258|0.6160512048176361|0|26|527|-80.737839|64|35.297134|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00072036880031|FRESH PRODUCE|PRODUCE|-80.737839|1.409141121495086|258|2
35.297134|dad2367b2dc5f7715d2354d05b3e4ca3d5c6e25d|1.69|2015-02-22 16:45:00|80.737901233649083|1|7203688003|258|35.35374439709836|0|46|527|-80.739|64|35.141204|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|35.349871187060224|00072036880031|FRESH PRODUCE|PRODUCE|-80.737839|80.737951987301685|171|1
35.297134|b6e5be271d9e51f7c2ee32eec4105b7d368fa5eb|2.59|2014-11-03 18:41:00|1.4094857484078087|1|7203663996|258|0.6160512048176361|0|26|342|-80.737839|57|35.297134|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00072036631299|MILK|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|5ea923522e03fd0a8bf6480b2e7f6aaf315a4d11|2.69|2014-09-22 19:18:00|1.4094857484078087|1|7203663996|258|0.6160512048176361|0|26|342|-80.737839|57|35.297134|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00072036631299|MILK|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|4ad03a5f83a3c8e462e6162b73ca70cd5b86dc83|2.69|2014-10-20 17:46:00|1.4094857484078087|1|7203663996|258|0.6160512048176361|0|26|342|-80.737839|57|35.297134|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00072036631299|MILK|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|240d6026ff9cbb5a5b0d38da6875f7c581564c8e|2.59|2014-11-23 15:37:00|1.4094857484078087|1|7203663996|258|0.6160512048176361|0|26|342|-80.737839|57|35.297134|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00072036631299|MILK|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|93121e6d751bfbf58ed4d75fa70c786191c9d29d|2.29|2015-02-26 19:38:00|1.4094857484078087|1|7203663996|258|0.6160512048176361|0|26|342|-80.737839|57|35.297134|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00072036631299|MILK|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|01c4ee678aab79e0d464b0c587dd64faaf5ef68b|2.29|2015-01-23 16:35:00|1.4094857484078087|1|7203663996|258|0.6160512048176361|0|26|342|-80.737839|57|35.297134|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00072036631299|MILK|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|dc0c515d109f4734c44b249964e44ebfcedc411b|3.15|2015-03-04 15:58:00|1.4094857484078087|1|4060034500|258|0.6160512048176361|0|26|313|-80.737839|51|35.297134|MARGARINE|0.0|3|ICBINB SPREAD BOWL|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00040600345002|BUTTER & MARGARINE|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|55e9986a9c71431182949a055a7b443037b23627|3.15|2015-01-25 17:45:00|80.737901233649083|1|4060034500|258|35.353744434231245|0|46|313|-80.70901|51|35.17335|MARGARINE|0.0|3|ICBINB SPREAD BOWL|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|35.349871187060224|00040600345002|BUTTER & MARGARINE|DAIRY|-80.737839|80.737919313662005|174|1
35.297134|ac1fd139b9518676e27087c64d7eb6a12aec164d|2.0|2015-03-07 15:26:00|1.4094857484078087|1|4300000953|258|0.6160512048176361|0|26|272|-80.737839|307|35.297134|TOPPINGS FROZEN|0.0|5|COOL WHIP WHIPPED TOPPING|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00043000009536|DESSERTS FROZEN|FROZEN|-80.737839|1.409141121495086|258|1
35.297134|413e75099f4fc2bf15c5bcc3d880110040b92094|4.99|2014-12-14 18:37:00|1.4094857484078087|1|4082201114|258|0.6160512048176361|0|26|1878|-80.737839|435|35.297134|HUMMUS|4.99|6|SPINACH ARTICHOKE HUMMUS|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00040822027540|SALADS|DELI|-80.737839|1.409141121495086|258|1
35.297134|2296ceb8df9073f2d4fce99a6089b7e175016f68|3.29|2014-11-01 15:14:00|1.4094857484078087|1|5210000444|258|0.6160512048176361|0|26|1245|-80.737839|34|35.297134|SINGLE SPICES|0.0|1|E  MC CINNAMON SUGAR|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00052100004440|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.737839|1.409141121495086|258|1
35.297134|19c26fa484fbe2e44a1c8c27cbc183b85756a6e1|2.99|2014-10-12 13:51:00|80.737901233649083|1|7203688212|258|35.353744434231245|0|46|555|-80.70901|64|35.17335|PACKAGED SALADS|0.49|4|HT SPRING MIX|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|35.349871187060224|00072036882127|FRESH PRODUCE|PRODUCE|-80.737839|80.737919313662005|174|1
35.297134|7c202aa5e712f2566399937b8712abe512831fad|2.69|2014-11-12 17:54:00|1.4094857484078087|1|7225001739|258|0.6160512048176361|0|26|1025|-80.737839|162|35.297134|WHITE|0.0|7|NATOWN WHITEWHEAT RTOP BRD|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00072250017398|SLICED BREAD|COMMERCIAL BAKERY|-80.737839|1.409141121495086|258|1
35.297134|b05619d7d7173b452575a83899eb1c1cfc764e61|1.77|2014-12-08 18:03:00|1.4094857484078087|1|7203698067|258|0.6160512048176361|0|26|365|-80.737839|56|35.297134|REFRIGERATED TEAS|0.74|3|HARRIS TEETER SWEET TEA|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00072036980670|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|be38935b2fa344e561536bdb664725e0bae95c53|1.77|2014-09-14 15:25:00|1.4094857484078087|1|7203698067|258|0.6160512048176361|0|26|365|-80.737839|56|35.297134|REFRIGERATED TEAS|0.0|3|HARRIS TEETER SWEET TEA|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00072036980670|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|3bd4577b8054c7c4273339ce4724b1e5799aaa45|1.77|2014-12-07 18:22:00|1.4094857484078087|1|7203698067|258|0.6160512048176361|0|26|365|-80.737839|56|35.297134|REFRIGERATED TEAS|0.0|3|HARRIS TEETER SWEET TEA|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00072036980670|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|1a7dfb1ca35880a0072aa6d87be62e80a57a51ec|2.69|2014-12-27 19:48:00|1.4094857484078087|1|7225001739|258|0.6160512048176361|0|26|1025|-80.737839|162|35.297134|WHITE|0.5|7|NATOWN WHITEWHEAT RTOP BRD|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00072250017398|SLICED BREAD|COMMERCIAL BAKERY|-80.737839|1.409141121495086|258|1
35.297134|dbbd5d7f32c5cf1d6d9058d67f5b0cdeecea5af8|3.99|2014-12-24 12:41:00|1.4094857484078087|1|4157005982|258|0.6160512048176361|0|26|1148|-80.737839|21|35.297134|ALMONDS|0.5|1|BLUE DIAMOND WHOLE NAT ALMOND|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00041570003831|NUTS|G1 GROCERY|-80.737839|1.409141121495086|258|1
35.297134|00c2388d5ad9ba7e089485c80e942865b9f484f3|3.99|2014-09-28 15:46:00|80.737901233649083|1|4400002854|258|35.353744434231245|0|46|1248|-80.70901|12|35.17335|SANDWICH COOKIES|1.49|1|OREO GOLDEN|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|35.349871187060224|00044000032586|COOKIES|G1 GROCERY|-80.737839|80.737919313662005|174|1
35.297134|6c2f4ebee1e4782fd83030a851f67f04670d8aba|52.35000000000002|2014-09-10 09:31:00|1.4094857484078087|1|6484939120|258|0.6160512048176361|0|26|7194|-80.737839|1600|35.297134|SPRING/SUMMER TOYS|2.62|18|I/O POOL NOODLE|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00064849391200|SEASONAL MERCHANDISE|GM|-80.737839|1.409141121495086|258|15
35.297134|405167804b4d7509df23be3daee502a82b396504|2.49|2014-12-17 17:35:00|1.4094857484078087|1|5040073942|258|0.6160512048176361|0|26|1033|-80.737839|163|35.297134|HAMBURGER|0.0|7|BALL PARK WHITE HAMS 8PK PP|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00050400739420|BUNS/ROLLS|COMMERCIAL BAKERY|-80.737839|1.409141121495086|258|1
35.297134|16ab9b999f4c5cf24390c0e187e26bc99bee85d8|1.25|2015-03-08 22:18:00|1.4094857484078087|1|5100002421|258|0.6160512048176361|0|26|214|-80.737839|33|35.297134|BROTH|0.0|1|SWANSON BROTH CHICKEN|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00051000024312|SOUP|G1 GROCERY|-80.737839|1.409141121495086|258|1
35.297134|d75362631e24d2669ab28e9885ff7440cb0c2147|2.49|2015-01-02 17:15:00|1.4094857484078087|1|5040073942|258|0.6160512048176361|0|26|1033|-80.737839|163|35.297134|HAMBURGER|0.0|7|BALL PARK WHITE HAMS 8PK PP|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00050400739420|BUNS/ROLLS|COMMERCIAL BAKERY|-80.737839|1.409141121495086|258|1
35.297134|bde3f3bb3ff4ee1e38f16738787a92a911e9d926|5.99|2014-12-29 16:48:00|80.737901233649083|1|7756725423|258|35.353744434231245|0|46|252|-80.70901|45|35.17335|PREMIUM ICE CREAM|1.41|5|BREYERS H'MADE VANILLA I/C|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|35.349871187060224|00077567226006|ICE CREAM|FROZEN|-80.737839|80.737919313662005|174|1
35.297134|bcd85ad5be0e0527e81f8a49438bfa7e365ad2c8|3.49|2015-01-09 18:32:00|1.4094857484078087|1|7203663995|258|0.6160512048176361|0|26|342|-80.737839|57|35.297134|FRESH MILK|0.0|3|HARRIS TEETER 1/2% MILK GALL|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00072036632012|MILK|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|76462680b6d62a8e1dcadcaa903d15a57517e85e|5.99|2014-11-25 21:17:00|1.4094857484078087|1|7756725423|258|0.6160512048176361|0|26|252|-80.737839|45|35.297134|PREMIUM ICE CREAM|3.0|5|BREYERS EX CREAMY VANILLA|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00077567250049|ICE CREAM|FROZEN|-80.737839|1.409141121495086|258|1
35.297134|dc544f03a27c2cb030280ed1830c9632866a8460|4.78|2015-02-10 13:32:00|1.4094857484078087|1|7357013000|258|0.6160512048176361|0|26|1267|-80.737839|53|35.297134|DIPS AND SPREADS|0.0|3|HELUVA GOOD FRENCH ONION DIP|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00073570130002|CULTURES|DAIRY|-80.737839|1.409141121495086|258|2
35.297134|72ee9276dae9fee1780ee29083df2aed5162f96d|1.99|2014-10-14 16:45:00|1.4094857484078087|1|7203688083|258|0.6160512048176361|0|26|526|-80.737839|64|35.297134|FRESH MUSHROOMS|0.0|4|HT WHITE MUSHROOMS, 8 OZ WHOLE|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00072036880833|FRESH PRODUCE|PRODUCE|-80.737839|1.409141121495086|258|1
35.297134|e417a2f262b3b486481798d60b7fe3265190f203|1.99|2015-02-07 13:31:00|1.4094857484078087|1|7203688083|258|0.6160512048176361|0|26|526|-80.737839|64|35.297134|FRESH MUSHROOMS|0.0|4|HT WHITE MUSHROOMS, 8 OZ WHOLE|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00072036880833|FRESH PRODUCE|PRODUCE|-80.737839|1.409141121495086|258|1
35.297134|beb70bfa8da337d5b8cce92d3aec13568c67311a|0.99|2015-01-30 20:01:00|1.4094857484078087|1|7203698291|258|0.6160512048176361|0|26|245|-80.737839|39|35.297134|VEGETABLES-CORE|0.39|1|HT PEAS SWEET|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00072036410214|VEGETABLES-CAN/JAR|G1 GROCERY|-80.737839|1.409141121495086|258|1
35.297134|a2e20fdd1730cf381c6b1ebc6a6ec7a8f8613edd|2.49|2014-09-20 18:48:00|1.4094857484078087|1|7203603104|258|0.6160512048176361|0|26|757|-80.737839|3|35.297134|BAKING NUTS|0.0|1|HT PECAN CHIPS PEG|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00072036031044|BAKING SUPPLIES|G1 GROCERY|-80.737839|1.409141121495086|258|1
35.297134|8c5422237a390bc8a117fb4b0aa1e184cd2d3d7b|2.0|2014-11-17 14:41:00|1.4094857484078087|1|2500004748|258|0.6160512048176361|0|26|338|-80.737839|56|35.297134|OTHER FRUIT JUICES|0.0|3|MINUTE MAID LEMONADE|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00025000047480|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|127d2c1df8f70c9b4cb03a3e9f7b189efd007fe4|3.19|2014-12-19 20:45:00|1.4094857484078087|1|2100012281|258|0.6160512048176361|0|26|320|-80.737839|53|35.297134|COTTAGE CHEESE|0.0|3|BREAKSTONE LRG CURD 4% COTTGE|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00021000122813|CULTURES|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|c23566f3871c1dcdeb07d39b34846135e3e0a59c|4.29|2014-11-22 16:43:00|1.4094857484078087|1|2100004007|258|0.6160512048176361|0|26|332|-80.737839|52|35.297134|STRING/SNACK|0.0|3|CRACKER BARREL CHEESE STICK 2|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00021000040087|CHEESE|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|77c06bb2cedcbde9ab01ca9718d99a5ca62a0e43|3.99|2014-09-14 15:19:00|1.4094857484078087|1|7203695676|258|0.6160512048176361|0|26|1656|-80.737839|381|35.297134|CUP CAKES|0.0|14|FFM MINI VANILLA CUPCAKES|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00072036956767|CAKES|BAKERY|-80.737839|1.409141121495086|258|1
35.297134|e3f674cf1e160675b48d3f8905ea3c81985b3336|1.69|2014-10-05 18:02:00|80.737901233649083|1|4900000044|258|35.353744434231245|0|46|54|-80.70901|8|35.17335|DIET|0.0|23|CB C/F DIET COKE CONTOUR|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|35.349871187060224|00049000000467|CARBONATED BEVERAGES|BEVERAGE|-80.737839|80.737919313662005|174|1
35.297134|9a52fddc4946082f14543326d9c44d10c44fb97e|3.99|2015-02-11 13:30:00|1.4094857484078087|1|3338300084|258|0.6160512048176361|0|26|500|-80.737839|64|35.297134|FRESH APPLES|0.0|4|GOLD DEL APPLE 3LB BAG|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00072036880277|FRESH PRODUCE|PRODUCE|-80.737839|1.409141121495086|258|1
35.297134|4b6c3a60bc9c44e34371824321d7bd51cf194d7a|3.99|2015-01-20 17:47:00|1.4094857484078087|1|3338300084|258|0.6160512048176361|0|26|500|-80.737839|64|35.297134|FRESH APPLES|0.0|4|GOLD DEL APPLE 3LB BAG|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00072036880277|FRESH PRODUCE|PRODUCE|-80.737839|1.409141121495086|258|1
35.297134|49c9f49bf11a470bb3e7e029822e1f902029210f|4.99|2014-11-14 16:45:00|1.4094857484078087|1|7144830025|258|0.6160512048176361|0|26|2021|-80.737839|505|35.297134|FRESH CHEESE|1.49|6|ALOUETTE GARLIC & HERB|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00071448300144|SPECIALTY CHEESE|DELI|-80.737839|1.409141121495086|258|1
35.297134|fb28885daff57f25a8e6d020af46deee5fa26591|3.19|2014-09-27 09:02:00|1.4094857484078087|1|4400000055|258|0.6160512048176361|0|26|88|-80.737839|13|35.297134|FLAKED SODA CRACKERS|0.69|1|NABISCO PREMIUMS|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00044000000578|CRACKERS|G1 GROCERY|-80.737839|1.409141121495086|258|1
35.297134|7256c3a3a52f2de2b41cff2c875f5947f8752cb5|11.69|2014-10-04 19:27:00|1.4094857484078087|1|20858800000|258|0.6160512048176361|0|26|648|-80.737839|154|35.297134|FISH FLTS/STK FARM RAISD|0.0|12|FRESH BONELESS SALMON FILLET|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00208588000003|FISH FILLETS/STEAKS|SEAFOOD|-80.737839|1.409141121495086|258|1
35.297134|023ce78762b7b81bca05044c82fd0726f4a77ce1|3.29|2014-09-29 18:26:00|1.4094857484078087|1|3000005040|258|0.6160512048176361|0|26|12|-80.737839|2|35.297134|PANCAKE MIXES|0.0|1|AJEMIMA COMP B-MILK P-CAKE|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00030000053003|BAKING MIXES|G1 GROCERY|-80.737839|1.409141121495086|258|1
35.297134|f639f4d18e7603faef2f1d6d85108c1f3a73f218|2.58|2014-12-03 18:30:00|1.4094857484078087|1|4920005675|258|0.6160512048176361|0|26|226|-80.737839|35|35.297134|SUGAR-POWDERED|0.6|1|DOMINO 10X CONF.SUGAR-BOX|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00049200051009|SUGAR/SUBSTITUTES|G1 GROCERY|-80.737839|1.409141121495086|258|2
35.297134|ae736dade7d897be6a2022660072df3a5d92f932|2.69|2015-01-13 18:05:00|1.4094857484078087|1|7294570544|258|0.6160512048176361|0|26|1025|-80.737839|162|35.297134|WHITE|0.0|7|SL S&S  W.G. WHITE BREAD|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00072945705449|SLICED BREAD|COMMERCIAL BAKERY|-80.737839|1.409141121495086|258|1
35.297134|ab584cdba09f64d07896e595e50656c58d10e159|2.59|2015-01-17 23:44:00|1.4094857484078087|1|7203695298|258|0.6160512048176361|0|26|1654|-80.737839|381|35.297134|DESSERT CAKES|0.0|14|OLD FASHION FUDGE CAKE SLICE|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00072036952981|CAKES|BAKERY|-80.737839|1.409141121495086|258|1
35.297134|de8277efe499814511c432dbcc7a08b552115e61|5.25|2014-11-26 11:01:00|1.4094857484078087|1||258|0.6160512048176361|0|26|538|-80.737839|64|35.297134|FRESH BEANS|0.52|4|COO GREEN BEANS, BULK|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00204066000008|FRESH PRODUCE|PRODUCE|-80.737839|1.409141121495086|258|1
35.297134|0b9096f27540f0483b98e4d51fe3d164639048b4|1.52|2014-10-28 19:32:00|1.4094857484078087|1|20897500000|258|0.6160512048176361|0|26|977|-80.737839|201|35.297134|FRESH HT CHICKEN|0.76|2|FRESH BONELESS CHICKEN BREAST|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00208975000005|POULTRY|MEAT|-80.737839|1.409141121495086|258|1
35.297134|a1acb337705cb1c50e2af13bd60ea4b6f57042c9|6.58|2015-03-05 17:48:00|1.4094857484078087|1|20897500000|258|0.6160512048176361|0|26|977|-80.737839|201|35.297134|FRESH HT CHICKEN|3.3|2|FRESH BONELESS CHICKEN BREAST|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00208975000005|POULTRY|MEAT|-80.737839|1.409141121495086|258|1
35.297134|98903fcf017a41b359c511b263b1280e61dc4b18|16.95|2014-12-24 11:34:00|1.4094857484078087|1|76211103160|258|0.6160512048176361|0|26|1598|-80.737839|369|35.297134|NFS MERCHANDISE|6.78|22|INK WAVES TMBLR HLDY14|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00762111031600|NFS STARBUCKS|COFFEE SHOP|-80.737839|1.409141121495086|258|1
35.297134|02e597849248b4fe0eb8c49de133c1d0586b4629|7.7|2015-01-14 13:57:00|1.4094857484078087|1||258|0.6160512048176361|0|26|503|-80.737839|64|35.297134|FRESH GRAPES|0.0|4|BLACK GRAPES, SEEDLESS 12/16|9c89f9d197f70fef83c51c18c98c672df4a2764d|3.911646916480473|0.61471665291522548|00204056000001|FRESH PRODUCE|PRODUCE|-80.737839|1.409141121495086|258|1
34.977331|478ea36f5050a3207cacacf44d72782e61bcc459|2.4|2014-11-02 09:34:00|1.41290891556208|1||149|0.6104695895098807|0|33|542|-81.027334|64|34.977331|FRESH VEGETABLES REMAIN|0.0|4|COO TURNIP ROOTS, BULK|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00204811000000|FRESH PRODUCE|PRODUCE|-81.027334|1.4141937624131469|149|1
34.977331|8edd28a6165b98d1f00bfce486e1bc8c4c6e7019|1.65|2015-02-22 10:16:00|1.41290891556208|1||149|0.6104695895098807|0|33|542|-81.027334|64|34.977331|FRESH VEGETABLES REMAIN|0.0|4|COO TURNIP ROOTS, BULK|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00204811000000|FRESH PRODUCE|PRODUCE|-81.027334|1.4141937624131469|149|1
34.977331|7ba42e71d8109553a322dbecd84eaa94decad8db|12.99|2014-11-17 16:24:00|1.41290891556208|1|36382400820|149|0.6104695895098807|0|33|4216|-81.027334|1200|34.977331|DECONGEST REMEDY-ADULT|3.0|17|MUCINEX EXPCTORANT 600MG 00820|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00363824008202|COUGH/COLD/SINUS|HBC|-81.027334|1.4141937624131469|149|1
34.977331|ddec907ad22ead8e0a93ef069e3bf376b2a951f7|4.99|2015-01-11 09:42:00|1.41290891556208|1|61611202795|149|0.6104695895098807|0|33|581|-81.027334|136|34.977331|FRESH SALSA|0.0|4|WHOLLY GUACAMOL CLASSIC 16OZ|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00616112027950|OTHER MERCHANDISE|PRODUCE|-81.027334|1.4141937624131469|149|1
34.977331|226453bdc9195733f532b8cdccbb57834342f082|7.18|2014-12-05 11:41:00|1.41290891556208|1|7027200216|149|0.6104695895098807|0|33|1132|-81.027334|55|34.977331|EGGS SUBSTITUTES|2.18|3|EGGBEATER CARTON|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00070272002163|EGGS FRESH|DAIRY|-81.027334|1.4141937624131469|149|2
34.977331|3c9a299c0fb16801a77ecc518d7914dd50d91020|4.49|2014-10-06 19:38:00|1.41290891556208|1|5210000373|149|0.6104695895098807|0|33|1245|-81.027334|34|34.977331|SINGLE SPICES|0.0|1|MC GOURMET PARSLEY FLAKES|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00052100003733|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|1141a86568e212d4fc60937d28c0bed21b6283ef|3.19|2014-09-27 17:10:00|1.41290891556208|1|7027200216|149|0.6104695895098807|0|33|1132|-81.027334|55|34.977331|EGGS SUBSTITUTES|0.0|3|EGGBEATER CARTON|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00070272002163|EGGS FRESH|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|e7601c2007367608caa58518cb809da287d676a6|6.99|2014-12-21 10:04:00|1.41290891556208|1|5210000383|149|0.6104695895098807|0|33|1245|-81.027334|34|34.977331|SINGLE SPICES|1.0|1|MC GOURMET DILL WEED|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00052100003832|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|d4c32f16e841e7aa5a5c78207534f676b174adc5|3.59|2014-11-28 12:56:00|1.41290891556208|1|7027200216|149|0.6104695895098807|0|33|1132|-81.027334|55|34.977331|EGGS SUBSTITUTES|0.4|3|EGGBEATER CARTON|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00070272002163|EGGS FRESH|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|1c1650dc43bfa47f4b38848a02a783814e5f859a|3.98|2014-12-31 11:32:00|1.41290891556208|1|7044640000|149|0.6104695895098807|0|33|498|-81.027334|111|34.977331|PICKLES & SAUERKRAUT|0.49|19|BOARS HEAD SAUERKRAUT 16 OZ|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00070446400009|MISC. PACKAGED MEATS|CASE READY MEATS|-81.027334|1.4141937624131469|149|2
34.977331|c2978cd4589f4c619d1ef4c092ec6ecc3b006197|3.25|2015-03-06 11:04:00|1.41290891556208|1|7203656080|149|0.6104695895098807|0|33|318|-81.027334|52|34.977331|SHREDDED/GRATED CHEESE|0.0|3|HT FANCY SHRED SWISS CHEESE|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00072036000200|CHEESE|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|581d190fc6ef10ed55010e1e3ceb411bf44080c1|4.0|2014-10-10 16:36:00|1.41290891556208|1||149|0.6104695895098807|0|33|511|-81.027334|64|34.977331|FRESH AVOCADOS|0.5|4|AVOCADOS, HASS XL 36CT|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00204770000004|FRESH PRODUCE|PRODUCE|-81.027334|1.4141937624131469|149|2
34.977331|b742316eb719cc3c187c74dfd7ebab35ca0a18c4|10.0|2015-02-08 10:13:00|1.41290891556208|1|61611227958|149|0.6104695895098807|0|33|581|-81.027334|136|34.977331|FRESH SALSA|0.0|4|WHOLLY GUACAMOLE CLASSIC 8OZ|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00616112279588|OTHER MERCHANDISE|PRODUCE|-81.027334|1.4141937624131469|149|4
34.977331|5b959f4161a00570d23ac507ab89276622077e18|13.98|2015-01-04 10:49:00|1.41290891556208|1|3700013885|149|0.6104695895098807|0|33|389|-81.027334|66|34.977331|NFS-LAUNDRY DETERGENTS|1.0|1|TIDE ULTRA STAIN RELEASE 46OZ|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00037000875864|DETERGENTS|G1 GROCERY|-81.027334|1.4141937624131469|149|2
34.977331|2712ebae743dfb9b05ef7dcf7a2d98e17d2d2b56|4.99|2015-01-18 09:57:00|1.41290891556208|1|4260845977|149|0.6104695895098807|0|33|139|-81.027334|20|34.977331|REMAINING SHELF STABLE JUICES|0.5|1|LAKEWOOD ORG SMT HLTH TRT CHRY|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00042608459774|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|d3a018188bb52fc8643e9f3f2bf526977865616b|4.79|2014-09-14 10:33:00|1.41290891556208|1|4720015264|149|0.6104695895098807|0|33|312|-81.027334|51|34.977331|BUTTER|2.02|3|CHALLENGE SALTED BUTTER|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00047200152641|BUTTER & MARGARINE|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|6230c4ade494fddef39e8c593f6841d3b85f11c5|4.99|2015-02-01 09:59:00|1.41290891556208|1|4260845977|149|0.6104695895098807|0|33|139|-81.027334|20|34.977331|REMAINING SHELF STABLE JUICES|0.5|1|LAKEWOOD ORG SMT HLTH TRT CHRY|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00042608459774|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|809881e9e4438901e09ba758f2c45d841e9c7931|4.99|2015-02-27 11:26:00|1.41290891556208|1|4260845977|149|0.6104695895098807|0|33|139|-81.027334|20|34.977331|REMAINING SHELF STABLE JUICES|0.0|1|LAKEWOOD ORG SMT HLTH TRT CHRY|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00042608459774|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|1f4e1167af7b836ffcd93f0f689f97d767c15e9a|4.0|2014-11-20 11:33:00|1.41290891556208|1|4300000953|149|0.6104695895098807|0|33|272|-81.027334|307|34.977331|TOPPINGS FROZEN|2.02|5|COOL WHIP WHIPPED TOPPING|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00043000009536|DESSERTS FROZEN|FROZEN|-81.027334|1.4141937624131469|149|2
34.977331|6146e3db01abc98e83ddfedf4f221940dcb613c2|3.49|2014-09-16 17:10:00|1.41290891556208|1|4400004557|149|0.6104695895098807|0|33|89|-81.027334|12|34.977331|GRAHAM CRACKERS|0.99|1|TEDDY GRAHAMS CHOCOLATE CHIP|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00044000005979|COOKIES|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|e24beae910fa9d3867f49095cb5bfc345ac8db2e|2.89|2014-09-16 08:41:00|1.41290891556208|1|4400000055|149|0.6104695895098807|0|33|88|-81.027334|13|34.977331|FLAKED SODA CRACKERS|0.0|1|NABISCO PREMIUMS|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00044000000578|CRACKERS|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|9a3ac49f7615587974a568f3f8e96f6234565c53|11.27|2014-12-18 11:56:00|1.41290891556208|1|20140400000|149|0.6104695895098807|0|33|296|-81.027334|49|34.977331|RANCHER BEEF|4.7|2|BEEF LOIN NY STRIP STEAK BNLS|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00201404000003|BEEF|MEAT|-81.027334|1.4141937624131469|149|1
34.977331|bb4ec6715c403b01d8e8a25d10a8547708119be5|2.19|2014-10-19 09:28:00|1.41290891556208|1|2400016717|149|0.6104695895098807|0|33|110|-81.027334|16|34.977331|FRUIT-CORE|0.52|1|DEL MONTE PEACH CHUNKS HS|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00024000058168|FRUIT-CAN/JAR|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|f9669a212dd2210cf1f1aa4327a26a3674d18769|0.97|2015-01-18 10:07:00|1.41290891556208|1|7203671102|149|0.6104695895098807|0|33|1025|-81.027334|162|34.977331|WHITE|0.0|7|HT OLD FASHIONED BREAD|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00072036711021|SLICED BREAD|COMMERCIAL BAKERY|-81.027334|1.4141937624131469|149|1
34.977331|c6094cece84422839a24e897ab30d4775e6aa0d8|0.97|2014-10-26 13:00:00|1.41290891556208|1|7203671102|149|0.6104695895098807|0|33|1025|-81.027334|162|34.977331|WHITE|0.0|7|HT OLD FASHIONED BREAD|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00072036711021|SLICED BREAD|COMMERCIAL BAKERY|-81.027334|1.4141937624131469|149|1
34.977331|873ed6885fd303296557137e05ea13c42fd353ee|5.99|2014-11-13 09:46:00|1.41290891556208|1|7778200787|149|0.6104695895098807|0|33|355|-81.027334|104|34.977331|FRESH GRILLING SAUSAGE|0.0|19|JOHNSONVILLE HOT ITALIAN|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00077782008135|DINNER SAUSAGE|CASE READY MEATS|-81.027334|1.4141937624131469|149|1
34.977331|bdd2c5b67726d785a796d24e1fa4518023661b88|3.89|2014-09-28 08:39:00|1.41290891556208|1|7835470749|149|0.6104695895098807|0|33|318|-81.027334|52|34.977331|SHREDDED/GRATED CHEESE|1.89|3|CABOT SHARP WHT CHEDDAR SHREDS|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00078354710968|CHEESE|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|e7ddfcb13ce8187a2c08c40d0fc32b865f35d8d3|4.99|2014-09-30 14:19:00|1.41290891556208|1|2858580102|149|0.6104695895098807|0|33|663|-81.027334|154|34.977331|FISH FILLETS/STEAKS PKGD|0.0|12|STEAMER LEMON DILL SALMON|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00028585801027|FISH FILLETS/STEAKS|SEAFOOD|-81.027334|1.4141937624131469|149|1
34.977331|64c183d3055381ef37b936de4a5348a7b6bd6b27|2.99|2014-09-11 11:05:00|1.41290891556208|1|2066200002|149|0.6104695895098807|0|33|184|-81.027334|28|34.977331|SALAD DRESSINGS-LIQUID|0.0|1|NEWMANS DRS VIN PARM RST GARL|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00020662002082|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|e132f95edcaa6efce4565e434db6c1eb3b6d3ed5|7.49|2014-10-27 11:32:00|1.41290891556208|1|6456322572|149|0.6104695895098807|0|33|291|-81.027334|48|34.977331|FROZEN POUTLRY|1.5|5|YUMMY-DINO BUDDIES|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00064563226345|FROZEN MEALS|FROZEN|-81.027334|1.4141937624131469|149|1
34.977331|90cc9f8b5b0d8ce7f280e2c209bb3e02bb933ae1|3.29|2014-10-02 16:59:00|1.41290891556208|1|2016922233|149|0.6104695895098807|0|33|469|-81.027334|198|34.977331|POTATOES|1.65|3|SIMPLY O'BRIEN HASH BROWNS|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00020169222129|POTATOES|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|dcd5d828903d9b2bd53c9a251c0af47f903b261e|2.11|2014-11-21 11:34:00|1.41290891556208|1||149|0.6104695895098807|0|33|500|-81.027334|64|34.977331|FRESH APPLES|0.0|4|GOLD DEL APPLE, WA 72|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00204020000006|FRESH PRODUCE|PRODUCE|-81.027334|1.4141937624131469|149|1
34.977331|a52c54d28c4073b6d2fb3fb0a6b37e0cd7802300|3.99|2014-10-12 16:13:00|1.41290891556208|1|88491218062|149|0.6104695895098807|0|33|61|-81.027334|9|34.977331|RTE CEREAL ADULT|0.0|1|POST SHREDDED WHEAT SPOON SIZE|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00884912180629|CEREAL|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|0e6fd2c3c5eaff2908f0be3e718edaf3b20680b6|4.69|2014-12-11 16:23:00|1.41290891556208|1|5100007620|149|0.6104695895098807|0|33|264|-81.027334|307|34.977331|DESSERT CAKES FROZEN|0.0|5|PEP FARM CHOCOLATE FUDGE CAKE|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00051000076236|DESSERTS FROZEN|FROZEN|-81.027334|1.4141937624131469|149|1
34.977331|f486af8b76653dbee893ffab75abedcf142c6452|12.99|2015-02-15 14:21:00|1.41290891556208|1|8308530096|149|0.6104695895098807|0|33|9961|-81.027334|887|34.977331|NFS-S/PREM-MERLOT|0.0|13|ESTANCIA MERLOT 750 ML|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00083085300968|SUPER PREMIUM ($11-$14.99)|WINE|-81.027334|1.4141937624131469|149|1
34.977331|2f718d459ad0c829b21993ba4b8fc0316df289ed|10.99|2014-11-17 16:26:00|1.41290891556208|1|8600381385|149|0.6104695895098807|0|33|9935|-81.027334|885|34.977331|NFS POP CAB SAUV|0.0|13|WOODBRIDGE CABERNET SAUV 1.5L|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00086003813854|POPULAR (4-$7.99)|WINE|-81.027334|1.4141937624131469|149|1
34.977331|4b747f02655497e88aa8d0048bc567209e9fad93|12.99|2014-11-01 14:28:00|1.41290891556208|1|8289610013|149|0.6104695895098807|0|33|9935|-81.027334|885|34.977331|NFS POP CAB SAUV|0.0|13|FETZER VALLEY OAKS CAB 1.5L|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00082896100132|POPULAR (4-$7.99)|WINE|-81.027334|1.4141937624131469|149|1
34.977331|165583f62cb67595cda3f3b556554b71285dfa62|4.19|2014-11-25 11:20:00|1.41290891556208|1|7101201050|149|0.6104695895098807|0|33|101|-81.027334|15|34.977331|FLOUR-ALL PURPOSE|1.2|1|KING ARTHUR UNBLEACH FLOUR-PLN|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00071012010509|FLOUR|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|5bdd4c656cb0664bb78a786d2f80cec493539221|1.77|2014-12-17 07:15:00|81.02739863253349|1|4178900121|149|35.015557116240501|0|14|1203|-80.810056|33|35.219587|RAMEN|0.77|1|MARUCHAN INSTANT LUNCH CHICKEN|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|35.014943729270243|00041789001215|SOUP|G1 GROCERY|-81.027334|81.027497361254916|401|3
34.977331|29cd68b5dc4264e4e35638fde07ba196c8ee128c|1.77|2014-12-22 07:37:00|81.02739863253349|1|4178900121|149|35.015557116240501|0|14|1203|-80.810056|33|35.219587|RAMEN|0.77|1|MARUCHAN INSTANT LUNCH CHICKEN|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|35.014943729270243|00041789001215|SOUP|G1 GROCERY|-81.027334|81.027497361254916|401|3
34.977331|b9d89aed21c99e2847d368a96fcc55d9a661f73a|11.97|2014-12-07 09:55:00|1.41290891556208|1|20405400000|149|0.6104695895098807|0|33|504|-81.027334|64|34.977331|FRESH BERRIES|6.97|4|RED RASPBERRIES 6 OZ|9e338a7539b48c9117f2464464ed23ad5abe7da3|2.6413485053299173|0.61055446569467375|00715756100019|FRESH PRODUCE|PRODUCE|-81.027334|1.4141937624131469|149|3
35.006282|2e657bfd021695afb5dd0a7f02c2e9a279bac625|4.9|2014-10-21 20:23:00|1.4091206135396188|4|7203663217|60|0.6109748797816256|0|47|330|-80.562829|55|35.006282|EGGS|0.9|3|HT GRADE A LARGE EGGS 18 CT|9f47f509e8dfb1332e922eab5ab1dfde7ee28587|18.78011652433307|0.61242566243833529|00072036632173|EGGS FRESH|DAIRY|-80.562829|1.4060866207711706|60|2
35.006282|22b419ffecaea7748aa93094e47f0d627e3209cc|9.38|2014-10-18 00:23:00|80.6036218474908|4|1111112425|60|35.278073049516308|0|34|726|-80.847383|73|35.024464|NFS-BODY WASHES|0.0|1|DOVE COOL MOISTURE BODY WASH|9f47f509e8dfb1332e922eab5ab1dfde7ee28587|18.78011652433307|35.262263711360632|00011111123311|PERSONAL SOAP/BATH ADDITIVES|G1 GROCERY|-80.562829|80.563194494659427|317|2
35.006282|3f4a6369a78ecabfde906674d418ff78e0c221fb|11.67|2014-10-15 15:24:00|80.6036218474908|4|3666906138|60|35.278073049516308|0|34|499|-80.847383|110|35.024464|MEATBALLS|4.26|19|COOKED PERFECT HOMESTYLE MTBLS|9f47f509e8dfb1332e922eab5ab1dfde7ee28587|18.78011652433307|35.262263711360632|00036669061380|FROZEN CASE MEAT|CASE READY MEATS|-80.562829|80.563194494659427|317|3
35.006282|5269aba41931977b84910a2c268b73a87a0c3e08|6.49|2014-10-16 23:15:00|80.6036218474908|4|31254770152|60|35.278073126202052|0|34|4030|-80.848528|1080|35.053394|ORAL RINSE-ANTISEPTIC|2.0|17|LISTERINE AMBER MOUTHWASH ORIG|9f47f509e8dfb1332e922eab5ab1dfde7ee28587|18.78011652433307|35.262263711360632|00312547701525|ORAL HYGIENE|HBC|-80.562829|80.563095920329417|11|1
35.006282|e801c0e4a28cad861716c6eedd061b144adcb590|2.65|2015-01-07 14:12:00|80.6036218474908|4|4119640471|60|35.278073063622358|0|34|1201|-80.850065|33|35.030252|RTS CANNED|2.65|1|PROG LIGHT CRM CHICKEN POT PIE|9f47f509e8dfb1332e922eab5ab1dfde7ee28587|18.78011652433307|35.262263711360632|00041196440829|SOUP|G1 GROCERY|-80.562829|80.563178455527193|470|1
35.006282|822acfb6e7db1e43fd842e9202572b0e621386c8|3.87|2014-10-20 21:13:00|80.6036218474908|4|3940001810|60|35.278073049516308|0|34|242|-80.847383|39|35.024464|CANNED BEANS|0.8699999999999999|1|BUSH PEAS BLACKEYE|9f47f509e8dfb1332e922eab5ab1dfde7ee28587|18.78011652433307|35.262263711360632|00039400013686|VEGETABLES-CAN/JAR|G1 GROCERY|-80.562829|80.563194494659427|317|3
35.006282|cd5fcc01cfa3a741bb7b5bf9f85e9d4a6f91b442|13.98|2015-01-13 21:54:00|80.6036218474908|4|4132231141|60|35.278073049516308|0|34|1277|-80.847383|279|35.024464|FROZEN SNACKS|3.98|5|FARM RICH MARINARA MOZ CH STX|9f47f509e8dfb1332e922eab5ab1dfde7ee28587|18.78011652433307|35.262263711360632|00041322356529|FROZEN SANDWICH AND SNACKS|FROZEN|-80.562829|80.563194494659427|317|2
34.95459|f2c52efc5a33c5a7d6aa3caca837047071900e20|2.5|2014-09-19 14:09:00|1.4091206135396188|4|7203695204|182|0.6100726841846847|0|47|1603|-80.758228|371|34.95459|PRIVATE LABEL BREAD|0.0|14|BAND OF BAKERS BAGUETTE|a10c6eadd1549b039e1a14eaa9fe9a045483ff62|2.6686016645045343|0.61242566243833529|00072036952042|BREAD|BAKERY|-80.758228|1.4094969766762753|182|1
34.95459|190edfad62190b38653c10a7ab1c791d5e54d93d|3.99|2014-09-21 18:22:00|1.4091206135396188|4|20980000000|182|0.6100726841846847|0|47|1677|-80.758228|383|34.95459|INDIVIDUALS (PASTRY CASE)|0.0|14|MASCARPONE CUP/GLASS|a10c6eadd1549b039e1a14eaa9fe9a045483ff62|2.6686016645045343|0.61242566243833529|00209811000005|PASTRY CASE|BAKERY|-80.758228|1.4094969766762753|182|1
34.95459|c97b53627599a928c151b60dc7c7db248b4196b8|7.99|2014-11-01 19:39:00|1.4091206135396188|4|8981950145|182|0.6100726841846847|0|47|9957|-80.758228|886|34.95459|NFS-PREM-OTHER RED|0.0|13|GABBIANO CHIANTI|a10c6eadd1549b039e1a14eaa9fe9a045483ff62|2.6686016645045343|0.61242566243833529|00089819501458|PREMIUM ($8-$10.99)|WINE|-80.758228|1.4094969766762753|182|1
34.95459|b60e873d36a9dc0d78e8213eda9cea9b2b498467|1.99|2014-10-23 14:34:00|1.4091206135396188|4||182|0.6100726841846847|0|47|561|-80.758228|64|34.95459|FR PROD ORGANIC PRODUCE|0.2|4|ORG PARSLEY, CURLY|a10c6eadd1549b039e1a14eaa9fe9a045483ff62|2.6686016645045343|0.61242566243833529|00294900000004|FRESH PRODUCE|PRODUCE|-80.758228|1.4094969766762753|182|1
34.95459|44951619d7e88b716de4fb39fc73fe179451efd3|4.29|2015-01-03 21:16:00|1.4091206135396188|4|2840006399|182|0.6100726841846847|0|47|204|-80.758228|31|34.95459|TORTILLA CHIPS|0.29|1|TOSTITOS MULTIGRAIN SCOOPS|a10c6eadd1549b039e1a14eaa9fe9a045483ff62|2.6686016645045343|0.61242566243833529|00028400036337|SNACKS|G1 GROCERY|-80.758228|1.4094969766762753|182|1
34.95459|dfd11ff8e993279ce7db37710bfdbe5635bca663|6.98|2014-12-10 20:37:00|80.758271881003409|4|7203695203|182|34.993210730168933|0|28|1639|-80.78468|377|35.096737|BULK (DONUTS)|0.0|14|6CT FRESH ASSORTED DONUTS|a10c6eadd1549b039e1a14eaa9fe9a045483ff62|2.6686016645045343|34.992988447249964|00072036952035|DONUTS|BAKERY|-80.758228|80.758292198850924|30|2
34.95459|f783d5f983a3dfa3ef747c14dc7bb379b048cef6|1.29|2014-12-08 13:19:00|80.758271881003409|4|1657191030|182|34.993210760331891|0|28|30|-80.837892|4|34.937113|CARBONATED WATER|0.29|1|SPARKLING ICE CRISP APPLE|a10c6eadd1549b039e1a14eaa9fe9a045483ff62|2.6686016645045343|34.992988447249964|00016571940379|BOTTLED WATER|G1 GROCERY|-80.758228|80.758253526040889|372|1
35.297134|e0ca69a36196a41d0c41f6a6b08ab19dff8ea235|7.98|2015-01-19 12:43:00|80.737901233649083|4|1630016564|258|35.347701015345997|0|46|335|-80.78468|56|35.096737|ORANGE JUICE-REGRIGERATED|2.98|3|FL NAT W/PULP ORANGE JUICE|a1675edaf5f9231a9815c7734d14d749f66809ed|3.4940678745850184|35.349871187060224|00016300165653|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.737839|80.7379814476554|30|2
35.297134|cf0074c4931cb6d95373646ca7a2c0ce95bda259|5.39|2014-10-13 18:25:00|80.737901233649083|4|4470000881|258|35.347701116367197|0|46|839|-80.810056|102|35.219587|STACK PACKS|0.0|19|OSCAR MAYER BEEF BOLOGNA|a1675edaf5f9231a9815c7734d14d749f66809ed|3.4940678745850184|35.349871187060224|00044700008812|LUNCHMEATS|CASE READY MEATS|-80.737839|80.737909315757989|401|1
35.667941|de0849e4207f426ce2d3f4829e4105e9718d81dc|8.89|2015-02-18 12:34:00|1.4057311447477159|2|20165700000|178|0.6225230078570788|0|52|297|-80.497332|49|35.667941|GROUND BEEF|0.99|2|HT GROUND BEEF CHUCK 80% LEAN|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00201657000003|BEEF|MEAT|-80.497332|1.4049434824709919|178|1
35.667941|1d5cebe7c331ea7699eb4c86779f1a8c19ad77f3|3.71|2014-10-27 13:22:00|1.4057311447477159|2||178|0.6225230078570788|0|52|501|-80.497332|64|35.667941|FRESH PEARS|0.0|4|BARTLETT PEARS|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00204409000009|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|4c7d5a77f373bffca13ebd3f2abd09946732f1f6|13.3|2015-01-07 13:43:00|1.4057311447477159|2|20254300000|178|0.6225230078570788|0|52|299|-80.497332|49|35.667941|ANGUS BEEF|4.49|2|VALUE PK ANGUS STEW MEAT|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00202543000008|BEEF|MEAT|-80.497332|1.4049434824709919|178|1
35.667941|78fd14e0c16864ad30cec1fcb6fce15a80dd251f|29.4|2015-01-06 19:03:00|1.4057311447477159|2|20165700000|178|0.6225230078570788|0|52|297|-80.497332|49|35.667941|GROUND BEEF|0.57|2|HT GROUND BEEF CHUCK 80% LEAN|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00201657000003|BEEF|MEAT|-80.497332|1.4049434824709919|178|6
35.667941|e26b53e50abc493a2d5682fd4d5b20bdf12ffa85|7.59|2015-03-08 14:35:00|80.497482303704658|2|20165700000|178|35.7478645851604|0|6|297|-80.780702|49|35.318911|GROUND BEEF|1.69|2|HT GROUND BEEF CHUCK 80% LEAN|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|35.699188602026126|00201657000003|BEEF|MEAT|-80.497332|80.497816662899567|167|1
35.667941|60e4358a304c117eee1edb0c1b982f5a15bd8b8f|2.55|2014-10-12 15:53:00|1.4057311447477159|2||178|0.6225230078570788|0|52|501|-80.497332|64|35.667941|FRESH PEARS|0.26|4|BARTLETT PEARS|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00204409000009|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|707ed2219046691d42cb477d8fd582e59cca98f5|54.199999999999996|2015-03-08 16:49:00|1.4057311447477159|2|20140400000|178|0.6225230078570788|0|52|296|-80.497332|49|35.667941|RANCHER BEEF|22.6|2|BEEF LOIN NY STRIP STEAK BNLS|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00201404000003|BEEF|MEAT|-80.497332|1.4049434824709919|178|4
35.667941|fdbc86e6948e889244c1d2f158e9abd5bfeefb9c|6.62|2015-02-16 13:26:00|1.4057311447477159|2|20598600000|178|0.6225230078570788|0|52|1800|-80.497332|400|35.667941|FFM BEEF|1.53|6|HT ROAST  BEEF|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00205986000000|FFM MEAT|DELI|-80.497332|1.4049434824709919|178|1
35.667941|3c381601564acf9387b6c2a682851dab3490bbfa|6.23|2014-12-03 14:23:00|1.4057311447477159|2|20598600000|178|0.6225230078570788|0|52|1800|-80.497332|400|35.667941|FFM BEEF|0.0|6|HT ROAST  BEEF|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00205986000000|FFM MEAT|DELI|-80.497332|1.4049434824709919|178|1
35.667941|23f3b856c9c060db7da3bbc20e2d55697e2a0982|8.15|2014-12-01 19:42:00|1.4057311447477159|2|20598600000|178|0.6225230078570788|0|52|1800|-80.497332|400|35.667941|FFM BEEF|0.0|6|HT ROAST  BEEF|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00205986000000|FFM MEAT|DELI|-80.497332|1.4049434824709919|178|1
35.667941|7d2953aacd6f28f86da6d08df4be45c0810f72e0|12.35|2014-11-10 19:56:00|1.4057311447477159|2|20598600000|178|0.6225230078570788|0|52|1800|-80.497332|400|35.667941|FFM BEEF|2.06|6|HT ROAST  BEEF|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00205986000000|FFM MEAT|DELI|-80.497332|1.4049434824709919|178|1
35.667941|ee82c0b8ed6c16460d620e19c98f0e7ca9bb6abe|6.62|2015-02-23 12:52:00|1.4057311447477159|2|20598600000|178|0.6225230078570788|0|52|1800|-80.497332|400|35.667941|FFM BEEF|0.0|6|HT ROAST  BEEF|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00205986000000|FFM MEAT|DELI|-80.497332|1.4049434824709919|178|1
35.667941|f4951b955dcf756e31923643ed1708e3d2485973|6.35|2014-12-08 13:29:00|1.4057311447477159|2|20598600000|178|0.6225230078570788|0|52|1800|-80.497332|400|35.667941|FFM BEEF|0.0|6|HT ROAST  BEEF|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00205986000000|FFM MEAT|DELI|-80.497332|1.4049434824709919|178|1
35.667941|d5d06df28417a94abfdc556bfc60212a15f9d64b|7.55|2014-10-21 12:06:00|1.4057311447477159|2|20598600000|178|0.6225230078570788|0|52|1800|-80.497332|400|35.667941|FFM BEEF|0.0|6|HT ROAST  BEEF|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00205986000000|FFM MEAT|DELI|-80.497332|1.4049434824709919|178|1
35.667941|1c643537b8164655976640a26f73b93c0907fdac|1.79|2015-02-25 18:31:00|80.497482303704658|2|7203688032|178|35.7478645851604|0|6|555|-80.780702|64|35.318911|PACKAGED SALADS|0.0|4|HT SHREDDED ICEBERG LETTUCE|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|35.699188602026126|00072036880321|FRESH PRODUCE|PRODUCE|-80.497332|80.497816662899567|167|1
35.667941|85e03f8255cf490d6d5d336b05469cc1c545a816|0.97|2014-09-11 16:03:00|1.4057311447477159|2|7203688002|178|0.6225230078570788|0|52|527|-80.497332|64|35.667941|FRESH CARROTS|0.0|4|HT WHOLE CARROTS 2LB BAG|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00072036880024|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|111a92cfbd75f2d910b639c793f329c993fee799|0.97|2014-11-07 16:51:00|1.4057311447477159|2|7203688002|178|0.6225230078570788|0|52|527|-80.497332|64|35.667941|FRESH CARROTS|0.0|4|HT WHOLE CARROTS 2LB BAG|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00072036880024|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|75e4875dfa7354140212b846f0b88316889fb70a|0.97|2015-02-12 10:30:00|1.4057311447477159|2|7203688002|178|0.6225230078570788|0|52|527|-80.497332|64|35.667941|FRESH CARROTS|0.0|4|HT WHOLE CARROTS 2LB BAG|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00072036880024|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|a7e59ebb9ca88ef1d9167313ee94d6ae31dabfb0|0.97|2015-03-05 15:15:00|1.4057311447477159|2|7203688002|178|0.6225230078570788|0|52|527|-80.497332|64|35.667941|FRESH CARROTS|0.0|4|HT WHOLE CARROTS 2LB BAG|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00072036880024|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|b0c9ab0d1dc9f95b38890215c70736f25b3b3aca|9.18|2014-11-01 10:57:00|1.4057311447477159|2|5450019322|178|0.6225230078570788|0|52|484|-80.497332|101|35.667941|BEEF WIENERS|2.29|19|BALL PARK BUN SIZE BEEF FRANK|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00054500193298|WIENERS|CASE READY MEATS|-80.497332|1.4049434824709919|178|2
35.667941|05ef520d31645aeaa682c2b4fa4f1b339be8867b|5.35|2015-01-26 19:31:00|1.4057311447477159|2|5450019322|178|0.6225230078570788|0|52|484|-80.497332|101|35.667941|BEEF WIENERS|2.68|19|BALL PARK BUN SIZE BEEF FRANK|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00054500193298|WIENERS|CASE READY MEATS|-80.497332|1.4049434824709919|178|1
35.667941|c242a6b2d6fa82d3a5884aef5a1299b972fb8b26|5.35|2015-01-31 16:01:00|1.4057311447477159|2|5450019322|178|0.6225230078570788|0|52|484|-80.497332|101|35.667941|BEEF WIENERS|2.68|19|BALL PARK BUN SIZE BEEF FRANK|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00054500193298|WIENERS|CASE READY MEATS|-80.497332|1.4049434824709919|178|1
35.667941|7f3e3acecbc0e61f3c119f028d2a7903ab677ab6|5.35|2015-01-26 19:30:00|1.4057311447477159|2|5450019322|178|0.6225230078570788|0|52|484|-80.497332|101|35.667941|BEEF WIENERS|2.68|19|BALL PARK BUN SIZE BEEF FRANK|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00054500193298|WIENERS|CASE READY MEATS|-80.497332|1.4049434824709919|178|1
35.667941|621c53ccb0a1978e6745cb0525e8b1f634af78e2|2.68|2014-09-30 13:46:00|1.4057311447477159|2|7203625010|178|0.6225230078570788|0|52|145|-80.497332|22|35.667941|MILK-CANNED|0.0|1|HT  EVAPORATED MILK|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00072036250100|PACKAGED MILKS & MODIFIERS|G1 GROCERY|-80.497332|1.4049434824709919|178|4
35.667941|deee64dcfbe5ef5e952cc4039434e0accb8d05bf|3.99|2015-02-10 17:33:00|80.497482303704658|2||178|35.7478645851604|0|6|529|-80.780702|64|35.318911|FRESH ASPARAGUS|1.0|4|GREEN  ASPARAGUS|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|35.699188602026126|00204080000008|FRESH PRODUCE|PRODUCE|-80.497332|80.497816662899567|167|1
35.667941|e70db9fa0952d2a8956cb973f12cd5c7664bcbaa|3.18|2014-11-26 13:15:00|1.4057311447477159|2|7800023046|178|0.6225230078570788|0|52|54|-80.497332|8|35.667941|DIET|0.59|23|CANADA DRY DT G/ALE 2 LITER|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00078000148466|CARBONATED BEVERAGES|BEVERAGE|-80.497332|1.4049434824709919|178|2
35.667941|ab585d68c884adfb8a4f216b7fd7a4e5c6046410|9.77|2014-10-28 16:20:00|1.4057311447477159|2|7203698308|178|0.6225230078570788|0|52|194|-80.497332|30|35.667941|OLIVE OIL|0.0|1|HT EXTRA VIRGIN OLIVE OIL|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00072036983084|SHORTENING/OIL|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|d5bfc6a027196ee4f481a472a749bf63fc58f5e3|2.29|2015-01-15 13:32:00|1.4057311447477159|2|7203663996|178|0.6225230078570788|0|52|342|-80.497332|57|35.667941|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00072036631299|MILK|DAIRY|-80.497332|1.4049434824709919|178|1
35.667941|e3b24666f0d335738746923e5357e498a4695383|2.29|2015-02-19 09:54:00|1.4057311447477159|2|7203663996|178|0.6225230078570788|0|52|342|-80.497332|57|35.667941|FRESH MILK|0.0|3|HARRIS TEETER WHOLE MILK|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00072036639967|MILK|DAIRY|-80.497332|1.4049434824709919|178|1
35.667941|fbb02ef01a96138af3cba76cc5bad889a748a98d|2.69|2014-10-09 17:00:00|1.4057311447477159|2|7203663996|178|0.6225230078570788|0|52|342|-80.497332|57|35.667941|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00072036631299|MILK|DAIRY|-80.497332|1.4049434824709919|178|1
35.667941|38ecb2ea52949fc745ee80b30b3ab062aee5f58f|2.29|2015-02-25 10:42:00|1.4057311447477159|2|7203663996|178|0.6225230078570788|0|52|342|-80.497332|57|35.667941|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00072036631299|MILK|DAIRY|-80.497332|1.4049434824709919|178|1
35.667941|6bb8d56d6bf8cc87d2d2e49e9f3ed165fad75c73|6.99|2014-11-24 13:51:00|1.4057311447477159|2|3770032228|178|0.6225230078570788|0|52|423|-80.497332|72|35.667941|NFS-DISPOSE PLATES/BOWLS|3.49|1|CHINET DINNER PLATE 10 3/8IN|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00037700322262|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|e13f87574fa1f94cca7201850c02ac982f1622b5|3.49|2014-11-21 15:52:00|1.4057311447477159|2|7096900009|178|0.6225230078570788|0|52|543|-80.497332|64|35.667941|FRESH GARLIC|0.0|4|MINCED GARLIC, JAR|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00070969000090|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|17fd3338f62840bd769987b2610c05162d7fd081|31.21|2015-01-09 18:16:00|1.4057311447477159|2|20234100000|178|0.6225230078570788|0|52|299|-80.497332|49|35.667941|ANGUS BEEF|10.42|2|ANGUS BEEF SIRLOIN TIP ROAST|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00202341000002|BEEF|MEAT|-80.497332|1.4049434824709919|178|2
35.667941|d23921df23efdd74d2a910ea3fc102089701ae59|10.29|2014-12-15 19:49:00|1.4057311447477159|2|20600100000|178|0.6225230078570788|0|52|1802|-80.497332|400|35.667941|FFM HAM|3.09|6|VIRGINIA BAKED HAM|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00206001000005|FFM MEAT|DELI|-80.497332|1.4049434824709919|178|1
35.667941|234cce53717a80e697d4f2431cad5f12a9bc77df|1.78|2014-10-15 15:21:00|1.4057311447477159|2|7203698210|178|0.6225230078570788|0|52|257|-80.497332|39|35.667941|TOMATOES|0.0|1|HT TOMATO SAUCE 15 NO SALT|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00072036982100|VEGETABLES-CAN/JAR|G1 GROCERY|-80.497332|1.4049434824709919|178|2
35.667941|a5a2e7334a6aac5822bdd360db5ddf1c353ff715|2.77|2014-12-31 09:14:00|1.4057311447477159|2|3338353030|178|0.6225230078570788|0|52|523|-80.497332|64|35.667941|FRESH POTATOES|0.0|4|RUSSET POTATO 8LB BAG|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00033383530307|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|3395221f3149f95acc1c68b84db5123160c1188c|5.99|2015-02-19 10:42:00|80.497482303704658|2|1834175105|178|35.7478645851604|0|6|9934|-80.780702|885|35.318911|NFS POP CHARDONNAY|0.0|13|CB-BAREFOOT CHARDONNAY|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|35.699188602026126|00018341751055|POPULAR (4-$7.99)|WINE|-80.497332|80.497816662899567|167|1
35.667941|c708586bd6344f1e409987b5665cc9a03cfab333|3.79|2015-02-20 18:12:00|80.497482303704658|2|7684010015|178|35.7478645851604|0|6|275|-80.780702|45|35.318911|SUPER PREMIUM ICE CREAM|0.0|5|BEN & JERRY RED VELVET CAKE|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|35.699188602026126|00076840128358|ICE CREAM|FROZEN|-80.497332|80.497816662899567|167|1
35.667941|8af8a7d1cab364f974fe8337f6fc8446c78d7dd2|8.99|2015-01-24 17:08:00|1.4057311447477159|2|7488201060|178|0.6225230078570788|0|52|1213|-80.497332|272|35.667941|HISP DINNERS/SHELLS|0.0|1|RIO RANCHO TOSTADO BOWLS|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00074882010600|HISPANIC PREP. FOODS|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|518e087aaebce59a7f327122e6e5d01daf791052|7.94|2014-09-20 18:35:00|1.4057311447477159|2|7203659020|178|0.6225230078570788|0|52|312|-80.497332|51|35.667941|BUTTER|0.0|3|HARRIS TEETER UNSALTED BUTTER|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00072036590213|BUTTER & MARGARINE|DAIRY|-80.497332|1.4049434824709919|178|2
35.667941|cceb78a7b7ce38523b193faedcaa090002be9f59|31.76|2014-12-13 09:42:00|1.4057311447477159|2|7203659020|178|0.6225230078570788|0|52|312|-80.497332|51|35.667941|BUTTER|11.76|3|HARRIS TEETER UNSALTED BUTTER|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00072036590213|BUTTER & MARGARINE|DAIRY|-80.497332|1.4049434824709919|178|8
35.667941|350ed392dc4c35bd8cbcb30f3e54c645ae3d85da|6.94|2015-02-01 18:39:00|1.4057311447477159|2|7203659020|178|0.6225230078570788|0|52|312|-80.497332|51|35.667941|BUTTER|1.5|3|HARRIS TEETER UNSALTED BUTTER|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00072036590213|BUTTER & MARGARINE|DAIRY|-80.497332|1.4049434824709919|178|2
35.667941|7b38ee5acc6a20abb052c24d42a67bf50f6a0a50|3.69|2015-02-13 17:24:00|80.497482303704658|2|7203688073|178|35.7478645851604|0|6|523|-80.780702|64|35.318911|FRESH POTATOES|0.0|4|HT BAKER POTATO 4 CT PKG|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|35.699188602026126|00072036880734|FRESH PRODUCE|PRODUCE|-80.497332|80.497816662899567|167|1
35.667941|fdaeb08bf62c9eb862c8664c78539f66582fa2ff|17.13|2015-02-14 15:12:00|1.4057311447477159|2|20302700000|178|0.6225230078570788|0|52|652|-80.497332|141|35.667941|FRESH LAMB PRIMALS|0.0|2|LAMB SEASONED BUTTERFLIED LEG|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00203027000002|LAMB|MEAT|-80.497332|1.4049434824709919|178|1
35.667941|034a4e5d63da456c381d9c1bc3c61155c6ae1c9d|9.98|2015-01-25 14:37:00|1.4057311447477159|2|8265750406|178|0.6225230078570788|0|52|31|-80.497332|4|35.667941|NON CARBONATED WATER|2.98|1|(U)DEER PARK WATER 24PK .5LT|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00082657504063|BOTTLED WATER|G1 GROCERY|-80.497332|1.4049434824709919|178|2
35.667941|9d86d04720ac2039a8da8d16a6a432e78dd22774|4.35|2014-10-13 19:33:00|1.4057311447477159|2|4400002747|178|0.6225230078570788|0|52|91|-80.497332|13|35.667941|SPRAYED BUTTER CRACKERS|1.35|1|RITZ CRACKERS|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00044000031114|CRACKERS|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|0d04f72e92553c57760ed5dec7d44a109c4c8514|2.49|2015-03-09 16:06:00|1.4057311447477159|2|5040073942|178|0.6225230078570788|0|52|1033|-80.497332|163|35.667941|HAMBURGER|0.0|7|BALL PARK WHITE HAMS 8PK PP|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00050400739420|BUNS/ROLLS|COMMERCIAL BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|20e1abf3cd96dcda274e6c322f51c4e74bb41163|2.49|2014-12-20 14:14:00|1.4057311447477159|2|5040073942|178|0.6225230078570788|0|52|1033|-80.497332|163|35.667941|HAMBURGER|0.0|7|BALL PARK WHITE HAMS 8PK PP|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00050400739420|BUNS/ROLLS|COMMERCIAL BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|ab414c4dcfbe3f3b66401c31255fba07ed73daa9|1.91|2015-01-16 12:00:00|1.4057311447477159|2||178|0.6225230078570788|0|52|522|-80.497332|64|35.667941|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00204664000004|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|df14376b7320c77a8f85c04c5d2d88af230bd873|2.79|2014-12-11 12:15:00|1.4057311447477159|2|5150020441|178|0.6225230078570788|0|52|103|-80.497332|15|35.667941|REMAINING FLOUR|0.3|1|PILLSBURY BEST FLOUR-UNBLEACHD|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00051500222416|FLOUR|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|f6f86a8493c98944a1710efd5d87edd4e1f6dabc|3.49|2014-10-31 12:53:00|1.4057311447477159|2|4812127620|178|0.6225230078570788|0|52|1037|-80.497332|164|35.667941|ENGLISH MUFFINS|1.75|7|THOMAS 100% WHEAT ENG MUFN PP|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00048121184070|BREAKFAST|COMMERCIAL BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|00259e0ca666d74f5060a9f470893a3feda8f474|3.58|2015-02-21 14:30:00|1.4057311447477159|2|5100005977|178|0.6225230078570788|0|52|212|-80.497332|33|35.667941|CONDENSED SOUP|1.84|1|CAMP HLTHY REQ GOLDEN MUSHROOM|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00051000207852|SOUP|G1 GROCERY|-80.497332|1.4049434824709919|178|2
35.667941|f335429f050baff3de81db38c0d3ed8972262460|4.78|2014-11-16 19:01:00|1.4057311447477159|2|7203663217|178|0.6225230078570788|0|52|330|-80.497332|55|35.667941|EGGS|0.78|3|HT GRADE A LARGE EGGS 18 CT|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00072036632173|EGGS FRESH|DAIRY|-80.497332|1.4049434824709919|178|2
35.667941|6770f3aa2e17157022a43275004b75f0eac06a0e|3.49|2014-11-09 20:48:00|1.4057311447477159|2|2840008294|178|0.6225230078570788|0|52|201|-80.497332|31|35.667941|POTATO CHIPS|0.99|1|LAYS KETTLE JALAPENO|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00028400082907|SNACKS|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|e82254b0471247a5778a390732ecaa617e217bd7|1.5|2015-01-28 14:28:00|1.4057311447477159|2|20563700000|178|0.6225230078570788|0|52|1823|-80.497332|410|35.667941|BH HAM|0.0|6|BOARS HEAD SWEET SLICE HAM|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00205629000008|BH MEAT|DELI|-80.497332|1.4049434824709919|178|1
35.667941|a6528289ac4bbed73f17273231bee318d6b1426b|7.98|2015-03-09 19:26:00|1.4057311447477159|2|4470001120|178|0.6225230078570788|0|52|838|-80.497332|102|35.667941|PEGS|2.0|19|OSCAR MAYER BEEF SALAMI|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00044700011201|LUNCHMEATS|CASE READY MEATS|-80.497332|1.4049434824709919|178|2
35.667941|37290c9512c5ea602830b6d8235d0bc20ee94dbe|7.42|2014-11-03 19:31:00|1.4057311447477159|2||178|0.6225230078570788|0|52|500|-80.497332|64|35.667941|FRESH APPLES|3.73|4|BRAEBURN APPLES|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00204103000008|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|5b7c770eac0f6f8cf1c972ddaaa7dd7325b0cfdf|7.96|2015-01-12 19:45:00|1.4057311447477159|2|7203663220|178|0.6225230078570788|0|52|330|-80.497332|55|35.667941|EGGS|2.96|3|HT GRADE A    LARGE EGGS|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00072036632203|EGGS FRESH|DAIRY|-80.497332|1.4049434824709919|178|4
35.667941|712c836cd11be34983eb82f4ef48a8754f4ba10a|5.98|2015-02-28 17:57:00|80.497482303704658|2|3338365583|178|35.7478645851604|0|6|522|-80.780702|64|35.318911|FRESH TOMATOES|0.98|4|SWEET GRAPE TOMATO (PINT)|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|35.699188602026126|00814369011214|FRESH PRODUCE|PRODUCE|-80.497332|80.497816662899567|167|2
35.667941|e635ec739df754695fbde8990324ee2aa8c3df7d|27.17|2015-02-14 14:23:00|80.497482303704658|2|20302800000|178|35.7478645851604|0|6|652|-80.780702|141|35.318911|FRESH LAMB PRIMALS|0.0|2|LAMB BONELESS BUTTERFLIED LEG|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|35.699188602026126|00203028000001|LAMB|MEAT|-80.497332|80.497816662899567|167|1
35.667941|22b68080746f420e0226ba70caeff43f3754c312|7.58|2014-10-28 16:22:00|1.4057311447477159|2|2500005542|178|0.6225230078570788|0|52|335|-80.497332|56|35.667941|ORANGE JUICE-REGRIGERATED|0.79|3|SIMPLY ORANGE ORIGINAL|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00025000055423|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.497332|1.4049434824709919|178|2
35.667941|d8e4968663e5c4b84baeb1b76c2a5a5ff392956a|14.03|2014-12-29 15:24:00|1.4057311447477159|2|20576900000|178|0.6225230078570788|0|52|1820|-80.497332|410|35.667941|BH BEEF|0.0|6|BOARS HEAD DELUXE ROAST BEEF|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00205769000005|BH MEAT|DELI|-80.497332|1.4049434824709919|178|1
35.667941|81b134915ac1ea78b35af33ac8788b0d87355500|19.81|2015-01-20 19:28:00|1.4057311447477159|2|20894700000|178|0.6225230078570788|0|52|977|-80.497332|201|35.667941|FRESH HT CHICKEN|9.379999999999999|2|HT WHOLE CHICKEN|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00208947000002|POULTRY|MEAT|-80.497332|1.4049434824709919|178|2
35.667941|8dc2be31a54a9349afb7a15e0b73f3c26c391408|23.9|2014-10-13 19:34:00|1.4057311447477159|2|20894700000|178|0.6225230078570788|0|52|977|-80.497332|201|35.667941|FRESH HT CHICKEN|11.31|2|HT WHOLE CHICKEN|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00208947000002|POULTRY|MEAT|-80.497332|1.4049434824709919|178|3
35.667941|e681a80ce304aa07eec886d4e8c693e4473482a9|3.79|2014-11-24 13:50:00|1.4057311447477159|2|5210000698|178|0.6225230078570788|0|52|1245|-80.497332|34|35.667941|SINGLE SPICES|0.0|1|MC BAY LEAVES|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00052100006987|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|8cb3f0f3bebe798d8b21f48ebf2e97c03c3f53af|4.85|2014-12-26 13:38:00|1.4057311447477159|2|7790011553|178|0.6225230078570788|0|52|361|-80.497332|105|35.667941|BREAKFAST SAUSAGE|1.51|19|JIMMY DEAN HOT SAUSAGE|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00077900115639|BREAKFAST SAUSAGE|CASE READY MEATS|-80.497332|1.4049434824709919|178|1
35.667941|e6288be41679a168ace143eb30a8754ae5352862|3.59|2015-03-02 20:15:00|1.4057311447477159|2|3500046112|178|0.6225230078570788|0|52|725|-80.497332|66|35.667941|NFS-DISHWASHING LIQUID|0.0|1|PALMOLIVE LIQ DISH ORIGINAL|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00035000461124|DETERGENTS|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|e38af275df8f175bca80b94fc19ef5ec44818b86|9.7|2014-11-03 15:43:00|1.4057311447477159|2|3450015136|178|0.6225230078570788|0|52|312|-80.497332|51|35.667941|BUTTER|0.86|3|L O L UNSALTED BUTTER QUARTERS|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00034500151504|BUTTER & MARGARINE|DAIRY|-80.497332|1.4049434824709919|178|2
35.667941|9728e7388ab5911413edc933659ed970e826298d|4.49|2015-01-24 17:08:00|1.4057311447477159|2|4812127707|178|0.6225230078570788|0|52|1036|-80.497332|164|35.667941|BREAKFAST BAGELS|2.25|7|THOMAS  RAISIN BAGELS 6CT PP|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00048121292089|BREAKFAST|COMMERCIAL BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|428ab3f509faa600413b44173d7dea765a64fcf4|3.79|2014-10-31 13:01:00|1.4057311447477159|2|4138309010|178|0.6225230078570788|0|52|1263|-80.497332|57|35.667941|GOOD FOR YOU MILK|0.0|3|LACTAID CAL FORT F F HALF GAL|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00041383090219|MILK|DAIRY|-80.497332|1.4049434824709919|178|1
35.667941|325040db57e271b8abaaaef2c175bd223cb28b9b|4.99|2015-01-07 16:03:00|1.4057311447477159|2|7203688138|178|0.6225230078570788|0|52|500|-80.497332|64|35.667941|FRESH APPLES|0.0|4|HT CRIPPS PINK APPLE 3LB|a54094fdd3cc6a2abd74855f25d528634d68ad75|5.522593675939065|0.6209993146566879|00072036881380|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.116638|58c12784487f734ebb2367dd40a13677c5d8d998|9.97|2014-09-12 14:48:00|80.856688219393845|1|7214011020|204|35.136548651953511|0|15|3202|-80.825175|1015|35.152722|HAND & BODY THERAPEUTIC|0.0|17|EUCERIN SMTHING ESS BDY LOTION|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00072140634827|HAND & BODY LOTION/SUN CARE|HBC|-80.85753|80.857542703059863|160|1
35.116638|7ecccfa26f6925ffc24defc3e05abd81e6a40a73|3.49|2014-11-10 14:04:00|80.856688219393845|1|7341013546|204|35.136548651953511|0|15|1035|-80.825175|163|35.152722|SANDWICH ROLL|0.0|7|ARN HNY WHEAT SANDWICH THIN PP|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00073410135433|BUNS/ROLLS|COMMERCIAL BAKERY|-80.85753|80.857542703059863|160|1
35.116638|20e5830a98ddcbf46f94875d2f8c021cbc4cdd4f|4.99|2015-02-18 10:59:00|80.856688219393845|1|7203688143|204|35.136548651953511|0|15|561|-80.825175|64|35.152722|FR PROD ORGANIC PRODUCE|1.0|4|ORG HT SPRING MIX 11 OZ|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00072036881434|FRESH PRODUCE|PRODUCE|-80.85753|80.857542703059863|160|1
35.116638|1a53e757c85a9d6ea1639fe24c984a3563e8940c|2.0|2015-01-02 11:56:00|80.856688219393845|1||204|35.136548651953511|0|15|511|-80.825175|64|35.152722|FRESH AVOCADOS|0.11|4|AVOCADOS, HASS XL 36CT|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00204770000004|FRESH PRODUCE|PRODUCE|-80.85753|80.857542703059863|160|1
35.116638|9a23233fd4a57b40c39fa2c4b93541bddda837d7|2.0|2015-01-14 11:15:00|80.856688219393845|1||204|35.136548651953511|0|15|511|-80.825175|64|35.152722|FRESH AVOCADOS|0.11|4|AVOCADOS, HASS XL 36CT|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00204770000004|FRESH PRODUCE|PRODUCE|-80.85753|80.857542703059863|160|1
35.116638|4f8d2ecb23427401c2bc5057d8be3fd96325ce43|3.19|2014-12-03 11:18:00|80.856688219393845|1|2220094152|204|35.136548651953511|0|15|3876|-80.825175|1070|35.152722|SOLID-MALE|0.0|17|SPEED STK IRISH SPRING ORIG AP|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00022200950367|DEODORANT|HBC|-80.85753|80.857542703059863|160|1
35.116638|6f948c485ac843ba11a726cb8219576e8e65fea4|4.99|2014-09-16 14:02:00|80.856688219393845|1|3800031834|204|35.136548651953511|0|15|74|-80.825175|9|35.152722|RTE CEREAL ALL FAMILY|0.0|1|KELL MINI WHEATS BITE LG BOX|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00038000318344|CEREAL|G1 GROCERY|-80.85753|80.857542703059863|160|1
35.116638|56a5aaf7e43d2743d35d8cf1526e1bef7391767b|3.59|2015-03-03 13:21:00|80.856688219393845|1|4000024906|204|35.136548651953511|0|15|46|-80.825175|7|35.152722|PKG CHOC|0.0|1|M&M PEANUT BUTTER|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00040000250104|CANDY|G1 GROCERY|-80.85753|80.857542703059863|160|1
35.116638|da2568b69f0cc74c995fcfb9974866e973d12d83|6.78|2014-09-14 12:39:00|80.856688219393845|1|4000024906|204|35.136548651953511|0|15|46|-80.825175|7|35.152722|PKG CHOC|0.0|1|M&M PEANUT BUTTER|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00040000250104|CANDY|G1 GROCERY|-80.85753|80.857542703059863|160|2
35.116638|e0ed3d7f801c43df24286d4849e2c6262f7f7866|4.99|2014-11-28 12:11:00|80.856688219393845|1|7597140209|204|35.136548651953511|0|15|1845|-80.825175|425|35.152722|FFM PRESLICED CHEESE|0.0|6|F.F. MUENSTER CHEESE|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00072036010322|PRESLICED CHEESE|DELI|-80.85753|80.857542703059863|160|1
35.116638|a0b6be9f1073a2d71b33bc0c1b6c2f48665ebb00|2.4|2015-02-15 15:42:00|80.856688219393845|1|7047000641|204|35.136548650866018|0|15|687|-80.848528|61|35.053394|BLENDED|0.0|3|YOPLAIT T/C KEY LIME PIE|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00070470180823|YOGURT|DAIRY|-80.85753|80.857545036815822|11|4
35.116638|167a8578f1cd283769518cb2fa933205589517bf|3.35|2015-01-27 11:57:00|80.856688219393845|1|3700022205|204|35.136548651953511|0|15|725|-80.825175|66|35.152722|NFS-DISHWASHING LIQUID|0.0|1|DAWN LIQ DISH ANTIBAC APPLE BL|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00037000222026|DETERGENTS|G1 GROCERY|-80.85753|80.857542703059863|160|1
35.116638|f2ba0173e704967288e555e2cab1e973ffdafd55|5.98|2014-10-11 13:11:00|80.856688219393845|1|81204900640|204|35.136548651953511|0|15|504|-80.825175|64|35.152722|FRESH BERRIES|0.0|4|BLUEBERRIES 6 OZ|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00033383220222|FRESH PRODUCE|PRODUCE|-80.85753|80.857542703059863|160|2
35.116638|8c568a2d4172e7f63784a7561c9d62c9000e00cf|4.99|2015-01-23 13:13:00|80.856688219393845|1|3800001621|204|35.136548651953511|0|15|61|-80.825175|9|35.152722|RTE CEREAL ADULT|0.0|1|KELLOGG SPECIAL K 18|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00038000016219|CEREAL|G1 GROCERY|-80.85753|80.857542703059863|160|1
35.116638|67fd4680739982979b5f7d20cd836206009cab0a|6.99|2015-02-02 12:52:00|80.856688219393845|1|4900002890|204|35.136548651953511|0|15|54|-80.825175|8|35.152722|DIET|0.0|23|CF DIET COKE 12 OZ 12 PK FP CN|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00049000029345|CARBONATED BEVERAGES|BEVERAGE|-80.85753|80.857542703059863|160|1
35.116638|5373e7f8ec363efe7a68ef34054ebfab568a31e1|6.79|2014-10-17 14:44:00|80.856688219393845|1|4900002890|204|35.136548651953511|0|15|54|-80.825175|8|35.152722|DIET|1.8|23|CF DIET COKE 12 OZ 12 PK FP CN|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00049000029345|CARBONATED BEVERAGES|BEVERAGE|-80.85753|80.857542703059863|160|1
35.116638|24c415b4b36caba55ea2b79972b388798459a5be|6.79|2014-11-24 14:23:00|80.856688219393845|1|4900002890|204|35.136548651953511|0|15|54|-80.825175|8|35.152722|DIET|1.8|23|CF DIET COKE 12 OZ 12 PK FP CN|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00049000029345|CARBONATED BEVERAGES|BEVERAGE|-80.85753|80.857542703059863|160|1
35.116638|23634d2480ad195a33422b71681311ac18e2aecd|6.79|2014-12-17 11:44:00|80.856688219393845|1|4900002890|204|35.136548651953511|0|15|54|-80.825175|8|35.152722|DIET|0.0|23|CF DIET COKE 12 OZ 12 PK FP CN|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00049000029345|CARBONATED BEVERAGES|BEVERAGE|-80.85753|80.857542703059863|160|1
35.116638|b060b1a42827e9c6b76296fa14ef23b2b4b22204|6.99|2015-01-03 15:33:00|80.856688219393845|1|4900002890|204|35.136548651953511|0|15|54|-80.825175|8|35.152722|DIET|2.0|23|CF DIET COKE 12 OZ 12 PK FP CN|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00049000029345|CARBONATED BEVERAGES|BEVERAGE|-80.85753|80.857542703059863|160|1
35.116638|f3640b295d93f8fb75a755e983105842eeb3f76d|6.79|2014-10-07 14:22:00|80.856688219393845|1|4900002890|204|35.136548651953511|0|15|54|-80.825175|8|35.152722|DIET|1.8|23|CF DIET COKE 12 OZ 12 PK FP CN|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00049000029345|CARBONATED BEVERAGES|BEVERAGE|-80.85753|80.857542703059863|160|1
35.116638|f56080beb56da37754e2cee04f86418f0cab7d75|6.99|2015-01-07 11:02:00|80.856688219393845|1|4900002890|204|35.136548651953511|0|15|54|-80.825175|8|35.152722|DIET|2.0|23|CF DIET COKE 12 OZ 12 PK FP CN|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00049000029345|CARBONATED BEVERAGES|BEVERAGE|-80.85753|80.857542703059863|160|1
35.116638|05fbedae7e26b985630c71ba3fbf630dc59949df|6.79|2014-09-29 14:12:00|80.856688219393845|1|4900002890|204|35.136548651953511|0|15|54|-80.825175|8|35.152722|DIET|1.8|23|CF DIET COKE 12 OZ 12 PK FP CN|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00049000029345|CARBONATED BEVERAGES|BEVERAGE|-80.85753|80.857542703059863|160|1
35.116638|e8f7cd83ffadf3e9457805c8a679c4f5fdbed72d|6.99|2015-02-12 14:52:00|80.856688219393845|1|4900002890|204|35.136548651953511|0|15|54|-80.825175|8|35.152722|DIET|2.0|23|CF DIET COKE 12 OZ 12 PK FP CN|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00049000029345|CARBONATED BEVERAGES|BEVERAGE|-80.85753|80.857542703059863|160|1
35.116638|e1d0feace5804ab1c5877068d329dab563784919|6.79|2014-11-19 11:45:00|80.856688219393845|1|4900002890|204|35.136548651953511|0|15|54|-80.825175|8|35.152722|DIET|1.8|23|CF DIET COKE 12 OZ 12 PK FP CN|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00049000029345|CARBONATED BEVERAGES|BEVERAGE|-80.85753|80.857542703059863|160|1
35.116638|c7bbda38ef28a11dab66bf4306dcc6f5279fa526|6.79|2014-12-08 14:02:00|80.856688219393845|1|4900002890|204|35.136548652122933|0|15|54|-80.849471|8|35.161696|DIET|1.8|23|CF DIET COKE 12 OZ 12 PK FP CN|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00049000029345|CARBONATED BEVERAGES|BEVERAGE|-80.85753|80.857542299675529|35|1
35.116638|66a3f0b93f4d5e0f12cda81aae084a14877c7d51|6.79|2014-10-25 15:14:00|80.856688219393845|1|4900002890|204|35.136548651953511|0|15|54|-80.825175|8|35.152722|DIET|1.8|23|CF DIET COKE 12 OZ 12 PK FP CN|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00049000029345|CARBONATED BEVERAGES|BEVERAGE|-80.85753|80.857542703059863|160|1
35.116638|1d76ca8f0e070fde93072494903364153d2fff69|1.69|2014-11-17 15:50:00|80.856688219393845|1|3660207290|204|35.136548651953511|0|15|4207|-80.825175|1200|35.152722|COUGH DROP-ADULT|0.85|17|RICOLA ECH. HONEY LEMN -30146|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00036602301467|COUGH/COLD/SINUS|HBC|-80.85753|80.857542703059863|160|1
35.116638|c1589cc866f22e59652d519d0dc82b3914877069|3.49|2014-12-14 14:02:00|80.856688219393845|1|3800001611|204|35.136548652122933|0|15|61|-80.849471|9|35.161696|RTE CEREAL ADULT|0.0|1|KELLOGG SPECIAL K 12 OZ BOX|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00038000016110|CEREAL|G1 GROCERY|-80.85753|80.857542299675529|35|1
35.116638|83a8c9fc0435bdcc4642fa3a0f2e417bd04311fc|3.49|2015-02-06 10:06:00|80.856688219393845|1|3800001611|204|35.136548651953511|0|15|61|-80.825175|9|35.152722|RTE CEREAL ADULT|0.0|1|KELLOGG SPECIAL K 12 OZ BOX|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00038000016110|CEREAL|G1 GROCERY|-80.85753|80.857542703059863|160|1
35.116638|b6185da2545e29972db0b2c58101a5d1591b9839|2.79|2014-12-23 13:40:00|80.856688219393845|1|5100014880|204|35.136548652122933|0|15|1499|-80.849471|33|35.161696|RTS MICROWAVE|0.0|1|CHUNKY MW CHILI ROADHOUSE|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00051000159045|SOUP|G1 GROCERY|-80.85753|80.857542299675529|35|1
35.116638|849903541c3a3a6d0ca4d31bf98dfed4049b43f7|30.29|2014-11-12 14:25:00|80.856688219393845|1|35058072638|204|35.136548651953511|0|15|4189|-80.825175|1200|35.152722|ALLERGY REMEDY-CHILDREN|0.0|17|L ZYRTEC ALLERGY LIQUIGELS|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00300450204448|COUGH/COLD/SINUS|HBC|-80.85753|80.857542703059863|160|1
35.116638|a5df3979e90a1e0f91b54105ca683ab863e6600b|3.96|2014-09-22 14:11:00|80.856688219393845|1|20596200000|204|35.136548651953511|0|15|1821|-80.825175|410|35.152722|BH TURKEY|0.0|6|BOARS HEAD MAPLE HONEY TURKEY|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00205962000000|BH MEAT|DELI|-80.85753|80.857542703059863|160|1
35.116638|14a397959c037498fdbfe67aefee31caed4ba51b|2.97|2014-10-15 11:45:00|80.856688219393845|1|20596200000|204|35.136548651953511|0|15|1821|-80.825175|410|35.152722|BH TURKEY|0.0|6|BOARS HEAD MAPLE HONEY TURKEY|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00205962000000|BH MEAT|DELI|-80.85753|80.857542703059863|160|1
35.116638|217ad4d3e92f9f6a9389aeb418a5ca1951abc2d8|5.06|2014-10-27 11:04:00|80.856688219393845|1|20596200000|204|35.136548651953511|0|15|1821|-80.825175|410|35.152722|BH TURKEY|0.92|6|BOARS HEAD MAPLE HONEY TURKEY|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00205962000000|BH MEAT|DELI|-80.85753|80.857542703059863|160|1
35.116638|c82908c59f7f57579b8722e7c4c4b63bf1127fb9|1.03|2014-10-30 14:22:00|80.856688219393845|1||204|35.136548651953511|0|15|502|-80.825175|64|35.152722|FRESH BANANAS|0.0|4|BANANAS, YELLOW|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00204011000008|FRESH PRODUCE|PRODUCE|-80.85753|80.857542703059863|160|1
35.116638|f7a32681ca3fc17821c802d877758d3d10277afa|0.64|2014-09-25 11:33:00|80.856688219393845|1||204|35.136548651953511|0|15|502|-80.825175|64|35.152722|FRESH BANANAS|0.0|4|BANANAS, YELLOW|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00204011000008|FRESH PRODUCE|PRODUCE|-80.85753|80.857542703059863|160|1
35.116638|4bff112d41eb9e38e21f7e942c086f4571d5c9fa|0.67|2014-10-01 11:07:00|80.856688219393845|1||204|35.136548651953511|0|15|502|-80.825175|64|35.152722|FRESH BANANAS|0.0|4|BANANAS, YELLOW|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00204011000008|FRESH PRODUCE|PRODUCE|-80.85753|80.857542703059863|160|1
35.116638|e332a1624d7c1f70baf6fd707508740f6d857e22|3.99|2014-11-05 13:14:00|80.856688219393845|1|71575620002|204|35.136548651953511|0|15|504|-80.825175|64|35.152722|FRESH BERRIES|0.2|4|STRAWBERRIES 1LB CLAM|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00715756200023|FRESH PRODUCE|PRODUCE|-80.85753|80.857542703059863|160|1
35.116638|f1b5259f1b53f59356a44129e7e11b9136c12588|5.98|2014-11-14 14:17:00|80.856688219393845|1|81204900640|204|35.136548651953511|0|15|504|-80.825175|64|35.152722|FRESH BERRIES|0.0|4|BLUEBERRIES 6 OZ|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00033383222288|FRESH PRODUCE|PRODUCE|-80.85753|80.857542703059863|160|2
35.116638|989de0c7643417841758125a1871b5abac924940|4.58|2014-10-21 11:28:00|80.856688219393845|1|3660207290|204|35.136548651953511|0|15|4207|-80.825175|1200|35.152722|COUGH DROP-ADULT|1.4|17|RICOLA SF LEMON MINT -19210|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00036602192102|COUGH/COLD/SINUS|HBC|-80.85753|80.857542703059863|160|2
35.116638|cded653231b1b6788118be5d059f10fb7128145d|5.07|2014-10-04 13:34:00|80.856688219393845|1|3660207290|204|35.136548651953511|0|15|4207|-80.825175|1200|35.152722|COUGH DROP-ADULT|0.0|17|RICOLA SF LEMON MINT -19210|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00036602192102|COUGH/COLD/SINUS|HBC|-80.85753|80.857542703059863|160|3
35.116638|723096d5a0a1db141b82f4467014c33d6706c456|3.19|2015-01-24 11:40:00|80.856688219393845|1|5113199525|204|35.136548651953511|0|15|4816|-80.825175|1235|35.152722|FIRST AID ADHESIVE BANDG|0.0|17|NEXCARE WATERPROOF CLR ONE SZE|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00051131995253|FIRST AID|HBC|-80.85753|80.857542703059863|160|1
35.116638|adc03b9483e5549fd86ea3243a2e0e82fa07a549|1.01|2015-02-20 11:35:00|80.856688219393845|1||204|35.136548651953511|0|15|502|-80.825175|64|35.152722|FRESH BANANAS|0.0|4|BANANAS, YELLOW|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00204011000008|FRESH PRODUCE|PRODUCE|-80.85753|80.857542703059863|160|1
35.116638|3e3bb640a4f8b5795f3e65ff03a1bb4de9545582|4.49|2014-11-12 14:19:00|80.856688219393845|1|7203001339|204|35.136548651953511|0|15|1685|-80.825175|385|35.152722|ENTENMANNS (SWEET GOODS)|0.0|14|ENT LB MINI FUDGE BROWNIES PP|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00072030013428|SWEET GOODS|BAKERY|-80.85753|80.857542703059863|160|1
35.116638|c2bb8412487af805e8cb618ec75a03bd50c3d205|2.29|2015-02-04 16:53:00|80.856688219393845|1|7203663996|204|35.136548652122933|0|15|342|-80.849471|57|35.161696|FRESH MILK|0.0|3|HARRIS TEETER 1%  MILK|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00072036631305|MILK|DAIRY|-80.85753|80.857542299675529|35|1
35.116638|6dedd71a497fae9eb2a680fc3e1572fb1c8f48fb|3.99|2015-02-25 09:55:00|80.856688219393845|1|7433610006|204|35.136548651953511|0|15|342|-80.825175|57|35.152722|FRESH MILK|0.0|3|HUNTER 1%  MILK  GALLON|a7bdd9d485ca9712eae0ec1f97820f0d2a0f189c|1.375778154788002|35.134355925261694|00074336100291|MILK|DAIRY|-80.85753|80.857542703059863|160|1
35.667941|a99b761712d66fb3db5a51e1dd5a8fe4f7c8c090|3.97|2015-03-08 19:50:00|1.4057311447477159|4|7203625034|178|0.6225230078570788|0|52|144|-80.497332|229|35.667941|CEAMERS-POWDERED|0.0|1|(U)HT NON DAIRY CREAMER|a9ef6aa9bcc45165f791c18fde47c679ada911a0|5.395443491535754|0.6209993146566879|00072036250346|COCOAS CREAMERS SYRUPS|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|de2e125c6966ee0dff541fb0e07c6fe9d4691558|3.19|2014-10-08 16:46:00|1.4057311447477159|4|7203656061|178|0.6225230078570788|0|52|320|-80.497332|53|35.667941|COTTAGE CHEESE|0.69|3|HT COTTAGE CHEESE|a9ef6aa9bcc45165f791c18fde47c679ada911a0|5.395443491535754|0.6209993146566879|00072036560612|CULTURES|DAIRY|-80.497332|1.4049434824709919|178|1
35.667941|a8d01fd11df0f9d6995655c0ab770a2c875abe12|0.97|2014-11-23 13:02:00|1.4057311447477159|4|7203637031|178|0.6225230078570788|0|52|212|-80.497332|33|35.667941|CONDENSED SOUP|0.17|1|HT SP HLTHY CRM MUSHROOM|a9ef6aa9bcc45165f791c18fde47c679ada911a0|5.395443491535754|0.6209993146566879|00072036370389|SOUP|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|5b41856ddabe3a9fc20dc08614f481d4be908846|14.7|2014-12-20 14:53:00|1.4057311447477159|4|4470002268|178|0.6225230078570788|0|52|358|-80.497332|100|35.667941|REGULAR BACON|3.68|19|OSCAR MAYER SLICED BACON|a9ef6aa9bcc45165f791c18fde47c679ada911a0|5.395443491535754|0.6209993146566879|00044700019887|BACON|CASE READY MEATS|-80.497332|1.4049434824709919|178|2
35.667941|d8e5da36352da4c2d4765052c11ca239852f600d|2.29|2015-01-31 15:09:00|1.4057311447477159|4|7203663996|178|0.6225230078570788|0|52|342|-80.497332|57|35.667941|FRESH MILK|0.82|3|HARRIS TEETER 2%   MILK|a9ef6aa9bcc45165f791c18fde47c679ada911a0|5.395443491535754|0.6209993146566879|00072036639998|MILK|DAIRY|-80.497332|1.4049434824709919|178|1
35.667941|25a3ad58e3d192ce1c9160f0fb02f5793ad69d87|4.19|2014-11-16 20:09:00|1.4057311447477159|4|1862770366|178|0.6225230078570788|0|52|61|-80.497332|9|35.667941|RTE CEREAL ADULT|2.22|1|KASHI HEART TO HEART BLUEBERRY|a9ef6aa9bcc45165f791c18fde47c679ada911a0|5.395443491535754|0.6209993146566879|00018627510031|CEREAL|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|5b4bf8781e28372604f51adeaeb47029fc20eab8|7.16|2015-02-06 14:03:00|1.4057311447477159|4|3600025824|178|0.6225230078570788|0|52|424|-80.497332|72|35.667941|NFS-FACIAL TISSUE|2.16|1|KLEENEX TISSUE WHITE 160CT|a9ef6aa9bcc45165f791c18fde47c679ada911a0|5.395443491535754|0.6209993146566879|00036000373905|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.497332|1.4049434824709919|178|4
35.667941|ca7937cecca3e53790b306b373581be76bf9eb93|2.45|2014-10-19 10:09:00|1.4057311447477159|4|7203663217|178|0.6225230078570788|0|52|330|-80.497332|55|35.667941|EGGS|0.45|3|HT GRADE A LARGE EGGS 18 CT|a9ef6aa9bcc45165f791c18fde47c679ada911a0|5.395443491535754|0.6209993146566879|00072036632173|EGGS FRESH|DAIRY|-80.497332|1.4049434824709919|178|1
35.024464|abc19f641f877551ad76aa900b9231b297ddcfc9|1.69|2014-11-20 16:38:00|80.848351720559364|3|7203688003|317|35.05275739545484|0|25|527|-80.994596|64|35.061685|FRESH CARROTS|0.0|4|HT BABY CARROTS 1LB BAG|ab3bc204996fad9f22c7b2f35d6c2708473c6ab8|1.9550053743548932|35.082633588753836|00072036880031|FRESH PRODUCE|PRODUCE|-80.847383|80.847392541820909|475|1
35.024464|b4361f69fa807d2ec80e64b7510787204fd190d1|3.99|2014-09-15 16:32:00|1.41290891556208|3|7127923100|317|0.6112922155462233|0|33|555|-80.847383|64|35.024464|PACKAGED SALADS|0.0|4|F.E. BABY SPRING SALAD MIX|ab3bc204996fad9f22c7b2f35d6c2708473c6ab8|1.9550053743548932|0.61055446569467375|00071279231006|FRESH PRODUCE|PRODUCE|-80.847383|1.4110530249708906|317|1
35.024464|8f31816302570d7192483bfb179cca27e6a3a430|2.29|2014-12-11 18:02:00|1.41290891556208|3|3250004281|317|0.6112922155462233|0|33|100|-80.847383|15|35.024464|CORN MEAL|0.0|1|WHITE LILY BTRMILK CORNMEAL SR|ab3bc204996fad9f22c7b2f35d6c2708473c6ab8|1.9550053743548932|0.61055446569467375|00032500042815|FLOUR|G1 GROCERY|-80.847383|1.4110530249708906|317|1
35.024464|9a8dc33aa6dd1bf0d61f963291c630d406778b79|4.49|2014-09-27 16:11:00|80.848351720559364|3|87989000001|317|35.052757393683848|0|25|1982|-80.97058|480|35.03469|DRY GOODS CRACKERS|0.0|6|ORIGINAL MULTI-SEED CRACKERS|ab3bc204996fad9f22c7b2f35d6c2708473c6ab8|1.9550053743548932|35.082633588753836|00879890000014|DRY GOODS|DELI|-80.847383|80.847398509238786|82|1
35.024464|8cdff01542746f3054a1d348724b93cde8ced293|1.99|2014-11-05 15:46:00|80.848351720559364|3|7044640000|317|35.05275739545484|0|25|498|-80.994596|111|35.061685|PICKLES & SAUERKRAUT|0.49|19|BOARS HEAD SAUERKRAUT 16 OZ|ab3bc204996fad9f22c7b2f35d6c2708473c6ab8|1.9550053743548932|35.082633588753836|00070446400009|MISC. PACKAGED MEATS|CASE READY MEATS|-80.847383|80.847392541820909|475|1
35.024464|43f98514af916d9f6aa8578932b8a6816f81f91f|1.82|2014-10-10 13:17:00|80.848351720559364|3|20575500000|317|35.052757385888057|0|25|1603|-80.837892|371|34.937113|PRIVATE LABEL BREAD|0.0|14|WHEAT BAGUETTE ROUNDS|ab3bc204996fad9f22c7b2f35d6c2708473c6ab8|1.9550053743548932|35.082633588753836|00205760000004|BREAD|BAKERY|-80.847383|80.847412976374386|372|1
35.024464|0c667586be011aef5db5b78e0ed8d465d8ee0ccc|2.53|2014-11-24 14:53:00|1.41290891556208|3||317|0.6112922155462233|0|33|500|-80.847383|64|35.024464|FRESH APPLES|0.0|4|GOLD DEL APPLE, WA 56|ab3bc204996fad9f22c7b2f35d6c2708473c6ab8|1.9550053743548932|0.61055446569467375|00233285000001|FRESH PRODUCE|PRODUCE|-80.847383|1.4110530249708906|317|1
35.024464|48158dc2e6a65eacde3e41133391346946f2f886|3.75|2015-02-28 15:36:00|80.848351720559364|3|97074|317|35.052757385888057|0|25|1597|-80.837892|369|34.937113|NFS BEVERAGE BLEND|0.0|22|MOCHA LIGHT FRAPPUCCINO TALL|ab3bc204996fad9f22c7b2f35d6c2708473c6ab8|1.9550053743548932|35.082633588753836|00000000970740|NFS STARBUCKS|COFFEE SHOP|-80.847383|80.847412976374386|372|1
35.024464|256a27dd21fe65f9cc7353ab29c37b2b465b877e|3.99|2014-12-28 17:02:00|1.41290891556208|3|5783602064|317|0.6112922155462233|0|33|522|-80.847383|64|35.024464|FRESH TOMATOES|0.0|4|CAMPARI TOMATO 16 OZ|ab3bc204996fad9f22c7b2f35d6c2708473c6ab8|1.9550053743548932|0.61055446569467375|00057836020641|FRESH PRODUCE|PRODUCE|-80.847383|1.4110530249708906|317|1
35.024464|fa5074f8d5d79cefb392a1b38dbba075d4e36bcb|2.69|2015-02-28 16:40:00|80.848351720559364|3|7225001739|317|35.052757385888057|0|25|1025|-80.837892|162|34.937113|WHITE|0.5|7|NATOWN WHITEWHEAT RTOP BRD|ab3bc204996fad9f22c7b2f35d6c2708473c6ab8|1.9550053743548932|35.082633588753836|00072250017398|SLICED BREAD|COMMERCIAL BAKERY|-80.847383|80.847412976374386|372|1
35.024464|b4d219e23184b8a619e500bdac243238859c40cf|3.99|2014-10-17 13:46:00|80.848351720559364|3|85609100102|317|35.052757393683848|0|25|3303|-80.97058|1025|35.03469|BATH ACCESSORIES|0.0|17|CLEAN LOGIC BATH BODY SCRUBBER|ab3bc204996fad9f22c7b2f35d6c2708473c6ab8|1.9550053743548932|35.082633588753836|00856091001026|BATH PRODUCTS|HBC|-80.847383|80.847398509238786|82|1
35.024464|a5670d4e702bce083470846f956b0ca05d1967d4|3.49|2014-12-18 15:36:00|80.848351720559364|3|7203695248|317|35.052757393683848|0|25|1611|-80.97058|371|35.03469|PITA'S AND FLAT BREADS|0.0|14|FFM WHITE FLATBREADS ROUNDS|ab3bc204996fad9f22c7b2f35d6c2708473c6ab8|1.9550053743548932|35.082633588753836|00072036954152|BREAD|BAKERY|-80.847383|80.847398509238786|82|1
35.442529|1f1c81d0cb452d828e3d6a69dd46236266ab2c06|1.2|2014-10-28 21:41:00|1.4102725052409182|2|3663203732|471|0.6185888262835733|0|1|685|-80.762919|61|35.442529|GREEK|0.2|3|DANNON LNF GREEK TSTED COCONUT|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00036632037374|YOGURT|DAIRY|-80.762919|1.4095788500714863|471|1
35.442529|ad32495dddcbbf8c0ed0694eec4f058c7c790b93|2.63|2014-12-12 17:55:00|1.4102725052409182|2||471|0.6185888262835733|0|1|500|-80.762919|64|35.442529|FRESH APPLES|1.32|4|BRAEBURN APPLES|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00204103000008|FRESH PRODUCE|PRODUCE|-80.762919|1.4095788500714863|471|1
35.442529|b72a60380ecda4ea24d81bf10a18fb3c33d75570|4.0|2014-10-24 18:21:00|1.4102725052409182|2||471|0.6185888262835733|0|1|511|-80.762919|64|35.442529|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00204770000004|FRESH PRODUCE|PRODUCE|-80.762919|1.4095788500714863|471|2
35.442529|c141466d50f1221e32aa7d7e90f769aa3a2202c8|3.69|2015-03-05 22:30:00|1.4102725052409182|2|38151905501|471|0.6185888262835733|0|1|3500|-80.762919|1045|35.442529|CONDITIONER-MID PRICE|0.7|17|HERBAL ESS CND HELLO HYDRATION|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00381519055027|HAIR & SCALP CARE|HBC|-80.762919|1.4095788500714863|471|1
35.442529|805dd3f1fbec74a8045a39525f621e440a970421|4.0|2015-01-05 18:27:00|1.4102725052409182|2||471|0.6185888262835733|0|1|511|-80.762919|64|35.442529|FRESH AVOCADOS|0.11|4|AVOCADOS, HASS XL 36CT|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00204770000004|FRESH PRODUCE|PRODUCE|-80.762919|1.4095788500714863|471|2
35.442529|72322061ea9a1f0a92c40bc110a531e103f49bb5|6.75|2014-12-09 21:05:00|80.749667378538092|2|20576400000|471|35.462678055724602|0|3|1820|-80.662946|410|35.412407|BH BEEF|0.0|6|BOARS HEAD PASTRAMI|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|35.465179900649026|00205764000000|BH MEAT|DELI|-80.762919|80.762922535933214|68|1
35.442529|3af9b99fec3fcf795bc01cae39db90581a17db8e|6.37|2015-02-05 17:54:00|1.4102725052409182|2|20576400000|471|0.6185888262835733|0|1|1820|-80.762919|410|35.442529|BH BEEF|0.0|6|BOARS HEAD PASTRAMI|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00205764000000|BH MEAT|DELI|-80.762919|1.4095788500714863|471|1
35.442529|f7ad22b5457d5b27b7b63cb2149171f782bda8ba|5.19|2015-01-09 21:12:00|1.4102725052409182|2|79951201201|471|0.6185888262835733|0|1|276|-80.762919|45|35.442529|ICE MILK/SHERBET/YOGURT-FROZEN|0.0|5|CIAO BELLA BART PEAR HIBIS SOR|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00799512012167|ICE CREAM|FROZEN|-80.762919|1.4095788500714863|471|1
35.442529|a018f5ec2bc4925c782caeda3bb4095be2bf4eb6|6.38|2014-11-16 20:22:00|80.749667378538092|2|61126971646|471|35.462678055618937|0|3|97|-80.746334|8|35.41832|ENERGY DRINKS|1.38|23|CB RED BULL SF 12 OZ CAN|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|35.465179900649026|00611269716467|CARBONATED BEVERAGES|BEVERAGE|-80.762919|80.762923349742664|190|2
35.442529|5a776703070b4a54050768f7ad18bbb25552e7ea|14.27|2015-01-23 19:47:00|1.4102725052409182|2|20949900000|471|0.6185888262835733|0|1|883|-80.762919|145|35.442529|SHRIMP FARM RAISED|8.16|12|51/60 CT EZ PEEL WHITE SHRIMP|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00209499000007|SHRIMP|SEAFOOD|-80.762919|1.4095788500714863|471|1
35.442529|514a852eb9369ad81572101554003a6b1c2fab15|2.4|2015-01-11 14:02:00|80.749667378538092|2||471|35.462678055660284|0|3|531|-80.860108|64|35.500972|FRESH CORN|0.0|4|COO YELLOW CORN|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|35.465179900649026|00204078000003|FRESH PRODUCE|PRODUCE|-80.762919|80.762923050859683|268|3
35.442529|5bd904cf1f66b460b4f2ed0ef3b37007d0b90754|2.4|2015-03-06 20:35:00|80.749667378538092|2||471|35.462678055660284|0|3|531|-80.860108|64|35.500972|FRESH CORN|0.0|4|COO YELLOW CORN|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|35.465179900649026|00204078000003|FRESH PRODUCE|PRODUCE|-80.762919|80.762923050859683|268|4
35.442529|31ce630f2e0ceafdd53e351c9a4d64134f238268|4.0|2015-02-07 20:55:00|1.4102725052409182|2||471|0.6185888262835733|0|1|531|-80.762919|64|35.442529|FRESH CORN|0.0|4|COO YELLOW CORN|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00204078000003|FRESH PRODUCE|PRODUCE|-80.762919|1.4095788500714863|471|5
35.442529|42d31ccd0e384c66e294be3200170bfce039316d|7.14|2014-10-26 20:29:00|80.749667378538092|2|20557100000|471|35.462678055724602|0|3|1820|-80.662946|410|35.412407|BH BEEF|0.0|6|BOARS HEAD LONDON BROIL|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|35.465179900649026|00205571000002|BH MEAT|DELI|-80.762919|80.762922535933214|68|1
35.442529|f568e526acd16106d0984163f0062e0f93694869|12.99|2015-02-22 18:38:00|80.749667378538092|2|20557100000|471|35.462678055618937|0|3|1820|-80.746334|410|35.41832|BH BEEF|0.0|6|BOARS HEAD LONDON BROIL|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|35.465179900649026|00205571000002|BH MEAT|DELI|-80.762919|80.762923349742664|190|1
35.442529|6d94d7f567935ce6556669a799d8c39b0a9021e2|1.68|2015-02-25 20:02:00|80.749667378538092|2||471|35.462678055660284|0|3|522|-80.860108|64|35.500972|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|35.465179900649026|00204664000004|FRESH PRODUCE|PRODUCE|-80.762919|80.762923050859683|268|1
35.442529|1c980929efa175b2d5967e3ef40e9e2ec87f5cfa|1.74|2014-10-05 21:01:00|80.749667378538092|2||471|35.462678055724602|0|3|522|-80.662946|64|35.412407|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|35.465179900649026|00204664000004|FRESH PRODUCE|PRODUCE|-80.762919|80.762922535933214|68|1
35.442529|1534192136e45ba2817751c1e89f41c96c8cf083|1.82|2014-12-30 21:21:00|1.4102725052409182|2||471|0.6185888262835733|0|1|522|-80.762919|64|35.442529|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00204664000004|FRESH PRODUCE|PRODUCE|-80.762919|1.4095788500714863|471|1
35.442529|7a33001d31a3e053737351c58fb02f4d58b44282|0.67|2014-12-31 13:41:00|80.749667378538092|2|7203641111|471|35.462678055618937|0|3|242|-80.746334|39|35.41832|CANNED BEANS|0.05|1|HT PEAS BLACKEYE|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|35.465179900649026|00072036411143|VEGETABLES-CAN/JAR|G1 GROCERY|-80.762919|80.762923349742664|190|1
35.442529|0ed97f9c068aba4e685b7fd5884c0c3926a4fef7|2.5|2015-01-07 20:45:00|80.749667378538092|2|7203670633|471|35.462678055660284|0|3|184|-80.860108|28|35.500972|SALAD DRESSINGS-LIQUID|0.25|1|HT ORG DRS MISO GINGER|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|35.465179900649026|00072036706362|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.762919|80.762923050859683|268|1
35.442529|737b7de620f82c110b6fb724ed0edde8794c5c7d|2.39|2014-11-29 16:00:00|1.4102725052409182|2|7320900007|471|0.6185888262835733|0|1|163|-80.762919|25|35.442529|RELISHES|0.0|1|MRS CAMPBELL CHOW CHOW HOT|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00073209000058|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.762919|1.4095788500714863|471|1
35.442529|3757cc2a7c0f95f8915878b0b073b4e6f8923aa0|2.38|2015-02-09 19:35:00|1.4102725052409182|2|3940001747|471|0.6185888262835733|0|1|242|-80.762919|39|35.442529|CANNED BEANS|0.38|1|BUSH BEAN KIDNEY DK|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00039400017349|VEGETABLES-CAN/JAR|G1 GROCERY|-80.762919|1.4095788500714863|471|2
35.442529|4265ab266d694861f66b6434cfbf711dca6f56c3|1.99|2014-12-15 20:51:00|1.4102725052409182|2|4131301242|471|0.6185888262835733|0|1|217|-80.762919|34|35.442529|EXTRACTS FOOD COLORING|0.2|1|FLAVOR KING IMITATION VANILLA|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00041313012427|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.762919|1.4095788500714863|471|1
35.442529|933bc402fa345877c45be8c9251baaf2c0d59d27|3.99|2015-01-01 22:44:00|1.4102725052409182|2|5929057322|471|0.6185888262835733|0|1|92|-80.762919|13|35.442529|REMAINING CRACKERS|0.99|1|CARRS CRACK PEPPER TABLE CRACK|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00059290575927|CRACKERS|G1 GROCERY|-80.762919|1.4095788500714863|471|1
35.442529|39ce27d3035376933e90afa2965595904fef0dbd|9.99|2015-01-29 20:40:00|80.749667378538092|2|7023666067|471|35.462678055724602|0|3|751|-80.662946|87|35.412407|NFS-BOUQUETS|0.0|9|$9.99 ROSE/GERBERA BOUQUET|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|35.465179900649026|00070236660675|FLORAL|FLORAL|-80.762919|80.762922535933214|68|1
35.442529|5ed40b456d5d5ec5803d8268893c5ab96829c1dd|2.99|2014-12-05 18:17:00|1.4102725052409182|2|20443000000|471|0.6185888262835733|0|1|510|-80.762919|64|35.442529|FRESH PINEAPPLE|0.0|4|GOLD PINEAPPLES|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00643126072003|FRESH PRODUCE|PRODUCE|-80.762919|1.4095788500714863|471|1
35.442529|d979b2be9d240e847f4237b11f3c46465d2a87b4|3.39|2014-11-02 20:29:00|1.4102725052409182|2|7203661037|471|0.6185888262835733|0|1|840|-80.762919|102|35.442529|TUBS|0.3|19|HT SMOKED PASTRAMI|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00072036610492|LUNCHMEATS|CASE READY MEATS|-80.762919|1.4095788500714863|471|1
35.442529|2741b72201bb584dfdbf02fb24696bafc7511364|6.98|2015-02-16 17:34:00|1.4102725052409182|2|2500004786|471|0.6185888262835733|0|1|335|-80.762919|56|35.442529|ORANGE JUICE-REGRIGERATED|1.98|3|MINUTE MAID PULP FREE|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00025000047893|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.762919|1.4095788500714863|471|2
35.442529|0925bd7187571bf63a99e27de64d1caf72352ccd|3.99|2014-09-27 15:38:00|1.4102725052409182|2||471|0.6185888262835733|0|1|539|-80.762919|64|35.442529|FRESH CAULIFLOWER|0.0|4|GREEN CAULIFLOWER|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00204567000002|FRESH PRODUCE|PRODUCE|-80.762919|1.4095788500714863|471|1
35.442529|4b7e19fa128ae4d9fc19d5eee7ffdaba1390d9e0|3.49|2014-12-11 20:50:00|1.4102725052409182|2|4460000889|471|0.6185888262835733|0|1|400|-80.762919|69|35.442529|NFS-LIQUID CLEANERS|0.49|1|FORMULA 409 A/P ANTI/BAC KITCN|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00044600008882|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.762919|1.4095788500714863|471|1
35.442529|d96f1dc9da02676a60f246c5292beb2fd4696f3a|8.99|2015-03-02 19:30:00|1.4102725052409182|2|7203688113|471|0.6185888262835733|0|1|583|-80.762919|136|35.442529|NUTS|0.0|4|HT PECAN PIECES TRAY|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00072036881137|OTHER MERCHANDISE|PRODUCE|-80.762919|1.4095788500714863|471|1
35.442529|a4fdd7ab83a589e7888c92373928aa03164d7255|3.99|2014-12-16 21:08:00|1.4102725052409182|2|7203671361|471|0.6185888262835733|0|1|317|-80.762919|52|35.442529|CHUNK AND BAR CHEESE|0.3|3|HT TRDR COLBY JCK CRACKER CUTS|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00072036713629|CHEESE|DAIRY|-80.762919|1.4095788500714863|471|1
35.442529|fc08fef3730a7114330cba4d2c81f1da44eff70a|1.67|2014-12-14 14:04:00|1.4102725052409182|2|3120001605|471|0.6185888262835733|0|1|106|-80.762919|16|35.442529|CRANBERRY SAUCE|0.17|1|OS CRANBERRY SC WHOLE|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00031200016034|FRUIT-CAN/JAR|G1 GROCERY|-80.762919|1.4095788500714863|471|1
35.442529|1b07eb66ad1ac00d0b7805dc8234005a019beb8c|8.58|2014-11-04 18:38:00|80.749667378538092|2|2840016014|471|35.462678055660284|0|3|201|-80.860108|31|35.500972|POTATO CHIPS|3.58|1|LAYS CLASSIC|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|35.465179900649026|00028400160148|SNACKS|G1 GROCERY|-80.762919|80.762923050859683|268|2
35.442529|84546e1c1c874f6caede9ff0e3d5817c2afe43f7|2.69|2014-09-26 22:12:00|80.749667378538092|2|7225001739|471|35.462678055618937|0|3|1025|-80.746334|162|35.41832|WHITE|0.0|7|NATOWN WHITEWHEAT RTOP BRD|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|35.465179900649026|00072250017398|SLICED BREAD|COMMERCIAL BAKERY|-80.762919|80.762923349742664|190|1
35.442529|b6484d4e1e50d705e7a5b3fd2d93c6d569d44a1a|2.69|2014-10-19 20:10:00|1.4102725052409182|2|7225001739|471|0.6185888262835733|0|1|1025|-80.762919|162|35.442529|WHITE|0.5|7|NATOWN WHITEWHEAT RTOP BRD|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00072250017398|SLICED BREAD|COMMERCIAL BAKERY|-80.762919|1.4095788500714863|471|1
35.442529|48399cd8cf3d943b5070e3b3585c28ffe2d22c58|3.49|2014-12-18 11:27:00|1.4102725052409182|2|7675325877|471|0.6185888262835733|0|1|6821|-80.762919|1580|35.442529|J HOOK LAMI PROGRAM|0.0|18|"GC 12"" SELF LOCK TONGS S/S"|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00076753258777|J-HOOK|GM|-80.762919|1.4095788500714863|471|1
35.442529|b2a796337cdb4c348fe6d45a58d8ee86da4ddd01|5.98|2014-12-16 21:07:00|1.4102725052409182|2|7199800001|471|0.6185888262835733|0|1|1246|-80.762919|34|35.442529|SPICE BLENDS|0.0|1|TONY CHACHERE CREOLE SEASONG|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00071998000013|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.762919|1.4095788500714863|471|2
35.442529|d45df5ea753382ab746b52ed8ef3e844e9ed82fa|2.69|2014-10-11 21:31:00|1.4102725052409182|2|1113200681|471|0.6185888262835733|0|1|155|-80.762919|24|35.442529|NFS-DOG TREATS|0.0|1|ALPO VARIETY SNAPS|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00011132006815|PET FOOD/SUPPLIES|G1 GROCERY|-80.762919|1.4095788500714863|471|1
35.442529|a5d467929fbb0b61c554d875a979f199a95e8374|11.97|2014-11-23 20:18:00|1.4102725052409182|2|3338324028|471|0.6185888262835733|0|1|504|-80.762919|64|35.442529|FRESH BERRIES|2.32|4|BLACKBERRIES 5.6 OZ|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00881006001099|FRESH PRODUCE|PRODUCE|-80.762919|1.4095788500714863|471|3
35.442529|cac025fa69ce076a66c249df3be233d40c977b59|5.7|2014-09-22 22:30:00|80.749667378538092|2|8390000536|471|35.462678055618937|0|3|365|-80.746334|56|35.41832|REFRIGERATED TEAS|2.1|3|GOLD PEAK DIET TEA|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|35.465179900649026|00083900005382|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.762919|80.762923349742664|190|2
35.442529|9cf2b0dd0faf36c85ee23cf6c02b7cb8284ebb5f|3.34|2015-01-18 14:32:00|1.4102725052409182|2|7203698181|471|0.6185888262835733|0|1|276|-80.762919|45|35.442529|ICE MILK/SHERBET/YOGURT-FROZEN|0.33|5|HT FF VANILLA YOGURT|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00072036981813|ICE CREAM|FROZEN|-80.762919|1.4095788500714863|471|1
35.442529|630ff2933c0ed75998e9a7b3c5c656b63758fc9c|6.99|2014-11-14 18:25:00|1.4102725052409182|2|7203670967|471|0.6185888262835733|0|1|37|-80.762919|10|35.442529|PODS/CUPS/SINGLES|0.6|1|HT HOUSE BLEND DECAF K-CUPS|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00072036709691|COFFEE|G1 GROCERY|-80.762919|1.4095788500714863|471|1
35.442529|3fa36f28b857f4b8ac9ed7a7851bf75e0ca92a19|5.19|2014-10-30 21:15:00|1.4102725052409182|2|89162700903|471|0.6185888262835733|0|1|1278|-80.762919|48|35.442529|SINGLE SERVE NUTRITIONAL|0.0|5|EVOL TANDOORI CHICKEN|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00891627009084|FROZEN MEALS|FROZEN|-80.762919|1.4095788500714863|471|1
35.442529|4137ec8f20ce9d9a6e4845c9bcc9a88af39c858f|1.61|2014-09-30 22:26:00|1.4102725052409182|2||471|0.6185888262835733|0|1|502|-80.762919|64|35.442529|FRESH BANANAS|0.0|4|BANANAS, YELLOW|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.762919|1.4095788500714863|471|1
35.442529|4ac55f38dfcea18dc8f3041b5446f53e8aadbc1e|4.99|2014-10-07 19:40:00|1.4102725052409182|2|7343509330|471|0.6185888262835733|0|1|1613|-80.762919|371|35.442529|THAW & SELL (BREAD)|1.99|14|KING'S HAWAIIAN SLICED BREAD|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00073435093305|BREAD|BAKERY|-80.762919|1.4095788500714863|471|1
35.442529|fa83d214557a4244844cbcf5f51e94509ef1b183|2.79|2014-12-07 20:03:00|1.4102725052409182|2|85392300200|471|0.6185888262835733|0|1|686|-80.762919|61|35.442529|FRUIT ON BOTTOM|0.32|3|NOOSA YOGHURT PINEAPPLE|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00853923002169|YOGURT|DAIRY|-80.762919|1.4095788500714863|471|1
35.442529|6edb697911ac6c792ac717a64582c8754f5b4e16|5.99|2014-09-30 18:55:00|80.749667378538092|2|3160018401|471|35.462678055660284|0|3|5529|-80.860108|1506|35.500972|SHOE CARE-POLISH|0.0|18|KIWI EXPRESS SHINE BLACK|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|35.465179900649026|00031600184012|SHOE CARE/LACES/SEWING|GM|-80.762919|80.762923050859683|268|1
35.442529|9093d6a25748b19adf6251dbe1c7a8552788bf49|14.59|2014-11-27 10:54:00|80.749667378538092|2|30299391716|471|35.462678055618937|0|3|3202|-80.746334|1015|35.41832|HAND & BODY THERAPEUTIC|2.0|17|CETAPHIL MOISTURIZING CREAM|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|35.465179900649026|00302993917168|HAND & BODY LOTION/SUN CARE|HBC|-80.762919|80.762923349742664|190|1
35.442529|44a4c947e82c16dc8617293259e213b7077c9e98|5.99|2014-10-10 13:35:00|80.749667378538092|2|2301200011|471|35.462678054089814|0|3|1475|-80.861571|485|35.444615|SUSHI CLASSIC|0.0|6|VEGETABLE COMBO|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|35.465179900649026|00023012000110|SUSHI|DELI|-80.762919|80.762929572760186|340|1
35.442529|620fab0499d2f8f946326eb8ff3473ec3f7a57f8|3.65|2014-12-06 20:42:00|1.4102725052409182|2|3010067264|471|0.6185888262835733|0|1|91|-80.762919|13|35.442529|SPRAYED BUTTER CRACKERS|1.15|1|TOWN HOUSE FLATBRD SEASALT OLV|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00030100506560|CRACKERS|G1 GROCERY|-80.762919|1.4095788500714863|471|1
35.442529|675df03471293dc7d432ef58ffff9dc8f99e1581|1.99|2014-12-21 13:47:00|1.4102725052409182|2||471|0.6185888262835733|0|1|274|-80.762919|44|35.442529|ICE|0.2|5|HT BAGGED ICE|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00072036480118|ICE|FROZEN|-80.762919|1.4095788500714863|471|1
35.442529|9923f31b10a6e84e622bbc309fab341306b1456d|12.99|2014-12-07 18:50:00|80.749667378538092|2|20577400000|471|35.462678055660284|0|3|1820|-80.860108|410|35.500972|BH BEEF|0.0|6|BH MESQUITE BEEF BRISKET|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|35.465179900649026|00205774000007|BH MEAT|DELI|-80.762919|80.762923050859683|268|1
35.442529|8209ffef31caa789e7dbc59526f986645bee0bf2|7.99|2015-02-04 18:23:00|80.749667378538092|2|2301200207|471|35.462678055660284|0|3|1475|-80.860108|485|35.500972|SUSHI CLASSIC|0.0|6|CRUNCHY SHRIMP ROLL|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|35.465179900649026|00023012002077|SUSHI|DELI|-80.762919|80.762923050859683|268|1
35.442529|fbb641a6c13e839c6e309227a05709a0a8a7dd59|1.29|2014-11-28 18:52:00|1.4102725052409182|2|2200000899|471|0.6185888262835733|0|1|48|-80.762919|7|35.442529|REGISTER GUM|0.0|1|EXTRA POLAR ICE 15 PC|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00022000008985|CANDY|G1 GROCERY|-80.762919|1.4095788500714863|471|1
35.442529|e4b1bbdfc14af1cb58e78e82ee9692e531e0a76e|2.49|2015-02-13 19:20:00|80.749667378538092|2|5100012573|471|35.462678055618937|0|3|137|-80.746334|20|35.41832|TOMATO & VEGETABLE JUICE|0.3|1|V8 SPLASH STRAWBERRY LEMONADE|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|35.465179900649026|00051000212597|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.762919|80.762923349742664|190|1
35.442529|45dfd73be077d58d513a9d5e47b294956d156d45|4.29|2015-01-18 14:10:00|80.749667378538092|2|7343500004|471|35.462678055660284|0|3|1631|-80.860108|373|35.500972|THAW & SELL (ROLLS)|0.0|14|KING'S HAWAIIAN 12CT ROLLS|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|35.465179900649026|00073435000044|ROLLS|BAKERY|-80.762919|80.762923050859683|268|1
35.442529|bfd81cf11244f9e9d7cd88e1f5622462ee750455|4.99|2015-02-22 09:54:00|1.4102725052409182|2|7420003201|471|0.6185888262835733|0|1|6816|-80.762919|1572|35.442529|LADIES/GIRLS SOCKS|0.0|18|(JHK)L'EGGS SLK TGT SZ B 03201|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00074200032017|SOCKS|GM|-80.762919|1.4095788500714863|471|1
35.442529|1c9c2ac3c9bf3644973e3cec0c7d103079e027a4|3.25|2014-10-29 21:05:00|80.749667378538092|2|3120020007|471|35.462678054089814|0|3|130|-80.861571|20|35.444615|CRANBERRY JUICE/DRINKS-SHELF|0.0|1|OSPRAY LIGHTSTYLE CRANBERRY|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|35.465179900649026|00031200342270|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.762919|80.762929572760186|340|1
35.442529|0e3e15c63229111cb5ff672a99fe409efc80cf72|16.7|2015-02-07 20:57:00|1.4102725052409182|2|76211188813|471|0.6185888262835733|0|1|37|-80.762919|10|35.442529|PODS/CUPS/SINGLES|2.72|1|STARBUCKS VERANDA KCUP|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|0.61833652052202714|00762111895318|COFFEE|G1 GROCERY|-80.762919|1.4095788500714863|471|2
35.442529|2204f26b9df563ae97f79f6c3a86250c51ec791f|1.19|2015-01-06 15:15:00|80.749667378538092|2|4178900301|471|35.462678055660284|0|3|1203|-80.860108|33|35.500972|RAMEN|0.19|1|MARUCHAN BOWL HOTSPICY CHICKEN|b3578ac112de48e5e9f3282499f7cf954ea7e3b5|1.3922511065686183|35.465179900649026|00041789003028|SOUP|G1 GROCERY|-80.762919|80.762923050859683|268|1
35.037115|7698ae5d50a793fec7b776e9dca7ba96b0f5c9eb|1.99|2015-02-16 15:39:00|80.805842308733688|1|7680828073|27|35.050796166851271|0|49|149|-80.770346|23|35.052812|WHSE PASTA CORE|0.49|1|BARILLA PASTA ROTINI|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|35.053350220983141|00076808280982|PASTA|G1 GROCERY|-80.8062|80.806205440656484|40|1
35.037115|c8d63a8f3c5c7449fa5bc0109b372309e557aa5e|13.3|2014-10-29 10:44:00|1.4091206135396188|1|7320289451|27|0.611513017149893|0|47|1277|-80.8062|279|35.037115|FROZEN SNACKS|0.0|5|JOSE OLE CHICKEN NACHO BITES|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|0.61242566243833529|00073202895248|FROZEN SANDWICH AND SNACKS|FROZEN|-80.8062|1.4103342460250419|27|2
35.037115|8260ef420f90403035455d13da5f43883865c70f|7.99|2014-12-23 13:36:00|80.805842308733688|1|7203695817|27|35.050796167325586|0|49|1945|-80.816172|465|35.059823|SUPERFLAG CHEF CASE|2.0|6|QUICHE LORRAINE|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|35.053350220983141|00072036958174|COLD PREPARED FOODS|DELI|-80.8062|80.806203199785557|66|1
35.037115|cdc1da681690e9d8351e41816974eaa3ddb759d7|12.14|2014-12-09 12:10:00|1.4091206135396188|1|20253500000|27|0.611513017149893|0|47|299|-80.8062|49|35.037115|ANGUS BEEF|0.0|2|ANGUS BEEF SIRLOIN STIR FRY|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|0.61242566243833529|00202533000001|BEEF|MEAT|-80.8062|1.4103342460250419|27|2
35.037115|bbc7e8da283c225442894ffbb6d8a24435303342|11.83|2014-10-01 16:06:00|80.805842308733688|1|20322700000|27|35.050796167325586|0|49|644|-80.816172|137|35.059823|NATURAL PORK|0.0|2|NIMAN PORK BNLS CENTER LOIN|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|35.053350220983141|00203227000000|PORK|MEAT|-80.8062|80.806203199785557|66|1
35.037115|546c75eab4e5b67adbcff6cdab245df5c91652a8|8.99|2014-11-18 12:00:00|1.4091206135396188|1|8259266064|27|0.611513017149893|0|47|577|-80.8062|136|35.037115|OTHER MERCH FR MSC JUICE|0.0|4|NAKED BLUE MACHINE|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|0.61242566243833529|00082592727640|OTHER MERCHANDISE|PRODUCE|-80.8062|1.4103342460250419|27|1
35.037115|30bfb1f79cabec8f72d30f56ad928c4e95cd018a|3.96|2014-09-12 11:12:00|1.4091206135396188|1|20253500000|27|0.611513017149893|0|47|299|-80.8062|49|35.037115|ANGUS BEEF|0.0|2|ANGUS BEEF SIRLOIN STIR FRY|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|0.61242566243833529|00202533000001|BEEF|MEAT|-80.8062|1.4103342460250419|27|1
35.037115|80cbaa37c7fa763b951d8e3c78ad641641710cad|2.99|2014-11-03 16:45:00|80.805842308733688|1|7127913204|27|35.050796167325586|0|49|555|-80.816172|64|35.059823|PACKAGED SALADS|0.0|4|F.E. FLAT LEAF SPINACH,PKG|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|35.053350220983141|00071279132044|FRESH PRODUCE|PRODUCE|-80.8062|80.806203199785557|66|1
35.037115|58f8ccb2be27b42454461fb142adc6d40c800599|2.5|2014-11-26 15:38:00|80.805842308733688|1|7203603104|27|35.050796166851271|0|49|757|-80.770346|3|35.052812|BAKING NUTS|0.5|1|HT PECAN CHIPS PEG|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|35.053350220983141|00072036031044|BAKING SUPPLIES|G1 GROCERY|-80.8062|80.806205440656484|40|1
35.037115|d5b3b983fec43489832c689f9ef97f695bc2a242|4.19|2015-01-05 16:47:00|1.4091206135396188|1|7203663089|27|0.611513017149893|0|47|345|-80.8062|57|35.037115|ORGANIC MILK|0.0|3|HTO ORGANIC CRTN WHOLE MILK|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|0.61242566243833529|00072036763860|MILK|DAIRY|-80.8062|1.4103342460250419|27|1
35.037115|49ccb39868275df4300039298e4c8b4cca7eedec|3.85|2014-09-20 17:17:00|80.805842308733688|1|7203663089|27|35.050796047737641|0|49|345|-80.893784|57|35.478031|ORGANIC MILK|0.0|3|HTO ORGANIC CRTN WHOLE MILK|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|35.053350220983141|00072036763860|MILK|DAIRY|-80.8062|80.80626994283493|179|1
35.037115|c74cbb293ba2eac9ca5f72c3bc0f4f1e290b2580|5.99|2015-02-11 15:41:00|80.805842308733688|1|7203676366|27|35.050796167325586|0|49|228|-80.816172|36|35.059823|TABLE SYRUP|1.0|1|HTO MAPLE SYRUP|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|35.053350220983141|00072036763662|TABLE SYRUPS|G1 GROCERY|-80.8062|80.806203199785557|66|1
35.037115|a163e73cd0a04860fcb17b3e44c2578ca4432f23|1.39|2014-10-29 16:19:00|80.805842308733688|1|5210094269|27|35.050796167325586|0|49|80|-80.816172|34|35.059823|SEASONING PACKETS|0.83|1|MC MILD CHILI SEASONING MIX|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|35.053350220983141|00052100155203|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.8062|80.806203199785557|66|1
35.037115|ccf80cc6358fb71423fc41a8f0ffb456ca9becd5|3.57|2014-12-04 13:40:00|80.805842308733688|1|7203603100|27|35.050796167325586|0|49|757|-80.816172|3|35.059823|BAKING NUTS|0.0|1|HT WALNUT PIECES|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|35.053350220983141|00072036031006|BAKING SUPPLIES|G1 GROCERY|-80.8062|80.806203199785557|66|1
35.037115|ebefcd1b58b5d525dadc97956864b058a3fc467a|3.99|2014-11-23 16:37:00|1.4091206135396188|1|7203618378|27|0.611513017149893|0|47|887|-80.8062|152|35.037115|SALADS|1.02|12|JALAPENO CRAB QUESO|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|0.61242566243833529|00072036183781|SALADS/DIPS|SEAFOOD|-80.8062|1.4103342460250419|27|1
35.037115|1fbec39569e1c23479f2ee1a7c6bf2c142a3070c|5.99|2014-09-15 15:48:00|80.805842308733688|1|6205881797|27|35.050796167325586|0|49|79|-80.816172|273|35.059823|ASIAN SAUCES/SEASONINGS|0.0|1|SHARWOOD CHUTNEY MANGO GINGER|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|35.053350220983141|00062058817979|ASIAN PREP. FOODS|G1 GROCERY|-80.8062|80.806203199785557|66|1
35.037115|e6d4f2c4f8f2092eb3b1c3fc7dc4f25628190e50|3.19|2015-02-25 10:46:00|1.4091206135396188|1|2460001700|27|0.611513017149893|0|47|221|-80.8062|34|35.037115|SALT SALT SUBSTITUTES|0.0|1|MORTON COARSE KOSHER SALT|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|0.61242566243833529|00024600017008|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.8062|1.4103342460250419|27|1
35.037115|5b927f88202082395b82d8347a9500182d2d64a6|3.59|2014-11-13 14:54:00|1.4091206135396188|1|3377601120|27|0.611513017149893|0|47|313|-80.8062|51|35.037115|MARGARINE|1.8|3|SMART BAL W/OMEGA 3 BTRY SPRD|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|0.61242566243833529|00033776011031|BUTTER & MARGARINE|DAIRY|-80.8062|1.4103342460250419|27|1
35.037115|a3383665b7086bf13895253f5dd1c3a4dbe19b6a|2.99|2014-12-24 17:56:00|1.4091206135396188|1|7203663217|27|0.611513017149893|0|47|330|-80.8062|55|35.037115|EGGS|0.0|3|HT GRADE A LARGE EGGS 18 CT|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|0.61242566243833529|00072036632173|EGGS FRESH|DAIRY|-80.8062|1.4103342460250419|27|1
35.037115|d2d15f707ec528c1431280fa98fccd2693091fef|4.49|2014-09-24 15:50:00|80.805842308733688|1|7027710520|27|35.050796166851271|0|49|2020|-80.770346|505|35.052812|CHEESE SPECIALTIES|0.0|6|ATHENOS FETA TRADITIONAL CRMBD|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|35.053350220983141|00070277105203|SPECIALTY CHEESE|DELI|-80.8062|80.806205440656484|40|1
35.037115|fb0ca1dea6ae6741c57db09018c62eb1e7ab6dcd|1.69|2014-09-22 16:13:00|1.4091206135396188|1|5480005009|27|0.611513017149893|0|47|238|-80.8062|38|35.037115|RICE FLAVORED|0.69|1|UNCLE BENS C INN CHICKEN R/V|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|0.61242566243833529|00054800050093|RICE GRAINS AND BEANS|G1 GROCERY|-80.8062|1.4103342460250419|27|1
35.037115|246c4e6f6bea726e89acf7c485469aefae49e5d9|1.33|2014-10-18 11:07:00|1.4091206135396188|1|89470001004|27|0.611513017149893|0|47|685|-80.8062|61|35.037115|GREEK|0.33|3|CHOBANI SEASONAL GREEN TEA|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|0.61242566243833529|00818290013866|YOGURT|DAIRY|-80.8062|1.4103342460250419|27|1
35.037115|3465979aea5aeba97a7b150e5c6fc208797bbeb9|2.49|2014-10-04 18:28:00|1.4091206135396188|1|7203688048|27|0.611513017149893|0|47|526|-80.8062|64|35.037115|FRESH MUSHROOMS|0.0|4|HT SLICED BABY BELLAS|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|0.61242566243833529|00072036880482|FRESH PRODUCE|PRODUCE|-80.8062|1.4103342460250419|27|1
35.037115|0962141f771250266851122c363cd41dc5c34f26|3.99|2014-10-08 09:29:00|1.4091206135396188|1|7203695283|27|0.611513017149893|0|47|1663|-80.8062|381|35.037115|CREME CAKE|0.0|14|FFM SLICED POUND CAKE|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|0.61242566243833529|00072036952752|CAKES|BAKERY|-80.8062|1.4103342460250419|27|1
35.037115|0012cc902c579cb58a086d0ee6e9a27cbe686b39|3.99|2014-10-31 10:03:00|1.4091206135396188|1|7203695676|27|0.611513017149893|0|47|1656|-80.8062|381|35.037115|CUP CAKES|0.0|14|FFM MINI VANILLA CUPCAKES|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|0.61242566243833529|00072036956767|CAKES|BAKERY|-80.8062|1.4103342460250419|27|1
35.037115|945327768e61d868a4ad18a130c376245c77d708|3.65|2015-02-26 16:09:00|1.4091206135396188|1|7585600110|27|0.611513017149893|0|47|273|-80.8062|43|35.037115|PREMIUM NOVELTIES|0.0|5|KLONDIKE SLIM A BEAR VAN 8CT|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|0.61242566243833529|00075856012422|FROZEN NOVELTIES|FROZEN|-80.8062|1.4103342460250419|27|1
35.037115|31cb25bedc8167895229bd01ca2be5baa585c49e|4.29|2014-11-21 14:56:00|80.805842308733688|1|4400003037|27|35.050796167325586|0|49|90|-80.816172|13|35.059823|SNACK CRACKERS|2.15|1|WHEAT THINS ORIGINAL|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|35.053350220983141|00044000030377|CRACKERS|G1 GROCERY|-80.8062|80.806203199785557|66|1
35.037115|66a140ebd3196aed38a0275e957c4e0a72bfa673|4.59|2015-03-05 13:00:00|80.805842308733688|1|78142152423|27|35.050796167325586|0|49|1601|-80.816172|371|35.059823|BRANDED BREAD|1.15|14|LA BREA SUNFLOWER HONEY LOAF|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|35.053350220983141|00781421524237|BREAD|BAKERY|-80.8062|80.806203199785557|66|1
35.037115|28161cfed121cc5331767c472d33ca82788baf84|4.49|2014-10-03 13:43:00|80.805842308733688|1|71575620002|27|35.050796166851271|0|49|504|-80.770346|64|35.052812|FRESH BERRIES|0.5|4|STRAWBERRIES 1LB CLAM|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|35.053350220983141|00812049005102|FRESH PRODUCE|PRODUCE|-80.8062|80.806205440656484|40|1
35.037115|cc5d63c84acad26cb51721bd7b1172f9711e90ef|4.59|2014-12-30 13:22:00|1.4091206135396188|1|78142152423|27|0.611513017149893|0|47|1601|-80.8062|371|35.037115|BRANDED BREAD|0.0|14|LA BREA SUNFLOWER HONEY LOAF|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|0.61242566243833529|00781421524237|BREAD|BAKERY|-80.8062|1.4103342460250419|27|1
35.037115|75a5f7b6658c65eb4ff9076379409391bb04fa30|4.0|2014-10-09 17:33:00|1.4091206135396188|1|20506500000|27|0.611513017149893|0|47|2020|-80.8062|505|35.037115|CHEESE SPECIALTIES|0.0|6|SPECIALITY CHEESE BY COUNT|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|0.61242566243833529|00205065000006|SPECIALTY CHEESE|DELI|-80.8062|1.4103342460250419|27|1
35.037115|d1563fc02ff6da111a7e5395e03c0d4ad04789eb|8.1|2015-02-20 16:27:00|80.805842308733688|1||27|35.050796166851271|0|49|503|-80.770346|64|35.052812|FRESH GRAPES|1.16|4|RED GRAPES,SEEDLESS 12/16|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|35.053350220983141|00204023000003|FRESH PRODUCE|PRODUCE|-80.8062|80.806205440656484|40|1
35.037115|0c7e8b9a70992a8ad3f247f2a86842b5aed811f4|6.49|2014-10-24 09:24:00|1.4091206135396188|1|7203688056|27|0.611513017149893|0|47|562|-80.8062|64|35.037115|FRESH CUT FRUIT|0.0|4|HT MIXED FRUIT CHUNKS 32OZ|b4d20b1da85bfc3039818ad38fe90a1758be51e1|0.9453356406923101|0.61242566243833529|00072036880567|FRESH PRODUCE|PRODUCE|-80.8062|1.4103342460250419|27|1
35.412407|59ab9d0f0eb8de1c8db7d421f3e13f874e75a241|2.29|2015-02-01 15:48:00|1.4102725052409182|4|7203663996|68|0.6180630982062877|0|1|342|-80.662946|57|35.412407|FRESH MILK|0.82|3|HARRIS TEETER 2%   MILK|b6eb042482e7af7dedd459820abe420f93e4580c|0.7024097339377912|0.61833652052202714|00072036639998|MILK|DAIRY|-80.662946|1.40783399205839|68|1
35.412407|d6d5c98795524d960d22306f96ede02112b996c0|2.0|2015-01-04 20:15:00|1.4102725052409182|4|7203663159|68|0.6180630982062877|0|1|1134|-80.662946|57|35.412407|CARTON MILK|0.0|3|HARRIS TEETER CHOCOLATE MILK|b6eb042482e7af7dedd459820abe420f93e4580c|0.7024097339377912|0.61833652052202714|00072036631596|MILK|DAIRY|-80.662946|1.40783399205839|68|1
35.412407|eb0722228b3f8344ec929dba56acd9201c4d5827|1.06|2015-02-08 18:15:00|1.4102725052409182|4||68|0.6180630982062877|0|1|523|-80.662946|64|35.412407|FRESH POTATOES|0.11|4|COO SWEET POTATOES, BULK|b6eb042482e7af7dedd459820abe420f93e4580c|0.7024097339377912|0.61833652052202714|00204091000004|FRESH PRODUCE|PRODUCE|-80.662946|1.40783399205839|68|1
35.412407|daf5a16faeba57718e6482c119da2d1a28bbff6a|1.81|2014-09-21 17:07:00|1.4102725052409182|4||68|0.6180630982062877|0|1|523|-80.662946|64|35.412407|FRESH POTATOES|0.42|4|COO SWEET POTATOES, BULK|b6eb042482e7af7dedd459820abe420f93e4580c|0.7024097339377912|0.61833652052202714|00204091000004|FRESH PRODUCE|PRODUCE|-80.662946|1.40783399205839|68|1
35.412407|3a8ea29f16e02346551fc0a042e217363bb238ef|3.39|2015-01-25 17:51:00|1.4102725052409182|4|3800031829|68|0.6180630982062877|0|1|74|-80.662946|9|35.412407|RTE CEREAL ALL FAMILY|0.89|1|KELL MIN WH LIL BITES ORIG|b6eb042482e7af7dedd459820abe420f93e4580c|0.7024097339377912|0.61833652052202714|00038000596827|CEREAL|G1 GROCERY|-80.662946|1.40783399205839|68|1
35.412407|867e28e3360d96ffe1761e4da55f5d277b051ea0|1.89|2014-11-24 16:55:00|1.4102725052409182|4|7800023046|68|0.6180630982062877|0|1|55|-80.662946|8|35.412407|REGULAR|0.89|23|CHERRY SUNDROP 2 LTR|b6eb042482e7af7dedd459820abe420f93e4580c|0.7024097339377912|0.61833652052202714|00078000232462|CARBONATED BEVERAGES|BEVERAGE|-80.662946|1.40783399205839|68|1
35.412407|aa9cdff719c4619c5ed07e907759471d860b7bc7|0.69|2015-02-15 19:30:00|1.4102725052409182|4||68|0.6180630982062877|0|1|509|-80.662946|64|35.412407|FRESH CITRUS-REMAINING|0.0|4|LEMONS, MEDIUM|b6eb042482e7af7dedd459820abe420f93e4580c|0.7024097339377912|0.61833652052202714|00204958000000|FRESH PRODUCE|PRODUCE|-80.662946|1.40783399205839|68|1
35.412407|eb6a92a4e8f1bc78617b9e84d3d591243f9d2e07|2.42|2014-10-02 10:02:00|1.4102725052409182|4|20596200000|68|0.6180630982062877|0|1|1821|-80.662946|410|35.412407|BH TURKEY|0.0|6|BOARS HEAD MAPLE HONEY TURKEY|b6eb042482e7af7dedd459820abe420f93e4580c|0.7024097339377912|0.61833652052202714|00205962000000|BH MEAT|DELI|-80.662946|1.40783399205839|68|1
35.412407|908883fbaff2b4a7ca61f2856e7f369411c2f343|3.99|2014-12-18 18:42:00|1.4102725052409182|4|1090000015|68|0.6180630982062877|0|1|440|-80.662946|76|35.412407|NFS-ALUMINUM FOIL|0.99|1|REYNOLDS FOIL 75 FT|b6eb042482e7af7dedd459820abe420f93e4580c|0.7024097339377912|0.61833652052202714|00010900000154|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.662946|1.40783399205839|68|1
35.412407|cf18611a7cc3a3a3ef47d26c2373d263904b64c9|4.0|2015-02-28 17:34:00|1.4102725052409182|4||68|0.6180630982062877|0|1|511|-80.662946|64|35.412407|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|b6eb042482e7af7dedd459820abe420f93e4580c|0.7024097339377912|0.61833652052202714|00204770000004|FRESH PRODUCE|PRODUCE|-80.662946|1.40783399205839|68|2
35.412407|7ce75ecaf1f9703677e758ce472df9923731157f|2.99|2014-12-10 17:23:00|1.4102725052409182|4|7203698770|68|0.6180630982062877|0|1|176|-80.662946|72|35.412407|NFS-DISPOSE CUPS|0.99|1|YH CLEAR CUPS 9 OZ|b6eb042482e7af7dedd459820abe420f93e4580c|0.7024097339377912|0.61833652052202714|00072036987709|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.662946|1.40783399205839|68|1
35.412407|09ca0241e916da9200cd5cd1255a45097f433ae3|0.7|2015-02-16 12:22:00|80.66957994482128|4|7203625010|68|35.422572467162134|0|38|145|-80.764523|22|35.341927|MILK-CANNED|0.0|1|HT  EVAPORATED MILK|b6eb042482e7af7dedd459820abe420f93e4580c|0.7024097339377912|35.385064306269825|00072036250100|PACKAGED MILKS & MODIFIERS|G1 GROCERY|-80.662946|80.662960909514112|220|1
35.412407|8d5d18c5c6bef47136f9afa9a23e0e2d5a4177cd|1.77|2015-01-24 18:34:00|1.4102725052409182|4|7203657031|68|0.6180630982062877|0|1|322|-80.662946|53|35.412407|SOUR CREAM|0.5|3|HT SOUR CREAM|b6eb042482e7af7dedd459820abe420f93e4580c|0.7024097339377912|0.61833652052202714|00072036570314|CULTURES|DAIRY|-80.662946|1.40783399205839|68|1
35.412407|e6f302fb1321bfde414ecac27e5bb3cdfb2a6732|3.98|2014-12-23 22:32:00|1.4102725052409182|4|7127915101|68|0.6180630982062877|0|1|555|-80.662946|64|35.412407|PACKAGED SALADS|0.0|4|F.E. SHREDS|b6eb042482e7af7dedd459820abe420f93e4580c|0.7024097339377912|0.61833652052202714|00071279151014|FRESH PRODUCE|PRODUCE|-80.662946|1.40783399205839|68|2
35.412407|3a9fc78faf702254154f263103da59f1203a3118|0.95|2015-01-10 21:57:00|1.4102725052409182|4|4600028869|68|0.6180630982062877|0|1|77|-80.662946|272|35.412407|HISP SAUCES/SEASONINGS|0.2|1|E  OEP SEASONING TACO|b6eb042482e7af7dedd459820abe420f93e4580c|0.7024097339377912|0.61833652052202714|00046000288697|HISPANIC PREP. FOODS|G1 GROCERY|-80.662946|1.40783399205839|68|1
35.412407|542060d84937503854d70165bb7fea7f1146a76a|0.7|2015-01-11 21:07:00|1.4102725052409182|4|20543600000|68|0.6180630982062877|0|1|1832|-80.662946|415|35.412407|BH SLICING CHEESE|0.0|6|BOARS HEAD MONTEREY JACK CHSE|b6eb042482e7af7dedd459820abe420f93e4580c|0.7024097339377912|0.61833652052202714|00205436000000|SLICING CHEESE|DELI|-80.662946|1.40783399205839|68|1
35.412407|6e2d2103fa63aacb3cff5d5605ecc59fa842a973|1.79|2014-11-18 20:56:00|1.4102725052409182|4|7203663157|68|0.6180630982062877|0|1|1134|-80.662946|57|35.412407|CARTON MILK|0.0|3|HARRIS TEETER 2% MILK|b6eb042482e7af7dedd459820abe420f93e4580c|0.7024097339377912|0.61833652052202714|00072036631558|MILK|DAIRY|-80.662946|1.40783399205839|68|1
35.412407|bad99435276570127c44941598bd4ee73da3eb11|1.99|2014-10-05 13:53:00|1.4102725052409182|4|7203663120|68|0.6180630982062877|0|1|495|-80.662946|108|35.412407|NON REFRIGERATED|1.0|19|"HT 8"" BURRITO TORTILLA"|b6eb042482e7af7dedd459820abe420f93e4580c|0.7024097339377912|0.61833652052202714|00072036631206|TORTILLAS|CASE READY MEATS|-80.662946|1.40783399205839|68|1
35.412407|c98db259871640016aeb73028ef2685a8b6a6c91|2.19|2015-02-16 15:54:00|1.4102725052409182|4|1200000230|68|0.6180630982062877|0|1|55|-80.662946|8|35.412407|REGULAR|0.69|23|PEPSI COLA 2 LTR NR|b6eb042482e7af7dedd459820abe420f93e4580c|0.7024097339377912|0.61833652052202714|00012000002304|CARBONATED BEVERAGES|BEVERAGE|-80.662946|1.40783399205839|68|1
35.412407|54d0e45cd994964ac6ab13d2f321e7d2c20e48df|1.59|2014-09-18 17:33:00|1.4102725052409182|4|1600043054|68|0.6180630982062877|0|1|10|-80.662946|2|35.412407|LAYER CAKE MIX|0.0|1|BC SUPER MOIST DEVILS FOOD|b6eb042482e7af7dedd459820abe420f93e4580c|0.7024097339377912|0.61833652052202714|00016000409828|BAKING MIXES|G1 GROCERY|-80.662946|1.40783399205839|68|1
35.412407|7f53d6da089948b649686d2cad9cca1a29529d69|6.02|2015-01-18 15:00:00|1.4102725052409182|4|20897500000|68|0.6180630982062877|0|1|977|-80.662946|201|35.412407|FRESH HT CHICKEN|3.02|2|FRESH BONELESS CHICKEN BREAST|b6eb042482e7af7dedd459820abe420f93e4580c|0.7024097339377912|0.61833652052202714|00208975000005|POULTRY|MEAT|-80.662946|1.40783399205839|68|1
35.412407|7dce5c3f6cdf320360eca42d9fa1801bab20afe5|1.35|2015-02-22 18:22:00|1.4102725052409182|4|20543700000|68|0.6180630982062877|0|1|1832|-80.662946|415|35.412407|BH SLICING CHEESE|0.0|6|BOARS HEAD PEPPER JACK CHEESE|b6eb042482e7af7dedd459820abe420f93e4580c|0.7024097339377912|0.61833652052202714|00205437000009|SLICING CHEESE|DELI|-80.662946|1.40783399205839|68|1
35.412407|ea8e1d2d9d67ab26f411d697f3046787dfdcc11b|4.59|2014-10-16 17:44:00|1.4102725052409182|4|20897500000|68|0.6180630982062877|0|1|977|-80.662946|201|35.412407|FRESH HT CHICKEN|2.3|2|FRESH BONELESS CHICKEN BREAST|b6eb042482e7af7dedd459820abe420f93e4580c|0.7024097339377912|0.61833652052202714|00208975000005|POULTRY|MEAT|-80.662946|1.40783399205839|68|1
35.444615|3419de1652c44a61f6913d5c75c7f3473378addb|5.5|2015-01-07 16:29:00|80.86161257435397|1|20596200000|340|35.471245480410708|0|36|1821|-80.844274|410|35.204336|BH TURKEY|0.0|6|BOARS HEAD MAPLE HONEY TURKEY|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00205962000000|BH MEAT|DELI|-80.861571|80.861650033664503|61|1
35.444615|0b73992be8c88f3dd823fea30fc00922df027973|16.36|2014-11-16 13:53:00|80.86161257435397|1||340|35.471245480410708|0|36|562|-80.844274|64|35.204336|FRESH CUT FRUIT|0.0|4|MIXED FRUIT (IN-STORE)|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00204472000005|FRESH PRODUCE|PRODUCE|-80.861571|80.861650033664503|61|3
35.444615|93274a402d6efa06fee2e2f3ca73ef332cfd5715|5.5|2015-02-15 14:57:00|1.4102725052409182|1|20596200000|340|0.6186252338517699|0|1|1821|-80.861571|410|35.444615|BH TURKEY|1.0|6|BOARS HEAD MAPLE HONEY TURKEY|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|0.61833652052202714|00205962000000|BH MEAT|DELI|-80.861571|1.4113006522851637|340|1
35.444615|8502512fd8ad2233eac96939a6fee6517f85528e|3.99|2014-12-24 17:20:00|80.86161257435397|1|7203602701|340|35.471245480410708|0|36|1878|-80.844274|435|35.204336|HUMMUS|0.5|6|FFM ARTISAN RED PEPPER HUMMUS|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00072036027030|SALADS|DELI|-80.861571|80.861650033664503|61|1
35.444615|857abc9cd66ce315ba9d4943ca2658cde1d12487|3.99|2014-12-03 16:37:00|80.86161257435397|1|7203602701|340|35.471245480410708|0|36|1878|-80.844274|435|35.204336|HUMMUS|0.5|6|FFM ARTISAN RED PEPPER HUMMUS|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00072036027030|SALADS|DELI|-80.861571|80.861650033664503|61|1
35.444615|56c5a2211e8098f060b55ae9756601138086d6c4|6.29|2014-10-25 12:00:00|80.86161257435397|1|5113193681|340|35.471245480410708|0|36|729|-80.844274|69|35.204336|NFS-SCOUR PAD/STEEL WOOL|0.0|1|SCOTCH BRITE HEAVY DUTY SCB SP|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00051131936812|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.861571|80.861650033664503|61|1
35.444615|0af54b22fdf4fbf0d78208316b698b25447e514b|3.69|2014-09-10 21:39:00|1.4102725052409182|1|74447391204|340|0.6186252338517699|0|1|1266|-80.861571|57|35.444615|COCONUT MILK|0.0|3|SO DELICIOUS COCONUT UNSWEETEN|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|0.61833652052202714|00744473912056|MILK|DAIRY|-80.861571|1.4113006522851637|340|1
35.444615|a5e4d7fe40451aa5ebdfb9d839f600037d7d275c|17.89|2015-01-27 21:08:00|1.4102725052409182|1|82927450229|340|0.6186252338517699|0|1|152|-80.861571|24|35.444615|NFS-CAT FOOD DRY|3.9|1|MEOW MIX|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|0.61833652052202714|00829274502252|PET FOOD/SUPPLIES|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.444615|fe5b59494330e63c756ddd983e8a1dbf32e85715|3.79|2015-01-13 16:12:00|80.86161257435397|1|7127930100|340|35.471245555788776|0|36|555|-80.762919|64|35.442529|PACKAGED SALADS|0.0|4|F.E. CAESAR SALAD|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00071279301006|FRESH PRODUCE|PRODUCE|-80.861571|80.861584975270006|471|1
35.444615|12df55c29c5078074976fc5cf7b91a8c5b5c8753|6.99|2015-02-22 15:00:00|1.4102725052409182|1|7203602601|340|0.6186252338517699|0|1|1981|-80.861571|480|35.444615|CHIPS|0.0|6|HTT 18 OZ  PITA CHIPS|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|0.61833652052202714|00072036026019|DRY GOODS|DELI|-80.861571|1.4113006522851637|340|1
35.444615|1cb820fe46d9a0078cb295b7c02b41ca47d7bf0d|5.29|2014-10-20 14:41:00|80.86161257435397|1|5385200100|340|35.471245480410708|0|36|1211|-80.844274|272|35.204336|HISP SALSA/DIPS|1.3|1|GREEN MTN GR SALSA MED|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00053852004009|HISPANIC PREP. FOODS|G1 GROCERY|-80.861571|80.861650033664503|61|1
35.444615|c37ce7463dd676819d10fb951b88c8b8e466a450|4.49|2015-01-09 17:07:00|80.86161257435397|1|7203695206|340|35.471245555788776|0|36|1885|-80.762919|440|35.442529|PASTA SAUCE|0.0|6|ALFREDO SAUCE|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00072036952318|PASTA|DELI|-80.861571|80.861584975270006|471|1
35.444615|ae670cfc602113d06c1451b9ce90d263f1de48f7|4.19|2015-02-10 19:14:00|80.86161257435397|1|65638535600|340|35.471245474749971|0|36|1245|-80.80146|34|35.17739|SINGLE SPICES|0.0|1|D&A SPICE MILL ORG GARLIC|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00656385366004|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.861571|80.861652858036848|208|1
35.444615|f0a864367cea4979958c36b75e049b8ec082e216|4.49|2014-09-28 16:22:00|1.4102725052409182|1|74759930652|340|0.6186252338517699|0|1|62|-80.861571|7|35.444615|SPECIALTY BAR/BOX CHOCOLATE|0.5|1|GHIRARDELLI SEASALT SOIREE|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|0.61833652052202714|00747599313059|CANDY|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.444615|790bba0879496f3efe738dec593df553005a6044|2.52|2014-09-15 16:29:00|1.4102725052409182|1||340|0.6186252338517699|0|1|561|-80.861571|64|35.444615|FR PROD ORGANIC PRODUCE|0.0|4|COO ORG MEDJOOL DATES|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|0.61833652052202714|00204862000004|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|f6b3ba5a372c9e0d5904c3cf52959d14ec44de8b|8.69|2014-10-12 15:50:00|1.4102725052409182|1|7203653118|340|0.6186252338517699|0|1|1243|-80.861571|21|35.444615|MIXED NUTS CASHEWS|2.7|1|HT CASHEWS HALVES|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|0.61833652052202714|00072036531186|NUTS|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.444615|cc58cc8c152d471254fd0c6c740d7bc0328621ab|7.78|2015-01-22 19:47:00|1.4102725052409182|1|4610000012|340|0.6186252338517699|0|1|318|-80.861571|52|35.444615|SHREDDED/GRATED CHEESE|2.78|3|SARGENTO OTB 4 CHSE MEX FINE C|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|0.61833652052202714|00046100000922|CHEESE|DAIRY|-80.861571|1.4113006522851637|340|2
35.444615|66edf9de64ac4f44a282a52b795040edf8531318|5.38|2015-02-21 15:43:00|80.86161257435397|1|7008506010|340|35.471245474749971|0|36|1277|-80.80146|279|35.17739|FROZEN SNACKS|1.38|5|BAGEL BITES CHEESE & PEPP|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00070085060121|FROZEN SANDWICH AND SNACKS|FROZEN|-80.861571|80.861652858036848|208|2
35.444615|f8a4937daf44ede2a91d37beeec075f6ab3e1a4b|4.99|2015-01-05 22:18:00|1.4102725052409182|1|71575620002|340|0.6186252338517699|0|1|504|-80.861571|64|35.444615|FRESH BERRIES|0.2|4|STRAWBERRIES 1LB CLAM|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|0.61833652052202714|00769197404021|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|e1fc41a4c2e31dde4ad94b3b4d04d6fbd2f189c9|8.99|2015-02-19 18:53:00|80.86161257435397|1|89953900024|340|35.471245480410708|0|36|458|-80.844274|82|35.204336|CRAFT BEER|0.0|16|TERRAPIN HOPSECUTIONER 6PK|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00899539000243|DOMESTIC BEER|BEER|-80.861571|80.861650033664503|61|1
35.444615|df8c5c78ac5d8a6c0105852b7b5cedad00a846fe|4.99|2014-10-08 21:58:00|1.4102725052409182|1|7940006835|340|0.6186252338517699|0|1|3814|-80.861571|1070|35.444615|INVISIBLE-FEMALE|0.0|17|DOVE GO FRESH RESTORE|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|0.61833652052202714|00079400271778|DEODORANT|HBC|-80.861571|1.4113006522851637|340|1
35.444615|aa9324da986e3f18e9fd5153b28d7c503b6a093d|1.99|2015-01-18 13:36:00|80.86161257435397|1|7348450151|340|35.471245458247765|0|36|100|-80.85013|15|35.175855|CORN MEAL|0.0|1|HSE-AUTRY YELLOW S/R CORNMEAL|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00073484503015|FLOUR|G1 GROCERY|-80.861571|80.861660584923655|218|1
35.444615|599a65219ed923a36aae5be755f26881d612726e|8.98|2014-12-13 12:28:00|80.86161257435397|1|2840009237|340|35.471245458247765|0|36|1981|-80.85013|480|35.175855|CHIPS|0.0|6|STACYS GARLIC BAGEL CHIPS|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00028400092531|DRY GOODS|DELI|-80.861571|80.861660584923655|218|2
35.444615|e6c4d121d4807cb396724747348896f94e11e8f2|1.29|2014-10-27 11:46:00|80.86161257435397|1|8379152001|340|35.471245557378879|0|36|1981|-80.746334|480|35.41832|CHIPS|0.0|6|DIRTY POTATO CHIP BBQ|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00083791520049|DRY GOODS|DELI|-80.861571|80.861579225699984|190|1
35.444615|1fe3844926e4728550924befbd45366e5af0fae2|3.99|2014-10-29 16:59:00|1.4102725052409182|1|4000015140|340|0.6186252338517699|0|1|46|-80.861571|7|35.444615|PKG CHOC|0.99|1|SNICKERS FUN SIZE|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|0.61833652052202714|00040000151401|CANDY|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.444615|d605eeaf76216c359e7e9243959d319b48025669|1.39|2014-09-26 03:32:00|1.4102725052409182|1|4133103857|340|0.6186252338517699|0|1|1214|-80.861571|272|35.444615|AUTHENTIC HISPANIC|0.0|1|GOYA SC RED HOT|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|0.61833652052202714|00041331038577|HISPANIC PREP. FOODS|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.444615|03ed417242f8b78f14b7f0bae8605ddda031c226|3.49|2014-12-05 17:45:00|80.86161257435397|1|1410007712|340|35.471245480410708|0|36|1253|-80.844274|12|35.204336|ALL OTHER COOKIES|0.0|1|PF DESRT SHOP CHOCOLAT BROWNIE|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00014100042181|COOKIES|G1 GROCERY|-80.861571|80.861650033664503|61|1
35.444615|81782ae4817e0eef28d9f8f0f53498938d818749|3.99|2014-12-23 17:16:00|80.86161257435397|1|20980000000|340|35.471245480410708|0|36|1677|-80.844274|383|35.204336|INDIVIDUALS (PASTRY CASE)|0.0|14|CHOCOLATE MOUSSE|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00209804000005|PASTRY CASE|BAKERY|-80.861571|80.861650033664503|61|1
35.444615|5a83c47ae4f9037f493bd87fd38c0339c3eed9e6|2.29|2015-02-17 16:29:00|1.4102725052409182|1|7203695739|340|0.6186252338517699|0|1|1976|-80.861571|475|35.444615|COLD PIZZA OTHER|0.0|6|WHEAT PIZZA DOUGH BALLS|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|0.61833652052202714|00072036957405|PIZZA|DELI|-80.861571|1.4113006522851637|340|1
35.444615|6355af95ed6ef9c4cc7f84186521553d0aa25490|3.99|2015-02-27 18:25:00|80.86161257435397|1|7203695676|340|35.47124555768859|0|36|1656|-80.893784|381|35.478031|CUP CAKES|0.0|14|FFM MINI VANILLA CUPCAKES|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00072036956767|CAKES|BAKERY|-80.861571|80.861577542180754|179|1
35.444615|600cf7f747538cc5f352d881adac26536f46bc9d|4.99|2015-01-14 15:55:00|80.86161257435397|1|4082201114|340|35.471245480410708|0|36|1878|-80.844274|435|35.204336|HUMMUS|2.49|6|HUMMUS W/ ROASTED PINE NUTS|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00040822011747|SALADS|DELI|-80.861571|80.861650033664503|61|1
35.444615|320996bea390ee58f84231b4feaf3060dd5bf829|4.98|2015-02-18 16:44:00|80.86161257435397|1|7478063991|340|35.471245474749971|0|36|30|-80.80146|4|35.17739|CARBONATED WATER|0.49|1|PERRIER 1LT PET CITRON|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00074780643184|BOTTLED WATER|G1 GROCERY|-80.861571|80.861652858036848|208|2
35.444615|5d242fc547c15c71aad797d54fd63d467f3c8d7e|4.49|2014-12-10 18:25:00|1.4102725052409182|1|7203695649|340|0.6186252338517699|0|1|1699|-80.861571|387|35.444615|EVERYDAY (COOKIES)|0.0|14|HT PINK SOFT SUGAR COOKIES|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|0.61833652052202714|00072036956491|COOKIES|BAKERY|-80.861571|1.4113006522851637|340|1
35.444615|3dfd5410e62fc77981906ffdd675057d3f4ca168|4.99|2015-02-09 07:43:00|80.86161257435397|1|8265750406|340|35.471245474749971|0|36|31|-80.80146|4|35.17739|NON CARBONATED WATER|0.5|1|(U)DEER PARK WATER 24PK .5LT|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00082657504063|BOTTLED WATER|G1 GROCERY|-80.861571|80.861652858036848|208|1
35.444615|1df666c0f4b27136c092cdf6054d8847afcda8e2|3.49|2015-02-12 14:34:00|80.86161257435397|1|7146426040|340|35.471245480410708|0|36|577|-80.844274|136|35.204336|OTHER MERCH FR MSC JUICE|0.0|4|BOLTHOUSE PROTEIN PLUS COFFEE|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00071464016272|OTHER MERCHANDISE|PRODUCE|-80.861571|80.861650033664503|61|1
35.444615|3557f555ea240468fc2f86eb0dda9ce028f1a35a|9.98|2015-02-14 16:33:00|80.86161257435397|1|71575620002|340|35.471245474749971|0|36|504|-80.80146|64|35.17739|FRESH BERRIES|2.5|4|STRAWBERRIES 1LB CLAM|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00812049005102|FRESH PRODUCE|PRODUCE|-80.861571|80.861652858036848|208|2
35.444615|fa45ca0010baf115248e765603f99829895a1401|10.99|2014-09-25 20:17:00|80.86161257435397|1|8143406815|340|35.471245480410708|0|36|9957|-80.844274|886|35.204336|NFS-PREM-OTHER RED|0.0|13|RED GUITAR TEMRANILLO|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00081434068156|PREMIUM ($8-$10.99)|WINE|-80.861571|80.861650033664503|61|1
35.444615|3f62a539e5de19c3ce386a275cc008ab6f3f9513|17.490000000000002|2014-12-26 17:42:00|1.4102725052409182|1|27082900000|340|0.6186252338517699|0|1|973|-80.861571|201|35.444615|FRESH PERDUE CHICKEN|0.0|2|PERDUE BNLS CHICKEN BREAST|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|0.61833652052202714|00270829000004|POULTRY|MEAT|-80.861571|1.4113006522851637|340|2
35.444615|e668482783f5e3a9533c86109539510caa0e02ce|5.98|2015-02-26 15:04:00|1.4102725052409182|1|70601011292|340|0.6186252338517699|0|1|1219|-80.861571|275|35.444615|PASTA SC CORE|0.0|1|BARILLA SC TOM BASIL|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|0.61833652052202714|00706010112961|PASTA SAUCES|G1 GROCERY|-80.861571|1.4113006522851637|340|2
35.444615|784c492c24cb403d4ff56610833b26bb4c8e566d|6.99|2015-03-03 18:44:00|80.86161257435397|1|5000025117|340|35.471245532119084|0|36|341|-80.875654|57|35.585842|CREAMERS|0.81|3|COFFEE-MATE ITAL SWT CREAM LIQ|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00050000605354|MILK|DAIRY|-80.861571|80.861616775612248|99|1
35.444615|1b33815d6310234b318ae770ebdc54734a6c848b|2.29|2014-11-04 13:24:00|80.86161257435397|1|4133533217|340|35.471245392949903|0|36|184|-80.771677|28|35.066546|SALAD DRESSINGS-LIQUID|0.0|1|KENS DRS VIN ITALIAN ASIAGO|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00041335000273|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.861571|80.861686183584979|45|1
35.444615|a0e55fbb5e75c066d54d98b8521b8e85a0fa4051|12.99|2015-02-11 10:07:00|80.86161257435397|1|20310500000|340|35.471245480410708|0|36|1153|-80.844274|87|35.204336|NFS-FRESH CUT ARRANGE|0.0|9|*BUDVASE|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00203105000009|FLORAL|FLORAL|-80.861571|80.861650033664503|61|1
35.444615|06e3596d78c9b3b194ddb7711666f4994869ee1a|1.39|2014-12-29 14:07:00|80.86161257435397|1|8265750067|340|35.471245405230086|0|36|31|-80.85753|4|35.116638|NON CARBONATED WATER|0.39|1|DEER PARK WATER 1LT|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00082657500676|BOTTLED WATER|G1 GROCERY|-80.861571|80.861681821772635|204|1
35.444615|fbbea24296dce5da225c8439d1d8e8948c3ba3c2|5.98|2014-12-13 11:02:00|80.86161257435397|1|1111038388|340|35.471245458247765|0|36|6752|-80.85013|1564|35.175855|STAPLER|0.0|18|OW MINI STAPLER W/ STAPLES|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00011110383884|SCHOOL & OFFICE SUPPLY|GM|-80.861571|80.861660584923655|218|2
35.444615|90aaa691608512429f85d450bb2249bf3a4bb9af|1.69|2015-02-12 18:50:00|80.86161257435397|1|4900000044|340|35.471245474749971|0|36|55|-80.80146|8|35.17739|REGULAR|0.0|23|CB SPRITE PROPRIETARY 20 OZ|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00049000007640|CARBONATED BEVERAGES|BEVERAGE|-80.861571|80.861652858036848|208|1
35.444615|5c4329f987eedf6fcb9eaf96abfcbecc46a9870b|0.99|2015-02-10 14:00:00|80.86161257435397|1|7203695306|340|35.471245405230086|0|36|1895|-80.85753|450|35.116638|TEA|0.0|6|FFM GREEN TEA W/GINSENG & HONY|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00072036018908|BEVERAGES|DELI|-80.861571|80.861681821772635|204|1
35.444615|9fd74399700a35cf80deae011402a113fea7666a|1.94|2014-10-30 16:32:00|80.86161257435397|1|7203698758|340|35.471245447440438|0|36|31|-80.849471|4|35.161696|NON CARBONATED WATER|0.0|1|HT SPRING WATER|bb80191f034cd42ef241adf70901f397e0fb0d93|1.8401072626272876|35.472272108304431|00072036987587|BOTTLED WATER|G1 GROCERY|-80.861571|80.861665302809385|35|2
34.977331|a58d7fceab65ead2e02643a55c676e3034f07f9c|2.89|2014-10-01 17:09:00|1.41290891556208|4|1800052180|149|0.6104695895098807|0|33|325|-81.027334|54|34.977331|BISCUITS-REFRIGERATED|0.0|3|PILLSBURY BUTTERMILK BISC 4PK|bea1aab0a475ba6742f2c1e34750b6ef8ee8efda|1.5463774458749717|0.61055446569467375|00018000521807|DOUGH PRODUCTS|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|ea3167dbc16c248d1afbabbb8f6e8c3914a86b6c|8.58|2014-11-16 19:24:00|1.41290891556208|4|2840006399|149|0.6104695895098807|0|33|204|-81.027334|31|34.977331|TORTILLA CHIPS|0.29|1|TOSTITOS HINT OF LIME|bea1aab0a475ba6742f2c1e34750b6ef8ee8efda|1.5463774458749717|0.61055446569467375|00028400064040|SNACKS|G1 GROCERY|-81.027334|1.4141937624131469|149|2
34.977331|74f3d4030ebf9dfe3d894834dd1b1f16a2ef341e|3.19|2014-10-14 17:10:00|1.41290891556208|4|7203632016|149|0.6104695895098807|0|33|195|-81.027334|30|34.977331|SALAD & COOKING OIL|0.69|1|HT VEGETABLE OIL|bea1aab0a475ba6742f2c1e34750b6ef8ee8efda|1.5463774458749717|0.61055446569467375|00072036320223|SHORTENING/OIL|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|6efe5e1cc5a4626f9091abfdb72fd416ff78781f|6.1|2014-12-16 19:44:00|1.41290891556208|4||149|0.6104695895098807|0|33|500|-81.027334|64|34.977331|FRESH APPLES|0.0|4|HONEY CRISP APPLE|bea1aab0a475ba6742f2c1e34750b6ef8ee8efda|1.5463774458749717|0.61055446569467375|00233283000003|FRESH PRODUCE|PRODUCE|-81.027334|1.4141937624131469|149|1
34.977331|ee1b579b131dff194bf9e8195b83bb60d2b71a77|8.98|2014-09-19 18:56:00|1.41290891556208|4|2840009217|149|0.6104695895098807|0|33|1981|-81.027334|480|34.977331|CHIPS|4.49|6|STACY'S PITA CHIPS NAKED|bea1aab0a475ba6742f2c1e34750b6ef8ee8efda|1.5463774458749717|0.61055446569467375|00028400092173|DRY GOODS|DELI|-81.027334|1.4141937624131469|149|2
34.977331|d6aef68379edb2372293f5988fe9b473c925e89d|2.67|2014-09-28 17:18:00|1.41290891556208|4|7203698754|149|0.6104695895098807|0|33|1265|-81.027334|57|34.977331|ALMOND MILK|0.0|3|HT ALMOND DRINK VANILLA|bea1aab0a475ba6742f2c1e34750b6ef8ee8efda|1.5463774458749717|0.61055446569467375|00072036987556|MILK|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|5330814fea57c7910a02103ebc66f786ba985753|2.69|2015-01-04 18:23:00|1.41290891556208|4|7008506010|149|0.6104695895098807|0|33|1277|-81.027334|279|34.977331|FROZEN SNACKS|0.0|5|BAGEL BITES CHEESE & PEPP|bea1aab0a475ba6742f2c1e34750b6ef8ee8efda|1.5463774458749717|0.61055446569467375|00070085060121|FROZEN SANDWICH AND SNACKS|FROZEN|-81.027334|1.4141937624131469|149|1
34.977331|574fee9bef560876ea81312ad0d5e5d525cbd367|2.45|2014-12-14 17:54:00|1.41290891556208|4|1450000253|149|0.6104695895098807|0|33|1272|-81.027334|50|34.977331|BAG VEG STEAM|0.45|5|BE STMFRESH BABY BROCCOLI BLND|bea1aab0a475ba6742f2c1e34750b6ef8ee8efda|1.5463774458749717|0.61055446569467375|00014500012951|VEGETABLES-FROZEN|FROZEN|-81.027334|1.4141937624131469|149|1
34.977331|b70831629d8cc6ab83919d2bb3be380b6ddca3af|1.89|2014-11-24 21:07:00|1.41290891556208|4||149|0.6104695895098807|0|33|500|-81.027334|64|34.977331|FRESH APPLES|0.0|4|RED DEL APPLE, WA  48|bea1aab0a475ba6742f2c1e34750b6ef8ee8efda|1.5463774458749717|0.61055446569467375|00233284000002|FRESH PRODUCE|PRODUCE|-81.027334|1.4141937624131469|149|1
34.977331|76e2b34a147b9cba71cf412647c05aab8e9e52f9|3.38|2015-01-31 10:09:00|1.41290891556208|4|7203688003|149|0.6104695895098807|0|33|527|-81.027334|64|34.977331|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|bea1aab0a475ba6742f2c1e34750b6ef8ee8efda|1.5463774458749717|0.61055446569467375|00072036880031|FRESH PRODUCE|PRODUCE|-81.027334|1.4141937624131469|149|2
34.977331|3d6b0c8f947536d6cad565c6fd566b7ddba5b8e9|4.49|2014-09-18 15:41:00|1.41290891556208|4|7203695906|149|0.6104695895098807|0|33|1609|-81.027334|371|34.977331|TAKE & BAKE BREAD|0.0|14|FFM GARLIC TEAR & SHARE BREAD|bea1aab0a475ba6742f2c1e34750b6ef8ee8efda|1.5463774458749717|0.61055446569467375|00072036959065|BREAD|BAKERY|-81.027334|1.4141937624131469|149|1
34.977331|51b98d2bbde371dc4ad3c52e1166f2a8475b3dbf|2.19|2015-03-08 13:05:00|1.41290891556208|4|4900005010|149|0.6104695895098807|0|33|54|-81.027334|8|34.977331|DIET|0.2|23|DT CLASSIC 2 LITER|bea1aab0a475ba6742f2c1e34750b6ef8ee8efda|1.5463774458749717|0.61055446569467375|00049000050110|CARBONATED BEVERAGES|BEVERAGE|-81.027334|1.4141937624131469|149|1
34.977331|1cebe2b40b334a071f0026fc6c37b261c846a9f0|5.79|2014-10-28 18:38:00|1.41290891556208|4|3680036733|149|0.6104695895098807|0|33|4236|-81.027334|1200|34.977331|DEX ADULT/CHILDREN|0.0|17|TC DAYTIME CLD/FLU PE SOFTGELS|bea1aab0a475ba6742f2c1e34750b6ef8ee8efda|1.5463774458749717|0.61055446569467375|00036800367333|COUGH/COLD/SINUS|HBC|-81.027334|1.4141937624131469|149|1
34.977331|11fb0628086821546c46a39ce5dd079f75e4b9d2|3.49|2014-12-24 18:58:00|1.41290891556208|4|7433610102|149|0.6104695895098807|0|33|342|-81.027334|57|34.977331|FRESH MILK|0.0|3|HIGHLAND CREST SKIM MILK|bea1aab0a475ba6742f2c1e34750b6ef8ee8efda|1.5463774458749717|0.61055446569467375|00074336101083|MILK|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|bbd36ecf477866423edcb965cd8ed3c119fd3a74|27.73|2014-09-29 15:34:00|1.41290891556208|4|20897500000|149|0.6104695895098807|0|33|977|-81.027334|201|34.977331|FRESH HT CHICKEN|13.9|2|FRESH BONELESS CHICKEN BREAST|bea1aab0a475ba6742f2c1e34750b6ef8ee8efda|1.5463774458749717|0.61055446569467375|00208975000005|POULTRY|MEAT|-81.027334|1.4141937624131469|149|1
34.977331|ca1c5898e3df4e211f9464d0f0a0f4b76a16384d|9.82|2014-09-17 16:43:00|1.41290891556208|4|20897500000|149|0.6104695895098807|0|33|977|-81.027334|201|34.977331|FRESH HT CHICKEN|4.92|2|FRESH BONELESS CHICKEN BREAST|bea1aab0a475ba6742f2c1e34750b6ef8ee8efda|1.5463774458749717|0.61055446569467375|00208975000005|POULTRY|MEAT|-81.027334|1.4141937624131469|149|1
34.977331|ff3c48ba2c1426263c3a177525e83f90cd25e81d|46.64|2014-10-26 12:56:00|1.41290891556208|4|20897500000|149|0.6104695895098807|0|33|977|-81.027334|201|34.977331|FRESH HT CHICKEN|11.9|2|FRESH BONELESS CHICKEN BREAST|bea1aab0a475ba6742f2c1e34750b6ef8ee8efda|1.5463774458749717|0.61055446569467375|00208975000005|POULTRY|MEAT|-81.027334|1.4141937624131469|149|2
34.977331|0134f21ffedf700652ecb510ed061d22217fb03a|9.38|2015-01-18 17:22:00|1.41290891556208|4|1600043779|149|0.6104695895098807|0|33|1433|-81.027334|9|34.977331|GRANOLA|0.0|1|NV PROTEIN GRANLA OATS DK CHOC|bea1aab0a475ba6742f2c1e34750b6ef8ee8efda|1.5463774458749717|0.61055446569467375|00016000437784|CEREAL|G1 GROCERY|-81.027334|1.4141937624131469|149|2
34.977331|54dc388dea55a8a1709e646f87febb82935b3f81|5.29|2015-02-10 17:00:00|1.41290891556208|4|7008503535|149|0.6104695895098807|0|33|1277|-81.027334|279|34.977331|FROZEN SNACKS|0.0|5|BAGEL BITES THREE CHEESE|bea1aab0a475ba6742f2c1e34750b6ef8ee8efda|1.5463774458749717|0.61055446569467375|00070085035358|FROZEN SANDWICH AND SNACKS|FROZEN|-81.027334|1.4141937624131469|149|1
34.977331|4e59048b8e78636e5efb76fb18aa4d2ed07c12a2|9.38|2015-02-12 07:45:00|1.41290891556208|4|81829001308|149|0.6104695895098807|0|33|685|-81.027334|61|34.977331|GREEK|2.38|3|CHOBANI 100 VANILLA 4 PK|bea1aab0a475ba6742f2c1e34750b6ef8ee8efda|1.5463774458749717|0.61055446569467375|00818290013101|YOGURT|DAIRY|-81.027334|1.4141937624131469|149|2
34.977331|49143f2195c725b124d93762e66d119429f63e0c|5.38|2014-12-29 06:41:00|1.41290891556208|4|1380016610|149|0.6104695895098807|0|33|1278|-81.027334|48|34.977331|SINGLE SERVE NUTRITIONAL|0.0|5|LC FIESTA G. CHICKEN|bea1aab0a475ba6742f2c1e34750b6ef8ee8efda|1.5463774458749717|0.61055446569467375|00013800101648|FROZEN MEALS|FROZEN|-81.027334|1.4141937624131469|149|2
34.977331|5a92bc1a1da8a48a61ba0bc6e8bd253159cb6b7f|3.19|2015-02-01 21:46:00|1.41290891556208|4|1800081778|149|0.6104695895098807|0|33|326|-81.027334|54|34.977331|COOKIES/BROWNIES-REFRIGERATED|0.0|3|PILLSBURY DELUXE CHOC CHIP|bea1aab0a475ba6742f2c1e34750b6ef8ee8efda|1.5463774458749717|0.61055446569467375|00018000817733|DOUGH PRODUCTS|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|638d31cbf7c7f32a8aa0a7ed4b7eee027f1ae8f5|6.29|2014-10-07 17:57:00|1.41290891556208|4|89470001013|149|0.6104695895098807|0|33|685|-81.027334|61|34.977331|GREEK|0.0|3|CHOBANI 100 VANILLA BLEND|bea1aab0a475ba6742f2c1e34750b6ef8ee8efda|1.5463774458749717|0.61055446569467375|00818290013194|YOGURT|DAIRY|-81.027334|1.4141937624131469|149|1
35.066546|17cdfaf9ddabcaa3572fd5e74a64e9aa28efccc3|5.49|2015-02-25 11:14:00|1.4091206135396188|2|7597116682|45|0.6120266850020475|0|47|1837|-80.771677|420|35.066546|FFM PRESLICED MEATS|0.0|6|FRESH FO0D SMOKED TURKY BREAST|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|0.61242566243833529|00072036959874|PRESLICED MEAT|DELI|-80.771677|1.409731706007376|45|1
35.066546|32b153e3e87d5084dd2aeb636c00170021c3b076|2.65|2014-09-21 12:44:00|1.4091206135396188|2|1600041888|45|0.6120266850020475|0|47|42|-80.771677|6|35.066546|GRANOLA/YOGURT BARS|0.0|1|NV BAR THINS DARK CHOC|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|0.61242566243833529|00016000418882|BREAKFAST FOODS|G1 GROCERY|-80.771677|1.409731706007376|45|1
35.066546|41e6d1c62cadfa6351ab72a9cb99f104a886e73e|2.79|2015-02-03 14:13:00|1.4091206135396188|2|9256714170|45|0.6120266850020475|0|47|6787|-80.771677|1568|35.066546|MAGAZINES MONTHLY|0.0|18|FAMILY CIRCLE|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|0.61242566243833529|00092567141708|MAGAZINES|GM|-80.771677|1.409731706007376|45|1
35.066546|bbdd89eb1cc5e9812996683a3f5a013692a33d12|4.49|2014-10-15 16:03:00|1.4091206135396188|2|2840023847|45|0.6120266850020475|0|47|201|-80.771677|31|35.066546|POTATO CHIPS|0.5|1|SMARTFOOD VARIETY 10 CT|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|0.61242566243833529|00028400238533|SNACKS|G1 GROCERY|-80.771677|1.409731706007376|45|1
35.066546|08c4e9f49ceb1d9b9204d392336761038f5c9857|4.99|2014-10-10 14:31:00|80.782094729586973|2|7203671139|45|35.08115140968583|0|27|141|-80.732725|21|35.082768|TRAIL MIXES AND BLENDS|1.0|1|HT PEANUT LOVERS MOUNTAIN MIX|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|35.102887530186244|00072036711434|NUTS|G1 GROCERY|-80.771677|80.771683162138743|147|1
35.066546|fbfcdeba5782a8b5db9105891bb5b7446cd38daf|4.99|2014-11-03 15:07:00|80.782094729586973|2|7203671139|45|35.081151408993385|0|27|141|-80.8062|21|35.037115|TRAIL MIXES AND BLENDS|1.0|1|HT PEANUT LOVERS MOUNTAIN MIX|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|35.102887530186244|00072036711434|NUTS|G1 GROCERY|-80.771677|80.771685256560431|27|1
35.066546|22e79c874f9f6ae84aacb49a04d9002a288d994a|7.3|2014-12-13 13:28:00|80.782094729586973|2|3010003012|45|35.08115140968583|0|27|91|-80.732725|13|35.082768|SPRAYED BUTTER CRACKERS|2.3|1|KEEBLER CLUB REDUCED FAT|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|35.102887530186244|00030100100706|CRACKERS|G1 GROCERY|-80.771677|80.771683162138743|147|2
35.066546|f7c7ce088bc704c82e1ad22a0587ce9da50df3bf|3.65|2015-01-13 15:28:00|80.782094729586973|2|3010003012|45|35.081151409700041|0|27|91|-80.7007|13|35.06858|SPRAYED BUTTER CRACKERS|1.15|1|KEEBLER CLUB REDUCED FAT|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|35.102887530186244|00030100100706|CRACKERS|G1 GROCERY|-80.771677|80.771683111651782|273|1
35.066546|8dc5992a3c1038c2ec5a4e7fffd3c2e1db0258c2|3.65|2014-12-06 15:06:00|1.4091206135396188|2|3010003012|45|0.6120266850020475|0|47|91|-80.771677|13|35.066546|SPRAYED BUTTER CRACKERS|1.15|1|CLUB MINIS|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|0.61242566243833529|00030100490524|CRACKERS|G1 GROCERY|-80.771677|1.409731706007376|45|1
35.066546|d6fab7136bae35d0469d46da8853bbb9af517811|2.17|2014-11-18 15:32:00|80.782094729586973|2|7433610204|45|35.08115140968583|0|27|331|-80.732725|52|35.082768|NATURAL SLICED|0.0|3|HC MILD CHEDDAR SLICES|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|35.102887530186244|00074336102042|CHEESE|DAIRY|-80.771677|80.771683162138743|147|1
35.066546|363bd8ddd29212789f159f62b9c80e091f9b8295|2.17|2014-10-06 14:40:00|80.782094729586973|2|7433610204|45|35.08115140968583|0|27|331|-80.732725|52|35.082768|NATURAL SLICED|0.0|3|HC MILD CHEDDAR SLICES|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|35.102887530186244|00074336102042|CHEESE|DAIRY|-80.771677|80.771683162138743|147|1
35.066546|23faf3817c043d2f36a11674b080d728dc65d457|2.89|2015-01-20 12:05:00|1.4091206135396188|2|7203655029|45|0.6120266850020475|0|47|331|-80.771677|52|35.066546|NATURAL SLICED|1.22|3|HT MEDIUM CHEDDAR SLICES|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|0.61242566243833529|00072036983930|CHEESE|DAIRY|-80.771677|1.409731706007376|45|1
35.066546|ce651c3066c9be6861f14c86e4e864adcb51f735|8.67|2015-02-11 16:32:00|80.782094729586973|2|7203655029|45|35.08115140968583|0|27|331|-80.732725|52|35.082768|NATURAL SLICED|3.67|3|HT MEDIUM CHEDDAR SLICES|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|35.102887530186244|00072036983930|CHEESE|DAIRY|-80.771677|80.771683162138743|147|3
35.066546|43c8191e0ae15f142a6186d080c3fd64c14ebb5e|2.89|2014-12-28 14:12:00|80.782094729586973|2|7203655029|45|35.081151404764753|0|27|331|-80.709466|52|35.124987|NATURAL SLICED|1.22|3|HT MEDIUM CHEDDAR SLICES|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|35.102887530186244|00072036983930|CHEESE|DAIRY|-80.771677|80.77169289298493|157|1
35.066546|ad4788c344456461ed946bb71125933b6b5a004a|2.89|2015-03-07 18:21:00|80.782094729586973|2|7203655029|45|35.08115140968583|0|27|331|-80.732725|52|35.082768|NATURAL SLICED|0.92|3|HT MEDIUM CHEDDAR SLICES|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|35.102887530186244|00072036983930|CHEESE|DAIRY|-80.771677|80.771683162138743|147|1
35.066546|23211d05ceea0327f00b0935fe5a6b073f20fb94|2.89|2014-11-10 13:37:00|80.782094729586973|2|7203655029|45|35.08115140968583|0|27|331|-80.732725|52|35.082768|NATURAL SLICED|1.45|3|HT MEDIUM CHEDDAR SLICES|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|35.102887530186244|00072036983930|CHEESE|DAIRY|-80.771677|80.771683162138743|147|1
35.066546|09cde2c5f04238a4286ee7cfd8e05ad7f4e9df13|6.49|2014-09-23 08:59:00|80.782094729586973|2|7703401130|45|35.08115140968583|0|27|141|-80.732725|21|35.082768|TRAIL MIXES AND BLENDS|1.5|1|SECOND NATURE CHOC MEDLEY|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|35.102887530186244|00077034011494|NUTS|G1 GROCERY|-80.771677|80.771683162138743|147|1
35.066546|e4a4baec4e3be8b4e982a9a58b6e7b66efc050e9|4.97|2014-10-21 17:18:00|80.782094729586973|2|7229000227|45|35.08115140968583|0|27|1271|-80.732725|41|35.082768|PROTEIN BREAKFAST|0.0|5|TENN PRIDE SAUS&BTTRMLK BISC|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|35.102887530186244|00072290002279|BREAKFAST FOODS FROZEN|FROZEN|-80.771677|80.771683162138743|147|1
35.066546|775c9160faef99e52c10f4b2cb6ddb36e1cdb9f8|4.97|2015-02-21 16:26:00|80.782094729586973|2|7229000227|45|35.081151409700041|0|27|1271|-80.7007|41|35.06858|PROTEIN BREAKFAST|0.0|5|TENN PRIDE SAUS&BTTRMLK BISC|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|35.102887530186244|00072290002279|BREAKFAST FOODS FROZEN|FROZEN|-80.771677|80.771683111651782|273|1
35.066546|1f3d2d0a127236e71b673ff4da326f3d656fca82|5.99|2014-12-23 14:06:00|80.782094729586973|2|7244014076|45|35.081151404300165|0|27|6791|-80.739|1568|35.141204|MAGAZINES ANNUAL|0.0|18|14076 BHG: WEEKEND MAKEOVER|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|35.102887530186244|00072440140769|MAGAZINES|GM|-80.771677|80.771693518131428|171|1
35.066546|07787693f12033f698f027d316d3c897f6b41f77|13.98|2015-01-05 10:39:00|1.4091206135396188|2|8558201232|45|0.6120266850020475|0|47|84|-80.771677|11|35.066546|CONDIMENTS-DSD VENDORS|7.0|1|VIRGINIA DINER UNC SALTED|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|0.61242566243833529|00085582012320|CONDIMENTS|G1 GROCERY|-80.771677|1.409731706007376|45|2
35.066546|22c08f9fa179132de5cea68c2fec5a4d7b7fd636|9.98|2015-01-26 16:28:00|80.782094729586973|2|7756706153|45|35.08115140968583|0|27|273|-80.732725|43|35.082768|PREMIUM NOVELTIES|2.98|5|BREYERS CARB SMART ALMOND BAR|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|35.102887530186244|00077567061539|FROZEN NOVELTIES|FROZEN|-80.771677|80.771683162138743|147|2
35.066546|737a6f54f69ef83e6313725347d87adef5e742e8|2.9699999999999998|2015-01-01 12:35:00|80.782094729586973|2|7641090275|45|35.08115140968583|0|27|166|-80.732725|21|35.082768|FRONT END NUTS|0.30000000000000004|1|LANCESALTED PEANUTS PP .99|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|35.102887530186244|00076410902753|NUTS|G1 GROCERY|-80.771677|80.771683162138743|147|3
35.066546|1d45bf74ec346ee0706df1a23f9dbad53313a834|2.97|2015-03-07 18:29:00|80.782094729586973|2|7468812100|45|35.08115140968583|0|27|423|-80.732725|72|35.082768|NFS-DISPOSE PLATES/BOWLS|0.0|1|"EASY WAY 9"" PAPER PLATES"|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|35.102887530186244|00074688121005|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.771677|80.771683162138743|147|1
35.066546|e5f68bf9e0d1f64c7e5026b11386930c49950740|1.89|2014-11-26 11:14:00|80.782094729586973|2|1300079630|45|35.08115140968583|0|27|69|-80.732725|26|35.082768|CANNED GRAVY|0.55|1|HEINZ GRAVY CHICKEN|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|35.102887530186244|00013000798204|PREPARED FOODS-DRY MIXES|G1 GROCERY|-80.771677|80.771683162138743|147|1
35.066546|886be220193048df4ea790450e4dcbdb76b3eac6|3.49|2015-01-12 15:46:00|1.4091206135396188|2|2389649770|45|0.6120266850020475|0|47|200|-80.771677|31|35.066546|MICROWAVE POPCORN|0.0|1|POP SECRET JMBO POP MOVIE BUTR|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|0.61242566243833529|00023896362700|SNACKS|G1 GROCERY|-80.771677|1.409731706007376|45|1
35.066546|f8f9b2adaff49b35ee18d5927215809b6166cc14|2.5|2014-10-12 13:05:00|80.782094729586973|2|4480000102|45|35.08115140968583|0|27|223|-80.732725|35|35.082768|SUGAR SUBSTITUTES|0.0|1|SWEET-N-LOW GRANULATED 100 PK|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|35.102887530186244|00044800001027|SUGAR/SUBSTITUTES|G1 GROCERY|-80.771677|80.771683162138743|147|1
35.066546|93d40cb04a04df60ae16fce062e8d7a123db8357|4.79|2014-11-05 15:50:00|1.4091206135396188|2|2310010327|45|0.6120266850020475|0|47|155|-80.771677|24|35.066546|NFS-DOG TREATS|0.0|1|CESAR SOFTIES FILET MIGNON TRT|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|0.61242566243833529|00023100103273|PET FOOD/SUPPLIES|G1 GROCERY|-80.771677|1.409731706007376|45|1
35.066546|71fa0be6a9a82f37777708b4af7bee0f65276205|9.99|2015-01-01 12:41:00|80.782094729586973|2|7726009983|45|35.08115140968583|0|27|727|-80.732725|7|35.082768|SEASONAL CANDY-SINGLE FAC|5.0|1|I/O(C14)RS PECAN DELIGHT BOX|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|35.102887530186244|00077260099839|CANDY|G1 GROCERY|-80.771677|80.771683162138743|147|1
35.066546|6cc9a872e3a13057d29c9b37124e1f71b766f28d|15.98|2014-12-13 13:37:00|80.782094729586973|2|30031872120|45|35.08115140968583|0|27|4236|-80.732725|1200|35.082768|DEX ADULT/CHILDREN|6.0|17|ROBITUSSIN PEAKCLD CHST DM MAX|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|35.102887530186244|00300318738122|COUGH/COLD/SINUS|HBC|-80.771677|80.771683162138743|147|2
35.066546|cbdb6447030b56e6eca319bdcd00ff09b1f617e4|2.85|2014-09-25 14:39:00|80.782094729586973|2|1380010321|45|35.08115140968583|0|27|1279|-80.732725|48|35.082768|SINGLE SERVE FLAVOR|0.0|5|STOUFFER HOMESTYLE MEAT LOAF|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|35.102887530186244|00013800100726|FROZEN MEALS|FROZEN|-80.771677|80.771683162138743|147|1
35.066546|51ac24642d832ccf5d2369648a5926ba71b4e04e|6.49|2015-03-02 14:53:00|80.782094729586973|2|4154800385|45|35.08115140968583|0|27|252|-80.732725|45|35.082768|PREMIUM ICE CREAM|1.61|5|EDY'S SLOW CHURNED NEOPOLITA|bf638225bfb4a746db6775347e74cac19e7bf7f6|1.0091985986518812|35.102887530186244|00041548740867|ICE CREAM|FROZEN|-80.771677|80.771683162138743|147|1
35.04711|5b68265e48ef23788f80ea06e0254082ca7b3547|2.0|2014-12-19 18:35:00|80.648225123995502|3|2840019079|129|35.068866225888307|0|30|201|-80.562829|31|35.006282|POTATO CHIPS|0.0|1|MUNCHOS|c7b45e477813e8af1039d22973990f1e47eadaef|1.5033026706250208|35.078006462436761|00028400190794|SNACKS|G1 GROCERY|-80.64817|80.648171038438633|60|1
35.04711|9d2d7e764d08b0fdad60204f1138b68c99387a46|8.99|2014-10-10 20:18:00|80.648225123995502|3|8200072385|129|35.068866220600434|0|30|461|-80.699909|84|35.002628|FLAVORED MALT BEVERAGE|0.0|16|SMIRNOFF ICE 6PK BOTTLE|c7b45e477813e8af1039d22973990f1e47eadaef|1.5033026706250208|35.078006462436761|00082000723851|SPECIALTY|BEER|-80.64817|80.64818855973958|477|1
35.04711|b2f1fd7820458ba78f1e5aae82a5d4172394d243|3.89|2014-10-03 18:00:00|1.4091206135396188|3|3800039118|129|0.6116874628086298|0|47|81|-80.64817|9|35.04711|RTE CEREAL KIDS|1.9|1|KELLOGG FROOT LOOPS 12.2|c7b45e477813e8af1039d22973990f1e47eadaef|1.5033026706250208|0.61242566243833529|00038000391187|CEREAL|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|505cefc9580cf306bf70e63a27910ac51b028b03|1.77|2015-01-05 17:21:00|1.4091206135396188|3|7203657031|129|0.6116874628086298|0|47|322|-80.64817|53|35.04711|SOUR CREAM|0.52|3|HT SOUR CREAM|c7b45e477813e8af1039d22973990f1e47eadaef|1.5033026706250208|0.61242566243833529|00072036570314|CULTURES|DAIRY|-80.64817|1.407576102208115|129|1
35.04711|a72ca07b2fc4cad3a854aa6e3ac5f1364b730cf9|3.33|2015-01-08 18:22:00|1.4091206135396188|3|7203643010|129|0.6116874628086298|0|47|252|-80.64817|45|35.04711|PREMIUM ICE CREAM|0.0|5|HT SMTH & CRMY COFFEE IC|c7b45e477813e8af1039d22973990f1e47eadaef|1.5033026706250208|0.61242566243833529|00072036981769|ICE CREAM|FROZEN|-80.64817|1.407576102208115|129|1
35.04711|901b1e534ec8d3ab25ef7dfe227a0545940e41d9|5.99|2015-03-04 15:35:00|80.648225123995502|3|76108880156|129|35.068866220199766|0|30|1939|-80.699686|465|35.000049|COLD PREP FOODS SIDES|0.0|6|MACARONI & CHEESE FAMILY SIZE|c7b45e477813e8af1039d22973990f1e47eadaef|1.5033026706250208|35.078006462436761|00761088801568|COLD PREPARED FOODS|DELI|-80.64817|80.648189247923554|249|1
35.667941|0637f4e8940eddcdddb3c7e520f8a9446d17b9cc|2.69|2014-10-18 18:30:00|80.497482303704658|4|7225001125|178|35.748699262477309|0|6|1025|-80.605588|162|35.43259|WHITE|0.0|7|MERITA OLD FASHIONED 20 OZ|c9f9922d888cf1f9687cd7a88495f19d4945522e|5.580225084605056|35.699188602026126|00072250011259|SLICED BREAD|COMMERCIAL BAKERY|-80.497332|80.497624735461429|202|1
35.412407|db68c2a71c0b03773c5b5170cfc6f1691c16d820|8.3|2015-01-05 16:37:00|80.606823361882718|4|7203646021|68|35.495988310188714|0|57|1463|-80.66939|42|35.28326|REGULAR FROZEN FRUIT|0.0|5|HT BERRY MEDLEY|cc3f7f4fc134576ed9addf733b730c4bcad0f890|5.77527213742783|35.500309569604553|00072036460622|FROZEN FRUIT|FROZEN|-80.662946|80.66308689801113|46|2
35.412407|b8ea8f963311c7d82a54704c8f7bd9ac5f6411e8|2.49|2014-12-24 17:14:00|80.606823361882718|4|7203688048|68|35.495988310188714|0|57|526|-80.66939|64|35.28326|FRESH MUSHROOMS|0.0|4|HT SLICED BABY BELLAS|cc3f7f4fc134576ed9addf733b730c4bcad0f890|5.77527213742783|35.500309569604553|00072036880482|FRESH PRODUCE|PRODUCE|-80.662946|80.66308689801113|46|1
35.412407|2642372b05cdcf3cdb5773ed7185338f7aa8261a|3.39|2015-01-09 13:15:00|80.606823361882718|4|5260305445|68|35.495988310188714|0|57|214|-80.66939|33|35.28326|BROTH|0.0|1|PACIFIC ORG LS FR CHICKN BROTH|cc3f7f4fc134576ed9addf733b730c4bcad0f890|5.77527213742783|35.500309569604553|00052603054454|SOUP|G1 GROCERY|-80.662946|80.66308689801113|46|1
35.412407|002adab3823611d2c53cfdea2ffc249540dad516|4.59|2014-12-29 12:16:00|80.606823361882718|4||68|35.495988289841172|0|57|529|-80.737839|64|35.297134|FRESH ASPARAGUS|0.0|4|PURPLE ASPARAGUS|cc3f7f4fc134576ed9addf733b730c4bcad0f890|5.77527213742783|35.500309569604553|00203079000005|FRESH PRODUCE|PRODUCE|-80.662946|80.663104045303285|258|1
35.412407|88d78c7e7a4b60c5189443569f17172acca3a642|7.99|2014-12-11 16:54:00|80.606823361882718|4|70587510016|68|35.495988310188714|0|57|4522|-80.66939|1215|35.28326|SPLMNT-CARDIO/CHOLESTEROL|1.6|17|BARLEANS FORTI-FLAX|cc3f7f4fc134576ed9addf733b730c4bcad0f890|5.77527213742783|35.500309569604553|00705875100168|VITAMINS & SUPPLEMENTS|HBC|-80.662946|80.66308689801113|46|1
35.412407|d78fb43a78e0b06f33b4ab80f9cb777d1aa6ced0|4.47|2014-11-29 15:05:00|80.606823361882718|4|7203663085|68|35.495988310188714|0|57|1132|-80.66939|55|35.28326|EGGS SUBSTITUTES|0.0|3|HARRIS TEETER LIQUID EGG PROD|cc3f7f4fc134576ed9addf733b730c4bcad0f890|5.77527213742783|35.500309569604553|00072036630858|EGGS FRESH|DAIRY|-80.662946|80.66308689801113|46|1
34.977331|b7597e7d46f73e8d4a1a1b2e54870bfe54b01e0c|6.79|2014-10-31 13:44:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|31148677b4b5bfd2c945a4271f6073529d160b17|6.79|2014-12-30 12:03:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|477d890779a4f80bd84968a3aee137fb0216e980|6.79|2014-11-28 15:57:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|88fd5a662a43648791fe7ea417dc00e5834cdfda|6.79|2014-12-05 18:06:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|3cce3621e535eda5a043fb65be17ab9f92101746|6.79|2014-09-19 11:39:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|5b73e23b5f70ee0fb180f0777393e90b65bce639|6.79|2015-02-20 13:43:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|f7153413136f72b52a32ef9341b555c2c4c0948b|6.79|2014-11-14 13:18:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.8|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|10d1030ededc19f48902aa486e2c3f0bd3a6ec30|6.79|2015-02-27 16:27:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|677771174e2d3954dc8626d2194fd91af5d00647|6.79|2014-12-19 17:17:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|87b13d828924033837915679f38bf84554864754|6.79|2015-01-09 17:13:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|c93d10c4448f18d1117c81c5dbcb97bfbdcb5e0e|6.79|2015-01-23 15:14:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|7e87215bca05cd7e368db91ff998069a0c4fcfb9|6.79|2014-12-12 14:54:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.8|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|e97091f5f917f27986d730cfb9dd42084d6f172a|6.79|2015-02-06 15:11:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|6ebd060bafff58f7844eb8f1775f7b566b2f9c9b|6.79|2014-09-26 15:03:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|906301c8d76df28a4b342ff85c608b9e2e9ff06d|6.79|2015-01-16 12:43:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.8|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|b56db24e2685c7181ccc4173ed729b88ea48b2d7|6.79|2015-02-14 10:05:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.8|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|1085ac4325119b298d6c35de5a009413bdc6adc8|6.79|2015-01-30 16:30:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|64c45a0ea4bad21ccbc9b9e9ec041e5035cd191e|6.79|2014-10-03 12:55:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.8|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|02ef606566fa92550c061898640baf098955772c|6.79|2015-01-02 14:05:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|5a52a59239770e4facac513c673c0089782fd996|6.79|2014-10-10 16:10:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|01b8c549e08aaa6a0b1379512dca4602dcac1b6a|6.79|2014-12-26 15:45:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|f20d2445fff15d7d399a1e6ba2a31f74779fd618|6.79|2014-11-21 13:03:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|f32fc284ad970932c8e338424d55714d2399e6d6|6.79|2015-03-07 13:50:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|e58a7050039c9bd7aaf796fcc52271bad0c5967f|6.79|2014-10-25 11:21:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|1b9cce9a55f488fcbbd20044bfcea41e12486dd5|6.79|2014-11-07 12:52:00|1.41290891556208|2|4850001833|149|0.6104695895098807|1|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA ORIGINAL|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00048500018330|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|533578b5427de32a0bf53bd111fe69e8ade03ad0|2.99|2014-10-17 14:44:00|1.41290891556208|2|7062266666|149|0.6104695895098807|1|33|52|-81.027334|7|34.977331|PKG NON CHOC|0.4|1|GOETZE'S CARAMEL CREMES|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00070622666663|CANDY|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|1c8d9643dbea3e9e91b87c43833babdcc363de7c|2.99|2014-09-12 12:18:00|1.41290891556208|2|7062266666|149|0.6104695895098807|1|33|52|-81.027334|7|34.977331|PKG NON CHOC|0.6|1|GOETZE'S CARAMEL CREMES|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00070622666663|CANDY|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|04dd9438343f42ddac91f5d924a6ce0595f065a7|22.99|2014-12-14 18:14:00|1.41290891556208|2|3680024421|149|0.6104695895098807|0|33|4186|-81.027334|1200|34.977331|ALLERGY REMEDY-ADULT|7.99|17|TC A/D ALLRGY-CETIRIZINE 10MG|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00036800244214|COUGH/COLD/SINUS|HBC|-81.027334|1.4141937624131469|149|1
34.977331|2f4289ef224ceb7b0fbbf89630a9b34afcc4c549|8.67|2014-12-18 22:56:00|1.41290891556208|2|7203663102|149|0.6104695895098807|0|33|339|-81.027334|57|34.977331|EGGNOGS/DRINKS|2.67|3|I/O HARRIS TEETER EGG NOG|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00072036631022|MILK|DAIRY|-81.027334|1.4141937624131469|149|3
34.977331|eac901b1fa98b0ed2c49a18f78852eec35c31644|7.99|2014-12-27 10:12:00|1.41290891556208|2|4242150024|149|0.6104695895098807|1|33|1839|-81.027334|420|34.977331|BH PRESLICED MEATS|0.0|6|BH PRE-SLICED HONEY SMK TURKEY|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00042421500240|PRESLICED MEAT|DELI|-81.027334|1.4141937624131469|149|1
34.977331|bbc3ec7a1fc37db53f9f4f0a5fd5530d16f4045c|13.58|2015-02-21 18:06:00|1.41290891556208|2|7064003404|149|0.6104695895098807|0|33|252|-81.027334|45|34.977331|PREMIUM ICE CREAM|5.62|5|B BUNNY VANILLA ICE CREAM|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00070640034017|ICE CREAM|FROZEN|-81.027334|1.4141937624131469|149|2
34.977331|7843d132ab08496465d7c5e695fcb5c679527a22|7.16|2015-03-03 20:08:00|1.41290891556208|2|5200033875|149|0.6104695895098807|0|33|171|-81.027334|20|34.977331|ISOTONIC DRINKS|3.16|1|GATORADE FROST GLACIER FREEZE|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00052000320169|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-81.027334|1.4141937624131469|149|4
34.977331|7365e41f708b560abf3ecabce1e13362a6278c2d|7.18|2014-10-21 21:06:00|1.41290891556208|2|4400002734|149|0.6104695895098807|0|33|1253|-81.027334|12|34.977331|ALL OTHER COOKIES|0.0|1|NILLA WAFERS|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00044000027346|COOKIES|G1 GROCERY|-81.027334|1.4141937624131469|149|2
34.977331|538b9a5bd02c0c9644c61873dd4ece1bbda357f9|7.99|2014-12-30 14:17:00|1.41290891556208|2|30031872120|149|0.6104695895098807|0|33|4236|-81.027334|1200|34.977331|DEX ADULT/CHILDREN|3.0|17|ROBITUSSIN PEAKCLD CHST DM MAX|cd417bd757e2f6b232ace6b944b7e169c06e08eb|0.44054116033638774|0.61055446569467375|00300318738122|COUGH/COLD/SINUS|HBC|-81.027334|1.4141937624131469|149|1
35.372142|065beb7bde33ecc2cba4bcf499e983f6479d4cbf|2.49|2015-02-14 08:31:00|80.779636304526477|0|60504939530|122|35.385245021190308|0|17|509|-80.86175|64|35.40953|FRESH CITRUS-REMAINING|0.0|4|LEMONS, SMALL 1LB BAG|cde5133718177388c556cb0046d9a2d38769d901|0.9053871219799431|35.392509581117899|00605049395300|FRESH PRODUCE|PRODUCE|-80.782849|80.782849473627735|209|1
34.937113|0d88d7b8a18e1bc3051c04d1fd925a1a5cc9df62|8.99|2014-10-03 00:09:00|80.856688219393845|4|79327199036|372|35.132464164535428|0|15|458|-80.85753|82|35.116638|CRAFT BEER|0.0|16|DUCK RABBIT MILK STOUT|d2a5aaa1e7ffd96c648c9f8fab7a4a1b675c4366|13.498315172500552|35.134355925261694|00793271990360|DOMESTIC BEER|BEER|-80.837892|80.838317422080024|204|1
34.937113|a124f3f0185d948697f83865525b7f92fd9ce630|0.97|2014-09-28 18:59:00|80.856688219393845|4|7203608070|372|35.132464164535428|0|15|68|-80.85753|11|35.116638|BARBECUE SAUCES|0.0|1|HT BBQ SC ORIGINAL|d2a5aaa1e7ffd96c648c9f8fab7a4a1b675c4366|13.498315172500552|35.134355925261694|00072036080707|CONDIMENTS|G1 GROCERY|-80.837892|80.838317422080024|204|1
34.937113|ab5bb7abb8e4d78094340d0782e7679f9b7be296|2.99|2014-12-10 12:53:00|80.856688219393845|4|7203670325|372|35.132464456720307|0|15|444|-81.027334|76|34.977331|NFS-PLASTIC WRAPS|0.49|1|YH PLASTIC WRAP|d2a5aaa1e7ffd96c648c9f8fab7a4a1b675c4366|13.498315172500552|35.134355925261694|00072036703255|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.837892|80.837995494089057|149|1
34.937113|88b1a104cf971904b7f92404cd15e137088076ba|5.49|2015-01-18 18:04:00|80.856688219393845|4|827411111|372|35.132464164535428|0|15|55|-80.85753|8|35.116638|REGULAR|0.0|23|VIRGILS CREAM SODA|d2a5aaa1e7ffd96c648c9f8fab7a4a1b675c4366|13.498315172500552|35.134355925261694|00090341543212|CARBONATED BEVERAGES|BEVERAGE|-80.837892|80.838317422080024|204|1
34.937113|6ceeff46e7110b537518386736ab6130621bb305|6.19|2015-01-10 23:58:00|80.856688219393845|4|7214011047|372|35.132464164535428|0|15|4842|-80.85753|1235|35.116638|FIRST AID LOTION|0.0|17|AQUAPHOR HEALING OINTMENT|d2a5aaa1e7ffd96c648c9f8fab7a4a1b675c4366|13.498315172500552|35.134355925261694|00072140110475|FIRST AID|HBC|-80.837892|80.838317422080024|204|1
34.937113|f7776f5e3878b406c3a8d6f37dfbb6b7d0464c23|9.99|2014-12-20 15:59:00|80.856688219393845|4|7203678030|372|35.132464164535428|0|15|458|-80.85753|82|35.116638|CRAFT BEER|0.0|16|HT CREATE YOUR OWN SAMPLER|d2a5aaa1e7ffd96c648c9f8fab7a4a1b675c4366|13.498315172500552|35.134355925261694|00072036780300|DOMESTIC BEER|BEER|-80.837892|80.838317422080024|204|1
34.937113|b2a9d6008b69d572ef0ba4465b7bfd19544a48d3|3.79|2014-12-12 12:46:00|80.856688219393845|4|7203688014|372|35.132464456720307|0|15|581|-81.027334|136|34.977331|FRESH SALSA|0.0|4|HT FRESH MILD SALSA|d2a5aaa1e7ffd96c648c9f8fab7a4a1b675c4366|13.498315172500552|35.134355925261694|00072036880215|OTHER MERCHANDISE|PRODUCE|-80.837892|80.837995494089057|149|1
34.937113|dd7727a59ed76d082a40a1ffb63ef0d5e29857b9|4.49|2014-10-31 09:40:00|80.856688219393845|4|4100009003|372|35.132464164535428|0|15|233|-80.85753|37|35.116638|BLACK TEA|0.0|1|LIPTON TEA COLD BREW FAMILY|d2a5aaa1e7ffd96c648c9f8fab7a4a1b675c4366|13.498315172500552|35.134355925261694|00041000090035|TEA|G1 GROCERY|-80.837892|80.838317422080024|204|1
34.937113|d6e9065cd7b4911567fc0cc4dea39850c178d7e1|6.57|2015-02-27 14:56:00|80.856688219393845|4|4900005010|372|35.132464164535428|0|15|54|-80.85753|8|35.116638|DIET|0.8500000000000001|23|DT SPRITE ZERO  2 LITER|d2a5aaa1e7ffd96c648c9f8fab7a4a1b675c4366|13.498315172500552|35.134355925261694|00049000050172|CARBONATED BEVERAGES|BEVERAGE|-80.837892|80.838317422080024|204|3
34.937113|a8526dab99364ffb2e8b6a6c8bb0401a089f5736|4.38|2014-10-10 00:16:00|80.856688219393845|4|4900005010|372|35.132464164535428|0|15|54|-80.85753|8|35.116638|DIET|1.09|23|DT SPRITE ZERO  2 LITER|d2a5aaa1e7ffd96c648c9f8fab7a4a1b675c4366|13.498315172500552|35.134355925261694|00049000050172|CARBONATED BEVERAGES|BEVERAGE|-80.837892|80.838317422080024|204|2
34.937113|95a8949f2c580cd32181418db19a2bc4cf5142e7|9.99|2014-12-05 18:23:00|80.856688219393845|4|7203601062|372|35.132464164535428|0|15|640|-80.85753|201|35.116638|MARINATED POULTRY|0.0|2|HT ROTISSERIE TURKEY TENDER|d2a5aaa1e7ffd96c648c9f8fab7a4a1b675c4366|13.498315172500552|35.134355925261694|00072036010629|POULTRY|MEAT|-80.837892|80.838317422080024|204|1
34.937113|34efe59aedfb5ab74445b53c3a644ed577464ace|11.99|2014-11-22 18:46:00|80.856688219393845|4|3760025836|372|35.132464164535428|0|15|638|-80.85753|137|35.116638|MARINATED PORK|0.0|2|HRML MESQUITE PORK FILET|d2a5aaa1e7ffd96c648c9f8fab7a4a1b675c4366|13.498315172500552|35.134355925261694|00037600497671|PORK|MEAT|-80.837892|80.838317422080024|204|1
35.053394|d0669757cbb3d6c382f6a9fec6f15c4f455903ab|2.79|2015-01-16 17:29:00|80.848351720559364|4||11|35.077351214610943|0|25|522|-80.850065|64|35.030252|FRESH TOMATOES|0.0|4|RED H/H TOMATOES, BULK|d71d02122de125e7370b55201049d8124c0aca1c|1.6553857258971414|35.082633588753836|00204799000009|FRESH PRODUCE|PRODUCE|-80.848528|80.84853525720753|470|1
35.053394|82e5defa4425d96686b0054f768a8558e50d9aca|1.79|2014-11-02 11:10:00|80.848351720559364|4|7203688032|11|35.077351214610943|0|25|555|-80.850065|64|35.030252|PACKAGED SALADS|0.0|4|HT SHREDDED ICEBERG LETTUCE|d71d02122de125e7370b55201049d8124c0aca1c|1.6553857258971414|35.082633588753836|00072036880321|FRESH PRODUCE|PRODUCE|-80.848528|80.84853525720753|470|1
35.053394|edec6b0adc474c1fc608b00d9017f67f48ae400c|5.98|2014-11-28 10:16:00|80.848351720559364|4|1090000510|11|35.077351214610943|0|25|442|-80.850065|76|35.030252|NFS-COOKING-STORAGE BAGS|0.99|1|REYNOLDS OVEN BAGS-TURKEY|d71d02122de125e7370b55201049d8124c0aca1c|1.6553857258971414|35.082633588753836|00010900005104|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.848528|80.84853525720753|470|2
35.053394|8885df458efc81ee2fd6322014214e072699265e|2.69|2015-01-22 09:22:00|80.848351720559364|4|7225001125|11|35.077351214610943|0|25|1025|-80.850065|162|35.030252|WHITE|0.7|7|MERITA OLD FASHIONED 20 OZ|d71d02122de125e7370b55201049d8124c0aca1c|1.6553857258971414|35.082633588753836|00072250011259|SLICED BREAD|COMMERCIAL BAKERY|-80.848528|80.84853525720753|470|1
35.053394|36eee32d489ccb22a24063f4378f7fdd720affda|7.99|2014-11-02 11:11:00|80.848351720559364|4|2301200207|11|35.077351214610943|0|25|1475|-80.850065|485|35.030252|SUSHI CLASSIC|0.0|6|CRUNCHY SHRIMP ROLL|d71d02122de125e7370b55201049d8124c0aca1c|1.6553857258971414|35.082633588753836|00023012002077|SUSHI|DELI|-80.848528|80.84853525720753|470|1
35.053394|50bb3bb27bda9cce50d38e57ac4614fd2e56397d|3.97|2014-12-28 10:29:00|80.848351720559364|4|7203659020|11|35.077351214610943|0|25|312|-80.850065|51|35.030252|BUTTER|0.0|3|HARRIS TEETER BUTTER QUARTERS|d71d02122de125e7370b55201049d8124c0aca1c|1.6553857258971414|35.082633588753836|00072036590206|BUTTER & MARGARINE|DAIRY|-80.848528|80.84853525720753|470|1
35.444064|89bab7a5728404690ad2e20f2a4e850778af59c9|16.59|2015-01-11 13:10:00|1.4102725052409182|4|20254300000|121|0.6186156170875914|0|1|299|-80.995484|49|35.444064|ANGUS BEEF|5.59|2|VALUE PK ANGUS STEW MEAT|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|0.61833652052202714|00202543000008|BEEF|MEAT|-80.995484|1.413637875046387|121|1
35.444064|a4c5a2fa9b4f9c4ba2a3b14217f61036dd43f249|6.99|2015-01-25 12:46:00|1.4102725052409182|4|3320009553|121|0.6186156170875914|0|1|389|-80.995484|66|35.444064|NFS-LAUNDRY DETERGENTS|3.0|1|A&H CLEAN MEADOW W/OXI CLEAN|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|0.61833652052202714|00033200095545|DETERGENTS|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|61670cf0694c96fd8cd02d4fb19ba390e593e99c|13.98|2014-10-26 11:41:00|1.4102725052409182|4|3320009553|121|0.6186156170875914|0|1|389|-80.995484|66|35.444064|NFS-LAUNDRY DETERGENTS|3.5|1|A&H CLEAN MEADOW W/OXI CLEAN|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|0.61833652052202714|00033200095545|DETERGENTS|G1 GROCERY|-80.995484|1.413637875046387|121|2
35.444064|18042b32ff897293cb8355bf155c1f643589b271|12.58|2015-02-14 14:32:00|1.4102725052409182|4|3320009991|121|0.6186156170875914|0|1|389|-80.995484|66|35.444064|NFS-LAUNDRY DETERGENTS|3.15|1|A&H CLEAN BURST|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|0.61833652052202714|00033200099901|DETERGENTS|G1 GROCERY|-80.995484|1.413637875046387|121|2
35.444064|7829f28cfbeb2bd1bef156e83ba7efb230bb9284|6.38|2014-09-28 10:30:00|1.4102725052409182|4|2733100032|121|0.6186156170875914|0|1|495|-80.995484|108|35.444064|NON REFRIGERATED|1.6|19|LA BANDERITA TORTILLA 10 INCH|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|0.61833652052202714|00027331000363|TORTILLAS|CASE READY MEATS|-80.995484|1.413637875046387|121|2
35.444064|de50dde0f157c9af1a301906eb2a950dcfd6b7de|3.19|2015-01-20 13:39:00|1.4102725052409182|4|2733100032|121|0.6186156170875914|0|1|495|-80.995484|108|35.444064|NON REFRIGERATED|0.0|19|LA BANDERITA TORTILLA 10 INCH|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|0.61833652052202714|00027331000363|TORTILLAS|CASE READY MEATS|-80.995484|1.413637875046387|121|1
35.444064|6de428c9877984fc7f7ad26a7123763b503a7ae3|6.38|2015-03-08 14:31:00|1.4102725052409182|4|2733100032|121|0.6186156170875914|0|1|495|-80.995484|108|35.444064|NON REFRIGERATED|0.0|19|LA BANDERITA TORTILLA 10 INCH|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|0.61833652052202714|00027331000363|TORTILLAS|CASE READY MEATS|-80.995484|1.413637875046387|121|2
35.444064|58925894fb44740a4aaea25380df713c00194c09|3.99|2014-10-30 18:10:00|1.4102725052409182|4|7835470843|121|0.6186156170875914|0|1|317|-80.995484|52|35.444064|CHUNK AND BAR CHEESE|1.49|3|CABOT SERIOUSLY SHARP YELLOW|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|0.61833652052202714|00078354717288|CHEESE|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|db58abfc0dc63e67932505609eefcd7f0c5d5c59|15.48|2014-12-14 10:18:00|1.4102725052409182|4|20600100000|121|0.6186156170875914|0|1|1802|-80.995484|400|35.444064|FFM HAM|4.65|6|VIRGINIA BAKED HAM|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|0.61833652052202714|00206001000005|FFM MEAT|DELI|-80.995484|1.413637875046387|121|1
35.444064|7396aabf0f721d8352b6dcf35eca4d7ab86ca0e1|5.99|2014-11-16 12:52:00|1.4102725052409182|4|3338314605|121|0.6186156170875914|0|1|509|-80.995484|64|35.444064|FRESH CITRUS-REMAINING|0.0|4|CLEMENTINES 3LB|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|0.61833652052202714|00072240133817|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|b977814abf82b72fb5b24db1e3862ce549254aa8|7.99|2015-02-01 12:16:00|1.4102725052409182|4|4242150024|121|0.6186156170875914|0|1|1839|-80.995484|420|35.444064|BH PRESLICED MEATS|1.5|6|BH PRE-SLICED HONEY SMK TURKEY|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|0.61833652052202714|00042421500240|PRESLICED MEAT|DELI|-80.995484|1.413637875046387|121|1
35.444064|446e40d4bcc6e29a1a9779a345462c9e053f55e7|19.98|2015-02-22 13:24:00|1.4102725052409182|4|4200044517|121|0.6186156170875914|0|1|426|-80.995484|72|35.444064|NFS-PAPER TOWELS|4.49|1|BRAWNY 6 BIG ROLL PICK A SIZE|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|0.61833652052202714|00042000445177|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.995484|1.413637875046387|121|2
35.444064|fd1064738af83b95a197f2374429a2504f118b0d|7.98|2015-03-01 13:16:00|1.4102725052409182|4|4300000037|121|0.6186156170875914|0|1|228|-80.995484|36|35.444064|TABLE SYRUP|2.0|1|LOG CABIN SYRUP|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|0.61833652052202714|00043000000373|TABLE SYRUPS|G1 GROCERY|-80.995484|1.413637875046387|121|2
35.444064|8c33c9e8c5fd9626b2b4a67896578d4f868df240|4.49|2015-02-16 07:04:00|80.995508130988839|4|3338397021|121|35.449819467189094|0|40|741|-80.780702|87|35.318911|"NFS-3""- 8"" FOLIAGE"|0.0|9|"4"" IVY ASSORTMENT    ED"|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|35.466476270328783|00033383970219|FLORAL|FLORAL|-80.995484|80.995486287843732|167|1
35.444064|13b3e789cde8be360a67fcd6f5ed5d5b50b7bc54|1.9|2014-09-14 10:46:00|1.4102725052409182|4||121|0.6186156170875914|0|1|502|-80.995484|64|35.444064|FRESH BANANAS|0.0|4|BANANAS, YELLOW|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|cdf07b7341761b28bc4a44f674db110a8c42f2b5|0.62|2015-01-01 15:19:00|1.4102725052409182|4||121|0.6186156170875914|0|1|502|-80.995484|64|35.444064|FRESH BANANAS|0.0|4|BANANAS, YELLOW|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|8543c7d8afbf423d90b0f16d0d41840ac131564f|0.81|2014-10-05 12:28:00|1.4102725052409182|4||121|0.6186156170875914|0|1|502|-80.995484|64|35.444064|FRESH BANANAS|0.0|4|BANANAS, YELLOW|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|6f1dbc46e59bed45cef1d1fa1a1628ce96105e8b|3.1|2014-12-24 07:06:00|80.995508130988839|4|2920000212|121|35.449819467189094|0|40|149|-80.780702|23|35.318911|WHSE PASTA CORE|0.78|1|MUELLER ELBOW MACARONI|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|35.466476270328783|00029200002133|PASTA|G1 GROCERY|-80.995484|80.995486287843732|167|2
35.444064|dafb56d2ecea88f7362d5057b46be266f5daf3c1|0.87|2015-02-08 10:28:00|1.4102725052409182|4||121|0.6186156170875914|0|1|502|-80.995484|64|35.444064|FRESH BANANAS|0.0|4|BANANAS, YELLOW|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|0d6003438839d5f3fdcdfd74f3ef818d0a57679a|1.23|2015-01-04 12:20:00|1.4102725052409182|4||121|0.6186156170875914|0|1|502|-80.995484|64|35.444064|FRESH BANANAS|0.0|4|BANANAS, YELLOW|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|6a295f8af9b81c270ee1dd593335c9e72835194e|1.56|2014-09-21 11:46:00|1.4102725052409182|4||121|0.6186156170875914|0|1|502|-80.995484|64|35.444064|FRESH BANANAS|0.0|4|BANANAS, YELLOW|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|b7551a6b4df9cffc8e0699cacb6525357e2fef83|10.78|2014-11-07 16:20:00|1.4102725052409182|4|5543762275|121|0.6186156170875914|0|1|719|-80.995484|10|35.444064|NFS-COFFEE FILTERS|2.69|1|MELITTA #4 BROWN COFFEE FILTER|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|0.61833652052202714|00055437624602|COFFEE|G1 GROCERY|-80.995484|1.413637875046387|121|2
35.444064|099911ff2d456627ca716b9551af6055e72472fc|9.99|2014-10-19 11:51:00|1.4102725052409182|4|7818508540|121|0.6186156170875914|0|1|353|-80.995484|110|35.444064|FROZEN CASE MEAT|0.0|19|MRS. BUDD'S WHITE CHICKEN PIE|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|0.61833652052202714|00078185085402|FROZEN CASE MEAT|CASE READY MEATS|-80.995484|1.413637875046387|121|1
35.444064|daa850c1117d0a5b48e1c4150388fcd97aa0bede|16.59|2014-12-06 17:53:00|1.4102725052409182|4|20597500000|121|0.6186156170875914|0|1|1822|-80.995484|410|35.444064|BH CHICKEN|0.0|6|BOARS HEAD BLAZIN BUFFALO CHKN|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|0.61833652052202714|00205975000004|BH MEAT|DELI|-80.995484|1.413637875046387|121|1
35.444064|57b223352f81a6776f4b11a42fe3d33843cb929b|4.0|2015-02-04 07:06:00|80.995508130988839|4|87126000501|121|35.449819467189094|0|40|1165|-80.780702|87|35.318911|NFS-FRESH CONSUMER BUNCH|0.0|9|BUNCH- MINI CARNATION|d89e6e5ff5c1eee89177c8d77412b8fceee72239|0.3976889046626061|35.466476270328783|00871260005018|FLORAL|FLORAL|-80.995484|80.995486287843732|167|1
35.03469|6ed36b0bfb09eb8dac6821aaeee92f5736224d36|3.0|2014-12-04 14:56:00|1.4132775322775095|4|7203660080|82|0.6114706929155321|0|58|1268|-80.97058|54|35.03469|BAGELS AND MUFFINS|0.5|3|HT PIE CRUST|d99fceb7649d71b82ea1dc1b061e8dd3a2b46bf6|1.0062698086776272|0.61177642288969325|00072036600806|DOUGH PRODUCTS|DAIRY|-80.97058|1.4132032182494703|82|1
35.03469|c4501c58956ec5a6e232be8dc4d07c68d1621473|4.99|2015-02-25 19:02:00|1.4132775322775095|4|1780015039|82|0.6114706929155321|0|58|152|-80.97058|24|35.03469|NFS-CAT FOOD DRY|1.0|1|KIT N' KABOODLE ESSENTIALS|d99fceb7649d71b82ea1dc1b061e8dd3a2b46bf6|1.0062698086776272|0.61177642288969325|00017800148849|PET FOOD/SUPPLIES|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|e547fe055425debe64d66b6904186590a855c87b|2.99|2015-01-18 13:38:00|1.4132775322775095|4|7073400003|82|0.6114706929155321|0|58|230|-80.97058|37|35.03469|HERBAL TEA|0.49|1|CELESTIAL SLEEPYTIME|d99fceb7649d71b82ea1dc1b061e8dd3a2b46bf6|1.0062698086776272|0.61177642288969325|00070734000034|TEA|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|ca1c1b30447f779e8a2b1d24899ef741db9ff84d|9.99|2015-02-13 13:09:00|80.970593795509558|4|7674007012|82|35.04925302405384|0|4|62|-80.994596|7|35.061685|SPECIALTY BAR/BOX CHOCOLATE|5.0|1|WHITMAN SAMPLER BOX PP9.99|d99fceb7649d71b82ea1dc1b061e8dd3a2b46bf6|1.0062698086776272|35.073829668338668|00076740070122|CANDY|G1 GROCERY|-80.97058|80.970583071385605|475|1
35.03469|d5b353733fac6fe93cfb6e67d6f117ff1487da5e|11.99|2015-03-01 20:19:00|1.4132775322775095|4|8520000098|82|0.6114706929155321|0|58|9946|-80.97058|886|35.03469|NFS-PREM-BLUSH|0.0|13|SUTTER HOME PINK MOSCATO 1.5L|d99fceb7649d71b82ea1dc1b061e8dd3a2b46bf6|1.0062698086776272|0.61177642288969325|00085200000982|PREMIUM ($8-$10.99)|WINE|-80.97058|1.4132032182494703|82|1
35.03469|5ebfe4a58db62bbe7437f52765f898f694b6435f|1.99|2015-01-11 17:04:00|1.4132775322775095|4|7203648011|82|0.6114706929155321|0|58|274|-80.97058|44|35.03469|ICE|0.0|5|HT BAGGED ICE 10LB (456)|d99fceb7649d71b82ea1dc1b061e8dd3a2b46bf6|1.0062698086776272|0.61177642288969325|00000000004560|ICE|FROZEN|-80.97058|1.4132032182494703|82|1
35.03469|b5f2720d5262bac565d8a750afc99833622b2f44|5.69|2014-10-22 15:45:00|80.970593795509558|4|7756725423|82|35.04925302405384|0|4|252|-80.994596|45|35.061685|PREMIUM ICE CREAM|1.31|5|BREYERS NATURAL VANILLA I/C|d99fceb7649d71b82ea1dc1b061e8dd3a2b46bf6|1.0062698086776272|35.073829668338668|00077567254238|ICE CREAM|FROZEN|-80.97058|80.970583071385605|475|1
35.03469|e1b3adeec3afda1a90e87454c583d21efe6dcc98|2.99|2014-09-18 19:19:00|1.4132775322775095|4|7203698567|82|0.6114706929155321|0|58|199|-80.97058|31|35.03469|DIPS & SALSAS|0.49|1|HT FRENCH ONION DIP|d99fceb7649d71b82ea1dc1b061e8dd3a2b46bf6|1.0062698086776272|0.61177642288969325|00072036985651|SNACKS|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|4ea7de17378ed7a6708471df4bd042749668ca5e|2.99|2015-02-19 14:14:00|1.4132775322775095|4|31284313105|82|0.6114706929155321|0|58|4308|-80.97058|1205|35.03469|ASPIRIN|0.0|17|ASPIRIN REGIMEN BAYER 06132|d99fceb7649d71b82ea1dc1b061e8dd3a2b46bf6|1.0062698086776272|0.61177642288969325|00312843061323|PAIN RELIEF|HBC|-80.97058|1.4132032182494703|82|1
35.297134|9782c6e460caef8a15ad1f7b9856bf5b032c96c7|5.49|2015-02-14 20:12:00|80.728244613218536|4|1037418019|258|35.308582349913806|0|5|1673|-80.66939|383|35.28326|PASTRY CASE CAKES|0.0|14|NO SUGAR ADDED CHEESECAKE|d9c3e0fe0eb209f552f772ed45d283e2e44c182c|0.791053343304979|35.296297200616316|00010374180192|PASTRY CASE|BAKERY|-80.737839|80.737841343256775|46|1
35.297134|523ac5379a2cc0203c799354cd48458dbbc39cd1|40.510000000000005|2014-11-08 12:33:00|80.728244613218536|4|20140400000|258|35.308582336504948|0|5|296|-80.662946|49|35.412407|RANCHER BEEF|3.75|2|BEEF LOIN NY STRIP STEAK BNLS|d9c3e0fe0eb209f552f772ed45d283e2e44c182c|0.791053343304979|35.296297200616316|00201404000003|BEEF|MEAT|-80.737839|80.737860597598825|68|5
35.297134|97896e8d3263f3e8540d8e5b1288b50e266c2cd0|0.97|2015-03-01 13:15:00|80.728244613218536|4|7203671102|258|35.308582349913806|0|5|1025|-80.66939|162|35.28326|WHITE|0.0|7|HT OLD FASHIONED BREAD|d9c3e0fe0eb209f552f772ed45d283e2e44c182c|0.791053343304979|35.296297200616316|00072036711021|SLICED BREAD|COMMERCIAL BAKERY|-80.737839|80.737841343256775|46|1
35.23102|f46a415c1ff77d21802941d0c50558bb6fedecad|2.69|2014-09-29 18:32:00|80.843809562956082|4|3663202720|205|35.247129259498287|0|37|688|-80.844274|61|35.204336|LIGHT|0.69|3|DANNON L&F BLUEBERRY|dff16621afbfa48d91fec6becb5a814d0317d7a1|1.1131109723700134|35.255745041786184|00036632027238|YOGURT|DAIRY|-80.8438|80.843805514634255|61|1
35.23102|0500a3b336846b637bdaca9ce0d5e8e656f7b305|3.59|2015-02-14 18:32:00|80.843809562956082|4|7027200216|205|35.247129259498287|0|37|1132|-80.844274|55|35.204336|EGGS SUBSTITUTES|0.4|3|EGGBEATER CARTON|dff16621afbfa48d91fec6becb5a814d0317d7a1|1.1131109723700134|35.255745041786184|00070272002163|EGGS FRESH|DAIRY|-80.8438|80.843805514634255|61|1
35.23102|4e4225ccce73904dd60069ab26625c6d99ec8dea|6.98|2015-02-07 18:14:00|80.843809562956082|4|3600038587|205|35.247129259498287|0|37|426|-80.844274|72|35.204336|NFS-PAPER TOWELS|0.98|1|KLEENEX HAND TOWEL WHITE|dff16621afbfa48d91fec6becb5a814d0317d7a1|1.1131109723700134|35.255745041786184|00036000385878|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.8438|80.843805514634255|61|2
35.23102|a075110f24260baf36df80cc862549c735386b09|3.99|2014-09-19 16:52:00|80.843809562956082|4|4973309101|205|35.247129259498287|0|37|76|-80.844274|11|35.204336|MEAT SAUCES|1.0|1|ECHOLULA CHIPOTLE SAUCE|dff16621afbfa48d91fec6becb5a814d0317d7a1|1.1131109723700134|35.255745041786184|00049733830119|CONDIMENTS|G1 GROCERY|-80.8438|80.843805514634255|61|1
35.23102|3124b1002287bc8b174b93266c448018458a037a|0.7|2015-01-09 15:18:00|80.843809562956082|4||205|35.247129259498287|0|37|522|-80.844274|64|35.204336|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|dff16621afbfa48d91fec6becb5a814d0317d7a1|1.1131109723700134|35.255745041786184|00204664000004|FRESH PRODUCE|PRODUCE|-80.8438|80.843805514634255|61|1
35.23102|037ae51fffb283b09547aee7bf86dc06d7065534|4.47|2014-09-25 18:54:00|80.843809562956082|4||205|35.247129259498287|0|37|561|-80.844274|64|35.204336|FR PROD ORGANIC PRODUCE|0.7|4|COO ORG GREEN ONIONS|dff16621afbfa48d91fec6becb5a814d0317d7a1|1.1131109723700134|35.255745041786184|00294068000007|FRESH PRODUCE|PRODUCE|-80.8438|80.843805514634255|61|3
35.23102|d179d6922bf86238733f9ccf896820ab5470ed2f|2.19|2015-01-31 15:39:00|80.843809562956082|4|7675324446|205|35.247129259498287|0|37|5900|-80.844274|1538|35.204336|SKEWERS|0.0|18|"(PLR) BAMBOO SKEWERS 4"" 30CT"|dff16621afbfa48d91fec6becb5a814d0317d7a1|1.1131109723700134|35.255745041786184|00076753244466|KITCHEN GADGETS|GM|-80.8438|80.843805514634255|61|1
35.323246|361aa1d6d20e0fe39f4a71647253a854e64bbef6|1.49|2014-12-03 11:57:00|80.945255278477163|3|2840002819|166|35.379456702527264|0|13|206|-80.86175|31|35.40953|FRONT END SNACKS|0.0|1|LAYS BBQ|e06b21d571a3a1c81a2a5604eba09f333ef4463e|3.8840269541479318|35.37387923947206|00028400025904|SNACKS|G1 GROCERY|-80.945176|80.945263821754935|209|1
35.323246|77602dff7a203666223e2fd298380100a1d7c6b4|1.49|2014-10-03 11:37:00|80.945255278477163|3|2840002819|166|35.379456702527264|0|13|206|-80.86175|31|35.40953|FRONT END SNACKS|0.0|1|LAYS BBQ|e06b21d571a3a1c81a2a5604eba09f333ef4463e|3.8840269541479318|35.37387923947206|00028400025904|SNACKS|G1 GROCERY|-80.945176|80.945263821754935|209|1
35.323246|6ca2534f072548bc451ecd447037c845c61f002d|1.49|2014-11-18 11:28:00|80.945255278477163|3|2840002819|166|35.379456702527264|0|13|206|-80.86175|31|35.40953|FRONT END SNACKS|0.0|1|LAYS BBQ|e06b21d571a3a1c81a2a5604eba09f333ef4463e|3.8840269541479318|35.37387923947206|00028400025904|SNACKS|G1 GROCERY|-80.945176|80.945263821754935|209|1
35.323246|765587c4a8dcf5fd58108a00a670d4e77b6773f7|1.49|2014-10-21 12:20:00|80.945255278477163|3|2840002819|166|35.379456702527264|0|13|206|-80.86175|31|35.40953|FRONT END SNACKS|0.0|1|LAYS BBQ|e06b21d571a3a1c81a2a5604eba09f333ef4463e|3.8840269541479318|35.37387923947206|00028400025904|SNACKS|G1 GROCERY|-80.945176|80.945263821754935|209|1
35.323246|f018835fd7d8ee95f19acc83c7d0137a64cdae70|1.89|2014-10-01 10:52:00|80.945255278477163|3|8390000575|166|35.379456702527264|0|13|99|-80.86175|32|35.40953|LIQUID TEA|0.2|1|GOLD PEAK DIET|e06b21d571a3a1c81a2a5604eba09f333ef4463e|3.8840269541479318|35.37387923947206|00083900005764|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.945176|80.945263821754935|209|1
35.323246|350e62efb021c646926c4936cf4a63ce25464580|8.58|2014-11-29 10:11:00|80.945255278477163|3|1115605450|166|35.379456702527264|0|13|233|-80.86175|37|35.40953|BLACK TEA|0.0|1|TETLEY TEA BRITISH BLEND 80CT|e06b21d571a3a1c81a2a5604eba09f333ef4463e|3.8840269541479318|35.37387923947206|00011156054502|TEA|G1 GROCERY|-80.945176|80.945263821754935|209|2
35.323246|d1fa5c08bd230b2eb4f09a989998a8c83e77753b|4.29|2015-03-06 12:04:00|80.945255278477163|3|1115605450|166|35.379456702527264|0|13|233|-80.86175|37|35.40953|BLACK TEA|0.0|1|TETLEY TEA BRITISH BLEND 80CT|e06b21d571a3a1c81a2a5604eba09f333ef4463e|3.8840269541479318|35.37387923947206|00011156054502|TEA|G1 GROCERY|-80.945176|80.945263821754935|209|1
35.323246|199c18dbe2bd24b5586a0d62b2372e22b6ff0ba4|2.0|2015-01-01 12:59:00|80.945255278477163|3|4300000953|166|35.379456702527264|0|13|272|-80.86175|307|35.40953|TOPPINGS FROZEN|1.01|5|COOL WHIP WHIPPED TOPPING|e06b21d571a3a1c81a2a5604eba09f333ef4463e|3.8840269541479318|35.37387923947206|00043000009536|DESSERTS FROZEN|FROZEN|-80.945176|80.945263821754935|209|1
35.323246|519c77149db2bd9575c4b3675197597d3d6b299e|4.99|2014-11-20 07:26:00|80.945255278477163|3|7144830025|166|35.379456702527264|0|13|2021|-80.86175|505|35.40953|FRESH CHEESE|1.49|6|ALOUETTE GARLIC & HERB|e06b21d571a3a1c81a2a5604eba09f333ef4463e|3.8840269541479318|35.37387923947206|00071448300144|SPECIALTY CHEESE|DELI|-80.945176|80.945263821754935|209|1
35.323246|acb5548d1c072b20fbc7c6b5a15e8ba36272bf0e|2.65|2014-11-24 14:30:00|80.945255278477163|3|4119640471|166|35.379456702527264|0|13|1201|-80.86175|33|35.40953|RTS CANNED|0.65|1|PROG LIGHT BEEF POT ROAST|e06b21d571a3a1c81a2a5604eba09f333ef4463e|3.8840269541479318|35.37387923947206|00041196404814|SOUP|G1 GROCERY|-80.945176|80.945263821754935|209|1
35.323246|5c60bdf09607de99286c3e4262ff9b0ba048adbd|4.0|2015-01-22 12:27:00|80.945255278477163|3|7047043332|166|35.379456702527264|0|13|685|-80.86175|61|35.40953|GREEK|1.0|3|YOPLAIT GREEK 100 APPLE PIE|e06b21d571a3a1c81a2a5604eba09f333ef4463e|3.8840269541479318|35.37387923947206|00070470476384|YOGURT|DAIRY|-80.945176|80.945263821754935|209|3
35.323246|b99febadb7a0f3d476800c9c865276507ef3206b|3.79|2014-09-13 13:44:00|80.945255278477163|3|7020055044|166|35.379456702527264|0|13|580|-80.86175|136|35.40953|OTHER MERCH DRESSINGS|0.0|4|MARZ SIMPLY CAESAR DRESSING|e06b21d571a3a1c81a2a5604eba09f333ef4463e|3.8840269541479318|35.37387923947206|00070200550469|OTHER MERCHANDISE|PRODUCE|-80.945176|80.945263821754935|209|1
35.323246|7bf2f518c6b759f667913e399d7bb99018b0096c|1.0|2014-09-23 12:33:00|80.945255278477163|3|61300873089|166|35.379456686978969|0|13|99|-80.8955|32|35.4437|LIQUID TEA|0.0|1|PP ARIZONA ARNOLD PALMER|e06b21d571a3a1c81a2a5604eba09f333ef4463e|3.8840269541479318|35.37387923947206|00613008730895|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.945176|80.945277687001536|272|1
35.323246|f9e280bc0206f1151ae4f9bb73e63fb927907b58|2.99|2014-12-23 14:11:00|80.945255278477163|3|61300873513|166|35.379456686978969|0|13|99|-80.8955|32|35.4437|LIQUID TEA|0.0|1|ARNOLD PALMER ZERO HALF&HALF|e06b21d571a3a1c81a2a5604eba09f333ef4463e|3.8840269541479318|35.37387923947206|00613008730444|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.945176|80.945277687001536|272|1
35.323246|f6a895d09bab175cfd5c8f5cf031d05548f88ec3|1.0|2014-09-26 12:19:00|80.945255278477163|3|61300872573|166|35.379456686978969|0|13|99|-80.8955|32|35.4437|LIQUID TEA|0.0|1|PP ARIZONA SWEET TEA|e06b21d571a3a1c81a2a5604eba09f333ef4463e|3.8840269541479318|35.37387923947206|00613008725730|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.945176|80.945277687001536|272|1
35.323246|3953f041b6ef5334b38c784d6c9764c364278721|4.29|2014-10-17 09:29:00|80.945255278477163|3|70897111891|166|35.379456702527264|0|13|1703|-80.86175|387|35.40953|SEASONAL COOKIES|1.79|14|HARVEST ORANGE FRSTD CHOC COOK|e06b21d571a3a1c81a2a5604eba09f333ef4463e|3.8840269541479318|35.37387923947206|00708971118914|COOKIES|BAKERY|-80.945176|80.945263821754935|209|1
35.323246|fd222edacd2ed0f58ec4735b35e2724716fca0f7|4.99|2015-02-23 07:57:00|80.945255278477163|3|1111018700|166|35.379456702527264|0|13|1647|-80.86175|379|35.40953|PACKAGED MUFFINS|1.02|14|FFM 4 CT BLUEBERRY MUFFIN|e06b21d571a3a1c81a2a5604eba09f333ef4463e|3.8840269541479318|35.37387923947206|00011110187000|MUFFINS|BAKERY|-80.945176|80.945263821754935|209|1
35.323246|487212da0ce76a130c93d3081d51be796d24c871|49.78|2014-11-22 13:15:00|80.945255278477163|3|20000700000|166|35.379456702527264|0|13|974|-80.86175|201|35.40953|FRESH TURKEY|14.58|2|BUTTERBALL FRSH TOM TRKY 16-22|e06b21d571a3a1c81a2a5604eba09f333ef4463e|3.8840269541479318|35.37387923947206|00200007000007|POULTRY|MEAT|-80.945176|80.945263821754935|209|1
35.323246|4abfe7a54eae80b11f8445e7fb120bcaacbd2bc4|3.49|2015-01-07 12:53:00|1.4102725052409182|4|7797503405|166|0.6165069451919168|0|1|202|-80.945176|31|35.323246|PRETZELS|0.0|1|SNYDERS RODS PRETZEL|e1f0574196fc0f90390a38ff930088c6b2cb706b|4.438685104811772|0.61833652052202714|00077975034064|SNACKS|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|6e04a0b637a79079ff695a162ac8bb7b7e4ea4dd|3.89|2015-02-03 20:27:00|1.4102725052409182|4|7457000400|166|0.6165069451919168|0|1|275|-80.945176|45|35.323246|SUPER PREMIUM ICE CREAM|0.0|5|H DAZS WHITE CHOC RASP TRF|e1f0574196fc0f90390a38ff930088c6b2cb706b|4.438685104811772|0.61833652052202714|00074570650309|ICE CREAM|FROZEN|-80.945176|1.4127598348062935|166|1
35.323246|8cf69af1e520e9d75b8823b6a0c982307e242401|3.99|2014-12-08 12:38:00|1.4102725052409182|4|7457000400|166|0.6165069451919168|0|1|275|-80.945176|45|35.323246|SUPER PREMIUM ICE CREAM|0.0|5|H DAZS WHITE CHOC RASP TRF|e1f0574196fc0f90390a38ff930088c6b2cb706b|4.438685104811772|0.61833652052202714|00074570650309|ICE CREAM|FROZEN|-80.945176|1.4127598348062935|166|1
35.323246|a414eeef0ee3920d55505c471e3f4b8da039db88|5.18|2014-09-15 13:50:00|1.4102725052409182|4|2800021010|166|0.6165069451919168|0|1|16|-80.945176|3|35.323246|BAKING CHOCOLATE/CHIPS/MORSELS|0.0|1|NESTLE SEMISWEET MORSELS|e1f0574196fc0f90390a38ff930088c6b2cb706b|4.438685104811772|0.61833652052202714|00028000215804|BAKING SUPPLIES|G1 GROCERY|-80.945176|1.4127598348062935|166|2
35.323246|8a2b8a7c69e51c19aa6acd2be7be21a7c050b6b4|2.35|2014-09-10 13:49:00|1.4102725052409182|4|4112907700|166|0.6165069451919168|0|1|1219|-80.945176|275|35.323246|PASTA SC CORE|0.0|1|CLASSICO SC SPICY RED PEPPER|e1f0574196fc0f90390a38ff930088c6b2cb706b|4.438685104811772|0.61833652052202714|00041129077429|PASTA SAUCES|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|6d0f4cf883095b4382ab0737a296852a456ae5b5|2.45|2014-10-03 10:18:00|1.4102725052409182|4|7203663217|166|0.6165069451919168|0|1|330|-80.945176|55|35.323246|EGGS|0.0|3|HT GRADE A LARGE EGGS 18 CT|e1f0574196fc0f90390a38ff930088c6b2cb706b|4.438685104811772|0.61833652052202714|00072036632173|EGGS FRESH|DAIRY|-80.945176|1.4127598348062935|166|1
35.323246|099249e5ba9160520b016c87408889af3aa7a4b4|2.0|2015-01-06 13:18:00|1.4102725052409182|4||166|0.6165069451919168|0|1|511|-80.945176|64|35.323246|FRESH AVOCADOS|0.11|4|AVOCADOS, HASS XL 36CT|e1f0574196fc0f90390a38ff930088c6b2cb706b|4.438685104811772|0.61833652052202714|00204770000004|FRESH PRODUCE|PRODUCE|-80.945176|1.4127598348062935|166|1
35.323246|373caaef01121eb459238664c064f7d3203486fc|4.0|2015-01-13 17:04:00|1.4102725052409182|4||166|0.6165069451919168|0|1|511|-80.945176|64|35.323246|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|e1f0574196fc0f90390a38ff930088c6b2cb706b|4.438685104811772|0.61833652052202714|00204770000004|FRESH PRODUCE|PRODUCE|-80.945176|1.4127598348062935|166|2
35.323246|09a3f839aa87efa33a4a214dfe28dba8d9206c9d|7.99|2015-01-21 17:13:00|1.4102725052409182|4|20250700000|166|0.6165069451919168|0|1|642|-80.945176|49|35.323246|NATURAL/ORGANIC BEEF|1.0|2|NATURAL 90% LEAN GROUND BEEF|e1f0574196fc0f90390a38ff930088c6b2cb706b|4.438685104811772|0.61833652052202714|00202507000006|BEEF|MEAT|-80.945176|1.4127598348062935|166|1
35.323246|27fb6a7d4ba2d014bea2b3be274173e70555fa2b|1.99|2014-12-08 13:17:00|1.4102725052409182|4|7053807511|166|0.6165069451919168|0|1|727|-80.945176|7|35.323246|SEASONAL CANDY-SINGLE FAC|0.32|1|I/O(C15)BOB MINI CANE 40CT|e1f0574196fc0f90390a38ff930088c6b2cb706b|4.438685104811772|0.61833652052202714|00070538075115|CANDY|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|b863c5e004f485ce7d0b9a95aa648735567c4ee0|4.55|2015-02-24 10:29:00|1.4102725052409182|4||166|0.6165069451919168|0|1|529|-80.945176|64|35.323246|FRESH ASPARAGUS|2.51|4|GREEN  ASPARAGUS|e1f0574196fc0f90390a38ff930088c6b2cb706b|4.438685104811772|0.61833652052202714|00204080000008|FRESH PRODUCE|PRODUCE|-80.945176|1.4127598348062935|166|1
35.323246|837a9b55d517f0013a3ed4d845dbec642ff52c0a|5.99|2014-11-24 11:20:00|1.4102725052409182|4|72037950126|166|0.6165069451919168|0|1|117|-80.945176|17|35.323246|DRIED REMAINING FRUIT|1.0|1|MADE IN NAT ORG DRY PINEAPPLE|e1f0574196fc0f90390a38ff930088c6b2cb706b|4.438685104811772|0.61833652052202714|00720379501266|FRUIT-DRIED|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|a59762fceeb9ec597bfc34c7c0a8696e65eebab5|5.99|2014-11-30 20:29:00|1.4102725052409182|4|72037950126|166|0.6165069451919168|0|1|117|-80.945176|17|35.323246|DRIED REMAINING FRUIT|1.0|1|MADE IN NAT ORG DRY PINEAPPLE|e1f0574196fc0f90390a38ff930088c6b2cb706b|4.438685104811772|0.61833652052202714|00720379501266|FRUIT-DRIED|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|ac527b42fbb94fcbf65ac479934d88c2288d24ee|19.99|2014-10-03 10:12:00|1.4102725052409182|4|4116743104|166|0.6165069451919168|0|1|4234|-80.945176|1200|35.323246|PSE SOLID DOSE|0.0|17|(PSE)ALLEGRA D 12 HR E/R CAPS|e1f0574196fc0f90390a38ff930088c6b2cb706b|4.438685104811772|0.61833652052202714|00041167431047|COUGH/COLD/SINUS|HBC|-80.945176|1.4127598348062935|166|1
35.323246|c6344c85b6127191b12df81b37c2440b77de21dc|0.5|2015-01-28 11:41:00|1.4102725052409182|4||166|0.6165069451919168|0|1|543|-80.945176|64|35.323246|FRESH GARLIC|0.0|4|COO GARLIC, WHITE, BULK|e1f0574196fc0f90390a38ff930088c6b2cb706b|4.438685104811772|0.61833652052202714|00204608000008|FRESH PRODUCE|PRODUCE|-80.945176|1.4127598348062935|166|1
35.323246|c901b0549159096223a118fec88e61cd1173c2c9|3.0|2014-11-22 21:55:00|1.4102725052409182|4|7203670492|166|0.6165069451919168|0|1|117|-80.945176|17|35.323246|DRIED REMAINING FRUIT|0.0|1|HT YOGURT RAISINS|e1f0574196fc0f90390a38ff930088c6b2cb706b|4.438685104811772|0.61833652052202714|00072036704924|FRUIT-DRIED|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|aa929f19d3a3a4026e7c35130dee5a21f454a382|3.0|2014-12-20 16:48:00|1.4102725052409182|4|7203670492|166|0.6165069451919168|0|1|117|-80.945176|17|35.323246|DRIED REMAINING FRUIT|0.0|1|HT YOGURT RAISINS|e1f0574196fc0f90390a38ff930088c6b2cb706b|4.438685104811772|0.61833652052202714|00072036704924|FRUIT-DRIED|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|0d0c552a0af3b9d0fdbfb2b4aaa3bb2f5e6bc13e|3.75|2014-11-24 11:19:00|1.4102725052409182|4|4470000063|166|0.6165069451919168|0|1|359|-80.945176|101|35.323246|MEAT WIENERS|0.0|19|OSCAR MAYER BUNLENGTH TURKEY|e1f0574196fc0f90390a38ff930088c6b2cb706b|4.438685104811772|0.61833652052202714|00071871544641|WIENERS|CASE READY MEATS|-80.945176|1.4127598348062935|166|1
35.43259|cb9ee5b0144e89ef860e6c1ad3d621e7eeb1753f|4.99|2014-12-09 13:28:00|1.4057311447477159|4|7203688117|202|0.6184153580092175|0|52|583|-80.605588|136|35.43259|NUTS|0.0|4|HT FILBERTS IN SHELL 1LB|e5da976040773545056c57c5ddcaadbe97ed7951|9.073372822842245|0.6209993146566879|00072036881175|OTHER MERCHANDISE|PRODUCE|-80.605588|1.406832906106031|202|1
35.43259|d873de9ca3e75096c88640d5eb512cd690d6f07f|4.99|2014-11-24 13:43:00|1.4057311447477159|4|7203688117|202|0.6184153580092175|0|52|583|-80.605588|136|35.43259|NUTS|0.0|4|HT FILBERTS IN SHELL 1LB|e5da976040773545056c57c5ddcaadbe97ed7951|9.073372822842245|0.6209993146566879|00072036881175|OTHER MERCHANDISE|PRODUCE|-80.605588|1.406832906106031|202|1
35.43259|0f3b72b03f55d4379c282069c435d9d0c59a82fe|3.99|2014-12-24 17:57:00|80.606823361882718|4|7835470843|202|35.563902430097258|0|57|317|-80.662946|52|35.412407|CHUNK AND BAR CHEESE|1.49|3|CABOT SERIOUSLY SHARP YELLOW|e5da976040773545056c57c5ddcaadbe97ed7951|9.073372822842245|35.500309569604553|00078354717288|CHEESE|DAIRY|-80.605588|80.605664151521935|68|1
35.43259|c6355b3a9aab36494ddd62459914fbf80faff05e|2.99|2015-02-19 16:22:00|1.4057311447477159|4|7203670267|202|0.6184153580092175|0|52|176|-80.605588|72|35.43259|NFS-DISPOSE CUPS|0.0|1|YH PLASTIC CUPS 9 OZ|e5da976040773545056c57c5ddcaadbe97ed7951|9.073372822842245|0.6209993146566879|00072036702678|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.605588|1.406832906106031|202|1
35.43259|7ae90197e051428441ac851c80095bd280c6a8c2|5.58|2015-02-19 19:35:00|1.4057311447477159|4|7203698417|202|0.6184153580092175|0|52|423|-80.605588|72|35.43259|NFS-DISPOSE PLATES/BOWLS|0.0|1|"YH 7"" ELEGWARE OCTAGONAL PLAT"|e5da976040773545056c57c5ddcaadbe97ed7951|9.073372822842245|0.6209993146566879|00072036984173|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.605588|1.406832906106031|202|2
35.059823|f3523c07c21834abb46fa46ca02c4c784194fee3|1.49|2014-12-01 17:56:00|1.4091206135396188|3|3400000727|66|0.6119093465164359|0|47|727|-80.816172|7|35.059823|SEASONAL CANDY-SINGLE FAC|0.75|1|I/O(C14)HRSHY CHOC SANTA|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00034000007271|CANDY|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|ed3c9c6192aeda48329f62992df0bb645bcf9250|3.39|2015-03-08 21:47:00|1.4091206135396188|3|3800031829|66|0.6119093465164359|0|47|74|-80.816172|9|35.059823|RTE CEREAL ALL FAMILY|0.0|1|KELL MIN WH FROST RAISIN|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00038000102301|CEREAL|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|6f68006227bca741c5f3483cd7f4f8ef5e863df8|3.39|2014-10-26 19:27:00|1.4091206135396188|3|3800031829|66|0.6119093465164359|0|47|74|-80.816172|9|35.059823|RTE CEREAL ALL FAMILY|1.7|1|KELL MIN WH FROST RAISIN|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00038000102301|CEREAL|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|cd776aee819e02e8e02948946e6fb2a788eb2af9|6.78|2015-01-26 19:01:00|1.4091206135396188|3|3800031829|66|0.6119093465164359|0|47|74|-80.816172|9|35.059823|RTE CEREAL ALL FAMILY|1.78|1|KELL MIN WH FROST RAISIN|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00038000102301|CEREAL|G1 GROCERY|-80.816172|1.4105082902580508|66|2
35.059823|45534cf8baa5fa3812074b59427aeb022c9a4870|3.39|2015-01-03 21:40:00|1.4091206135396188|3|3800031829|66|0.6119093465164359|0|47|74|-80.816172|9|35.059823|RTE CEREAL ALL FAMILY|0.0|1|KELL MIN WH FROST RAISIN|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00038000102301|CEREAL|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|f94fa52cc10e737abf6a8878c5a74fda46ee1f62|3.39|2014-12-22 16:25:00|1.4091206135396188|3|3800031829|66|0.6119093465164359|0|47|74|-80.816172|9|35.059823|RTE CEREAL ALL FAMILY|0.0|1|KELL MIN WH FROST RAISIN|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00038000102301|CEREAL|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|473e814efc01481ca505d3c617fa03dd8212d643|3.39|2014-12-30 11:38:00|1.4091206135396188|3|3800031829|66|0.6119093465164359|0|47|74|-80.816172|9|35.059823|RTE CEREAL ALL FAMILY|0.0|1|KELL MIN WH FROST RAISIN|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00038000102301|CEREAL|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|f1c3cbbb4781f0e18ace3245dc80b76d3bff0848|3.39|2014-11-23 18:47:00|1.4091206135396188|3|3800031829|66|0.6119093465164359|0|47|74|-80.816172|9|35.059823|RTE CEREAL ALL FAMILY|0.0|1|KELL MIN WH FROST RAISIN|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00038000102301|CEREAL|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|1d34e7e69a8e6130d211f4108b7a347bdd414202|3.39|2015-01-10 21:38:00|1.4091206135396188|3|3800031829|66|0.6119093465164359|0|47|74|-80.816172|9|35.059823|RTE CEREAL ALL FAMILY|0.0|1|KELL MIN WH FROST RAISIN|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00038000102301|CEREAL|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|41cbe76f146ba51d62f6bd6e6cd741af31eef079|6.78|2015-02-23 18:48:00|1.4091206135396188|3|3800031829|66|0.6119093465164359|0|47|74|-80.816172|9|35.059823|RTE CEREAL ALL FAMILY|0.89|1|KELL MIN WH FROST RAISIN|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00038000102301|CEREAL|G1 GROCERY|-80.816172|1.4105082902580508|66|2
35.059823|81e753a0023fd954944e07b394244ff994349372|1.97|2015-03-02 19:00:00|1.4091206135396188|3|7203633023|66|0.6119093465164359|0|47|200|-80.816172|31|35.059823|MICROWAVE POPCORN|0.0|1|HT POPCORN - BAGGED  2 LB|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00072036330239|SNACKS|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|ff547e7c07ae82226bfaa44eb3de81b57ad06d0d|3.69|2015-01-15 17:13:00|1.4091206135396188|3|7127928100|66|0.6119093465164359|0|47|555|-80.816172|64|35.059823|PACKAGED SALADS|0.0|4|F.E. VEGGIE LOVERS SALAD|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00071279281001|FRESH PRODUCE|PRODUCE|-80.816172|1.4105082902580508|66|1
35.059823|ceee0c90c6ce428ef7689fbd012a938df4ab850c|3.69|2015-01-31 09:32:00|1.4091206135396188|3|7127928100|66|0.6119093465164359|0|47|555|-80.816172|64|35.059823|PACKAGED SALADS|0.0|4|F.E. VEGGIE LOVERS SALAD|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00071279281001|FRESH PRODUCE|PRODUCE|-80.816172|1.4105082902580508|66|1
35.059823|c997e9c8a755ee314c5107b1ce5d5d5286557fcb|3.69|2015-02-19 12:55:00|1.4091206135396188|3|7127928100|66|0.6119093465164359|0|47|555|-80.816172|64|35.059823|PACKAGED SALADS|0.0|4|F.E. VEGGIE LOVERS SALAD|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00071279281001|FRESH PRODUCE|PRODUCE|-80.816172|1.4105082902580508|66|1
35.059823|e25e86e050d1aee3b374083a1e799d3164239dfe|3.69|2015-01-18 15:31:00|1.4091206135396188|3|7127928100|66|0.6119093465164359|0|47|555|-80.816172|64|35.059823|PACKAGED SALADS|0.0|4|F.E. VEGGIE LOVERS SALAD|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00071279281001|FRESH PRODUCE|PRODUCE|-80.816172|1.4105082902580508|66|1
35.059823|cfa9e566c54419f75b050614fb2c0a3a5c6a531f|3.99|2015-01-11 19:40:00|1.4091206135396188|3|7127927100|66|0.6119093465164359|0|47|555|-80.816172|64|35.059823|PACKAGED SALADS|0.0|4|F.E. BABY SPINACH|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00071279271002|FRESH PRODUCE|PRODUCE|-80.816172|1.4105082902580508|66|1
35.059823|27696173789f53afaf43f5640bb04a82feee6886|3.69|2015-02-03 16:17:00|1.4091206135396188|3|7127928100|66|0.6119093465164359|0|47|555|-80.816172|64|35.059823|PACKAGED SALADS|0.0|4|F.E. VEGGIE LOVERS SALAD|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00071279281001|FRESH PRODUCE|PRODUCE|-80.816172|1.4105082902580508|66|1
35.059823|0cfb4a39772afa50caad4ff8ff16f1b907f20966|3.69|2015-01-05 16:48:00|1.4091206135396188|3|7127928100|66|0.6119093465164359|0|47|555|-80.816172|64|35.059823|PACKAGED SALADS|0.0|4|F.E. VEGGIE LOVERS SALAD|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00071279281001|FRESH PRODUCE|PRODUCE|-80.816172|1.4105082902580508|66|1
35.059823|04d54e7fa755c81008ae7daffc4bba5486e3324d|1.2|2014-11-20 17:10:00|1.4091206135396188|3|2400001738|66|0.6119093465164359|0|47|257|-80.816172|39|35.059823|TOMATOES|0.2|1|DEL MONTE TOMATO CHILI STYLE|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00024000012672|VEGETABLES-CAN/JAR|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|d7a9f213b6c83e7c4c36ba7063bc5d364e488b48|2.29|2014-11-07 16:48:00|1.4091206135396188|3|1800000260|66|0.6119093465164359|0|47|325|-80.816172|54|35.059823|BISCUITS-REFRIGERATED|0.0|3|GRANDS BUTTERMILK BISCUITS|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00018000001828|DOUGH PRODUCTS|DAIRY|-80.816172|1.4105082902580508|66|1
35.059823|74925f31bd33e263caf022cc26e3a951c0be72f1|2.77|2014-11-04 15:43:00|1.4091206135396188|3|3338353030|66|0.6119093465164359|0|47|523|-80.816172|64|35.059823|FRESH POTATOES|0.0|4|RUSSET POTATO 8LB BAG|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00033383530307|FRESH PRODUCE|PRODUCE|-80.816172|1.4105082902580508|66|1
35.059823|4f4d23838fb58d1df85bb03cd5acd88ad4b220fb|4.19|2014-11-26 16:50:00|1.4091206135396188|3|5210007086|66|0.6119093465164359|0|47|217|-80.816172|34|35.059823|EXTRACTS FOOD COLORING|1.26|1|E  MCCORMICK VANILLA EXTRACT|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00052100070865|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|5ee8ece35b8f9c88c8b3a768c9df048862b71361|3.29|2014-09-26 19:12:00|1.4091206135396188|3|7203670548|66|0.6119093465164359|0|47|318|-80.816172|52|35.059823|SHREDDED/GRATED CHEESE|0.0|3|HTT PARMESAN/ROMANO SHRED|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00072036705488|CHEESE|DAIRY|-80.816172|1.4105082902580508|66|1
35.059823|558e8593ac772d1470c9ea069c0f2f645d0f1480|1.79|2015-01-22 18:58:00|1.4091206135396188|3|7142901230|66|0.6119093465164359|0|47|238|-80.816172|38|35.059823|RICE FLAVORED|0.29|1|ZATARAINS RICE SPANISH.|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00071429012271|RICE GRAINS AND BEANS|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|cf5db05e524c0c6cff818c866058a0d95f54103d|1.79|2015-02-26 19:54:00|1.4091206135396188|3|7142901230|66|0.6119093465164359|0|47|238|-80.816172|38|35.059823|RICE FLAVORED|0.29|1|ZATARAINS RICE SPANISH.|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00071429012271|RICE GRAINS AND BEANS|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|57318acfc471ca87e2697b888f80bff5245ff2ff|1.79|2015-03-09 19:01:00|1.4091206135396188|3|7142901230|66|0.6119093465164359|0|47|238|-80.816172|38|35.059823|RICE FLAVORED|0.29|1|ZATARAINS RICE SPANISH.|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00071429012271|RICE GRAINS AND BEANS|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|79d9032b15f843edb925d4c1ad95ee733dc5e3fe|1.25|2015-02-15 21:57:00|1.4091206135396188|3|7203624020|66|0.6119093465164359|0|47|149|-80.816172|23|35.059823|WHSE PASTA CORE|0.25|1|HT PASTA PENNE RIGATE|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00072036240200|PASTA|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|fd84303effebbadd336ee7fe36395004285cb6da|4.49|2015-02-04 18:48:00|1.4091206135396188|3|4812127707|66|0.6119093465164359|0|47|1036|-80.816172|164|35.059823|BREAKFAST BAGELS|2.24|7|THOMAS SEASONAL BAGELS PP|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00048121251000|BREAKFAST|COMMERCIAL BAKERY|-80.816172|1.4105082902580508|66|1
35.059823|54b2aa80da6664fed2fef39aa6155bf4d8f6d12e|4.49|2015-02-10 18:40:00|1.4091206135396188|3|4812127707|66|0.6119093465164359|0|47|1036|-80.816172|164|35.059823|BREAKFAST BAGELS|2.24|7|THOMAS SEASONAL BAGELS PP|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00048121251000|BREAKFAST|COMMERCIAL BAKERY|-80.816172|1.4105082902580508|66|1
35.059823|dcf29a1630663fd427d06af031082a63285de4fb|2.49|2015-01-07 18:13:00|1.4091206135396188|3|2700037882|66|0.6119093465164359|0|47|257|-80.816172|39|35.059823|TOMATOES|0.0|1|HUNTS TOMATO DICED BGO 28|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00027000378908|VEGETABLES-CAN/JAR|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|8b9381cda83915992e2b1716b4029a59478c83eb|7.78|2015-02-06 18:30:00|1.4091206135396188|3|2265530615|66|0.6119093465164359|0|47|487|-80.816172|105|35.059823|PRECOOKED B/FAST SAUSAGE|2.78|19|BUTTERBALL COOKED TURK PATTIES|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00022655306160|BREAKFAST SAUSAGE|CASE READY MEATS|-80.816172|1.4105082902580508|66|2
35.059823|373b61cef46d0678016e3a1782675ade27e70d73|2.69|2014-12-08 18:35:00|1.4091206135396188|3|2700039023|66|0.6119093465164359|0|47|257|-80.816172|39|35.059823|TOMATOES|0.9|1|HUNTS TOMATO SAUCE 29|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00027000390238|VEGETABLES-CAN/JAR|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|10533826d6af93b7f2a3d0a35f95090a6f766c38|3.89|2015-02-11 19:16:00|1.4091206135396188|3|2265530615|66|0.6119093465164359|0|47|487|-80.816172|105|35.059823|PRECOOKED B/FAST SAUSAGE|0.92|19|BUTTERBALL COOKED TURK PATTIES|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00022655306160|BREAKFAST SAUSAGE|CASE READY MEATS|-80.816172|1.4105082902580508|66|1
35.059823|60fc47cdd21fed4644e2673e16299f3e722faf49|3.49|2014-09-23 20:31:00|1.4091206135396188|3|7203688133|66|0.6119093465164359|0|47|556|-80.816172|64|35.059823|PACKAGED VEGETABLES|0.0|4|HT FAJITA MIX|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00072036881335|FRESH PRODUCE|PRODUCE|-80.816172|1.4105082902580508|66|1
35.059823|8a16e880d74f22121ab01ebd9158c14c5cb56b05|3.49|2014-09-13 17:24:00|1.4091206135396188|3|7203688133|66|0.6119093465164359|0|47|556|-80.816172|64|35.059823|PACKAGED VEGETABLES|0.0|4|HT FAJITA MIX|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00072036881335|FRESH PRODUCE|PRODUCE|-80.816172|1.4105082902580508|66|1
35.059823|2eadef3fa8f37c336a1bdf0b414b65c9c9c4b594|9.98|2014-12-13 17:48:00|1.4091206135396188|3|1111018700|66|0.6119093465164359|0|47|1647|-80.816172|379|35.059823|PACKAGED MUFFINS|2.04|14|FFM 4 CT DBL CHOC CHIP MUFFIN|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00011110187024|MUFFINS|BAKERY|-80.816172|1.4105082902580508|66|2
35.059823|feea656189a5c3ffd64a58e98ca211337db1ad82|2.69|2014-10-28 16:09:00|1.4091206135396188|3|70935100013|66|0.6119093465164359|0|47|556|-80.816172|64|35.059823|PACKAGED VEGETABLES|0.69|4|APIO BROCCOLI FLORETS|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00709351000133|FRESH PRODUCE|PRODUCE|-80.816172|1.4105082902580508|66|1
35.059823|1c32254812d41dd572c334a3bfb02b3c004b7296|11.28|2014-12-05 17:46:00|1.4091206135396188|3|20895300000|66|0.6119093465164359|0|47|977|-80.816172|201|35.059823|FRESH HT CHICKEN|0.0|2|HT FRESH BNLS CHICKEN BREAST|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00208953000003|POULTRY|MEAT|-80.816172|1.4105082902580508|66|1
35.059823|057dc5f47508eee664eb3a0c989c5759b3ecaeba|8.98|2015-01-16 18:30:00|1.4091206135396188|3|20895300000|66|0.6119093465164359|0|47|977|-80.816172|201|35.059823|FRESH HT CHICKEN|0.0|2|HT FRESH BNLS CHICKEN BREAST|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00208953000003|POULTRY|MEAT|-80.816172|1.4105082902580508|66|1
35.059823|c617fb95aa1ebd0737b84d4c907ff54b11f9a5d0|9.68|2014-10-14 19:03:00|1.4091206135396188|3|20895300000|66|0.6119093465164359|0|47|977|-80.816172|201|35.059823|FRESH HT CHICKEN|0.0|2|HT FRESH BNLS CHICKEN BREAST|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00208953000003|POULTRY|MEAT|-80.816172|1.4105082902580508|66|1
35.059823|d1e86a46a4d3d9605fb98cc439c072a6471a8040|1.99|2014-10-20 15:52:00|1.4091206135396188|3|4600081101|66|0.6119093465164359|0|47|1213|-80.816172|272|35.059823|HISP DINNERS/SHELLS|0.0|1|OEP SHELL TACO STND STF|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00046000279183|HISPANIC PREP. FOODS|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|89b479e25c019397ab252c78b449a1950649fa7f|0.99|2015-02-12 18:06:00|1.4091206135396188|3|2700038815|66|0.6119093465164359|0|47|257|-80.816172|39|35.059823|TOMATOES|0.19|1|HUNTS TOMATO PASTE BSL GAR ORE|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00027000388235|VEGETABLES-CAN/JAR|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|266e430d4c819ba3b63ed95e044fd46ca0cda01b|3.15|2015-02-24 18:54:00|1.4091206135396188|3|3000001190|66|0.6119093465164359|0|47|60|-80.816172|9|35.059823|HOT CEREAL|0.65|1|QUAKER OATML RSN DATE WALNT|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00030000012406|CEREAL|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|3fef41b22b6a923e00ef90996e6c0bc8d1751b68|2.49|2014-10-15 19:20:00|1.4091206135396188|3|7203690022|66|0.6119093465164359|0|47|1035|-80.816172|163|35.059823|SANDWICH ROLL|0.0|7|HT PREM WHEAT SNDWCH BUN 8CT|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00072036900227|BUNS/ROLLS|COMMERCIAL BAKERY|-80.816172|1.4105082902580508|66|1
35.059823|7d8be3a38f5f418f26c93d536546e2824537087d|1.97|2014-10-06 16:33:00|1.4091206135396188|3|7203614993|66|0.6119093465164359|0|47|105|-80.816172|16|35.059823|FRUIT CUPS AND GELS|0.0|1|HT 4PK FRT CUP MANDARIN NSA|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00072036708052|FRUIT-CAN/JAR|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|0520e73a50ade19835fa1a0202df43c7a4e4881b|2.57|2014-09-11 10:06:00|1.4091206135396188|3||66|0.6119093465164359|0|47|523|-80.816172|64|35.059823|FRESH POTATOES|0.0|4|COO SWEET POTATOES, BULK|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00204091000004|FRESH PRODUCE|PRODUCE|-80.816172|1.4105082902580508|66|1
35.059823|663f8f3dbc3a6aaf928a56ebdbb9bf8cc90c3e72|4.49|2015-02-16 20:42:00|80.816179662140996|3|70897191697|66|35.080284602722699|0|41|1703|-80.8955|387|35.4437|SEASONAL COOKIES|1.5|14|RED VELVET FRSTD SUGAR COOKIES|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|35.070508771677183|00708971916978|COOKIES|BAKERY|-80.816172|80.816262761970094|272|1
35.059823|013988bc2d1d4d4fd58c71416c16d6a053f6923d|4.18|2014-11-11 17:50:00|1.4091206135396188|3|20165700000|66|0.6119093465164359|0|47|297|-80.816172|49|35.059823|GROUND BEEF|0.93|2|HT GROUND BEEF CHUCK 80% LEAN|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00201657000003|BEEF|MEAT|-80.816172|1.4105082902580508|66|1
35.059823|a0b3942b9e330e27d8b20219cf8c25e5d2ee84ef|7.99|2014-11-22 22:21:00|1.4091206135396188|3|8382010401|66|0.6119093465164359|0|47|459|-80.816172|83|35.059823|IMPORT BEER|0.0|16|GUINNESS DRAUGHT 6PK|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00083820104011|IMPORT BEER|BEER|-80.816172|1.4105082902580508|66|1
35.059823|ada133bb34c7741f2acfee145a35f1e56ac12715|8.99|2014-09-28 18:45:00|1.4091206135396188|3|8382010401|66|0.6119093465164359|0|47|459|-80.816172|83|35.059823|IMPORT BEER|0.0|16|GUINNESS DRAUGHT 6PK|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00083820104011|IMPORT BEER|BEER|-80.816172|1.4105082902580508|66|1
35.059823|0d5d57d2845135707ae1f7f5cf808231d7f803f0|4.59|2014-10-31 13:56:00|1.4091206135396188|3|4480000142|66|0.6119093465164359|0|47|225|-80.816172|35|35.059823|SUGAR-GRANULATED|0.0|1|SUGAR IN THE RAW|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00044800001423|SUGAR/SUBSTITUTES|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|b70b82fb9f3e5de6eed7ff0d9adf1e278fc2b0d4|2.79|2014-09-26 09:46:00|1.4091206135396188|3|1800000501|66|0.6119093465164359|0|47|328|-80.816172|54|35.059823|SWEET ROLLS-REFRIGERATED|0.79|3|PILLSBURY CINNAMON ROLLS|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00018000005017|DOUGH PRODUCTS|DAIRY|-80.816172|1.4105082902580508|66|1
35.059823|a43c84a736be65c3a8a516ee62d8720ebd89bf71|4.29|2015-02-07 17:28:00|1.4091206135396188|3|2840006399|66|0.6119093465164359|0|47|204|-80.816172|31|35.059823|TORTILLA CHIPS|0.29|1|TOSTITOS MULTIGRAIN SCOOPS|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00028400036337|SNACKS|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|c5fc14c5d7a9a916ec04377f1f80febbc8854233|1.49|2014-11-12 19:40:00|1.4091206135396188|3|7203688005|66|0.6119093465164359|0|47|555|-80.816172|64|35.059823|PACKAGED SALADS|0.0|4|HT GARDEN SALAD 16 OZ|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00072036880055|FRESH PRODUCE|PRODUCE|-80.816172|1.4105082902580508|66|1
35.059823|50275605d3c52abfb3f650448afa5847a7123be3|0.99|2014-10-03 14:16:00|1.4091206135396188|3|3400000031|66|0.6119093465164359|0|47|47|-80.816172|7|35.059823|REGISTER BARS|0.49|1|COOKIES CREME SINGLE BAR|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00034000002399|CANDY|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|30c67c3c422f85d1910912bdec67f9b87f2500b3|8.54|2014-12-15 13:05:00|1.4091206135396188|3|20332900000|66|0.6119093465164359|0|47|641|-80.816172|137|35.059823|PREMIUM PORK|0.0|2|PORK SIRLOIN ROAST BONELESS|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00203329000007|PORK|MEAT|-80.816172|1.4105082902580508|66|1
35.059823|c83ed22e70295139b30fb411139ff0303eeaa9de|10.98|2015-02-20 21:57:00|1.4091206135396188|3|4400003442|66|0.6119093465164359|0|47|91|-80.816172|13|35.059823|SPRAYED BUTTER CRACKERS|2.98|1|RITZ FAMILY SIZE|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00044000034429|CRACKERS|G1 GROCERY|-80.816172|1.4105082902580508|66|2
35.059823|88183d8ab0e45821905af53ea04b1b20d12bea28|1.69|2015-03-02 16:37:00|1.4091206135396188|3|4900000977|66|0.6119093465164359|0|47|31|-80.816172|4|35.059823|NON CARBONATED WATER|0.0|1|CB DASANI WATER 20 OZ SINGLES|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00049000009774|BOTTLED WATER|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|ddf35708a20d4272d2bcda53c6564e4494a59995|2.99|2015-01-20 18:52:00|1.4091206135396188|3|5100015339|66|0.6119093465164359|0|47|137|-80.816172|20|35.059823|TOMATO & VEGETABLE JUICE|1.0|1|V8 VFUSION POMEGRANTE BLUEBRY|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00051000169839|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|68c0193d5ebdb32a6a58e29b98001210982dcaa9|6.38|2014-12-03 18:15:00|1.4091206135396188|3|7203655010|66|0.6119093465164359|0|47|317|-80.816172|52|35.059823|CHUNK AND BAR CHEESE|0.69|3|HT 2% SHARP CHEDDAR CHEESE|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00072036705112|CHEESE|DAIRY|-80.816172|1.4105082902580508|66|2
35.059823|e18bf6e53a36a4054231ed10d8f5194efc90601e|4.49|2014-09-23 14:11:00|1.4091206135396188|3|7203695824|66|0.6119093465164359|0|47|2005|-80.816172|495|35.059823|BH GREEN SALADS|1.5|6|CHEF SALAD W/ BH MEAT|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00072036952073|GREEN SALADS|DELI|-80.816172|1.4105082902580508|66|1
35.059823|90b09927f0d0eefb0fe8f47531c86729e480f736|6.49|2015-02-27 21:55:00|1.4091206135396188|3|4154800385|66|0.6119093465164359|0|47|252|-80.816172|45|35.059823|PREMIUM ICE CREAM|1.61|5|EDY'S GRAND CHO CP CKIE DGH|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00041548550855|ICE CREAM|FROZEN|-80.816172|1.4105082902580508|66|1
35.059823|36c86f9d5a8a382a8f89a921fc345263c5c6f74c|3.29|2014-10-26 20:40:00|80.816179662140996|3|1410008786|66|35.080284734723769|0|41|1033|-80.78468|163|35.096737|HAMBURGER|0.0|7|PEP  WHEAT HAMBURGER BUNS PP|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|35.070508771677183|00014100087861|BUNS/ROLLS|COMMERCIAL BAKERY|-80.816172|80.816185171344543|30|1
35.059823|fa3e85d1bd8e1255fa4fbb359701f0f45f7e15d3|1.49|2014-12-06 14:15:00|1.4091206135396188|3|2840002819|66|0.6119093465164359|0|47|206|-80.816172|31|35.059823|FRONT END SNACKS|0.0|1|DORITOS NACHO CHEESE|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00028400028196|SNACKS|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|5310be065f87e52165df926ed9ccd706161f27eb|1.49|2014-12-01 15:19:00|1.4091206135396188|3|2840002819|66|0.6119093465164359|0|47|206|-80.816172|31|35.059823|FRONT END SNACKS|0.0|1|DORITOS NACHO CHEESE|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00028400028196|SNACKS|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|fd6ccf2fa7c46e2a5a9b005b11462b1b73fb1367|11.59|2015-01-17 23:44:00|1.4091206135396188|3|30045044909|66|0.6119093465164359|0|47|4296|-80.816172|1205|35.059823|ACETAMINOPHEN|2.6|17|L TYLENOL EX-ST CAPLET-44909|e656420b48b9329ea9c4b29668210b14aeea91da|1.4138566523078009|0.61242566243833529|00300450449092|PAIN RELIEF|HBC|-80.816172|1.4105082902580508|66|1
35.141204|7f2c9a1e6fe74fddae8b7e8ee08ee4395b198569|4.29|2015-01-11 19:43:00|80.739023103730261|2|2840015938|171|35.168699574318879|0|16|201|-80.771677|31|35.066546|POTATO CHIPS|2.15|1|RUFFLES REDUCED FAT|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00028400033978|SNACKS|G1 GROCERY|-80.739|80.739031129843468|45|1
35.141204|a0e2380c9ab8ef4c74f985703e7e781c88514147|4.29|2014-10-20 14:23:00|80.739023103730261|2|2840015938|171|35.168699586081864|0|16|201|-80.709466|31|35.124987|POTATO CHIPS|1.79|1|RUFFLES REDUCED FAT|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00028400033978|SNACKS|G1 GROCERY|-80.739|80.739001178142971|157|1
35.141204|fde01b5951828161ddd42a5d4334bb1b6a19958b|5.29|2014-10-09 17:28:00|80.739023103730261|2|4440018400|171|35.168699574318879|0|16|293|-80.771677|48|35.066546|FROZEN SEAFOOD|1.95|5|GORTON'S GRILLED TILAPIA|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00044400186506|FROZEN MEALS|FROZEN|-80.739|80.739031129843468|45|1
35.141204|b7a25c1e780d1176910c816d71bb45b2b2569550|5.58|2015-01-10 20:25:00|80.739023103730261|2|4310045388|171|35.168699574318879|0|16|6740|-80.771677|1564|35.066546|SCHOOL PAPER-OTHER|0.0|18|FIVE STAR FAT NTBK 200CT|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00043100453888|SCHOOL & OFFICE SUPPLY|GM|-80.739|80.739031129843468|45|2
35.141204|a7e50ef80eaf23c6dcf3fa0fe512403d48f17672|1.39|2015-03-06 16:56:00|80.739023103730261|2|4144310303|171|35.168699574318879|0|16|242|-80.771677|39|35.066546|CANNED BEANS|0.0|1|M HOLMES SND PINTO BEANS|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00041443119539|VEGETABLES-CAN/JAR|G1 GROCERY|-80.739|80.739031129843468|45|1
35.141204|be214092743bdc7ecccc6c6787adba2c85dd13b0|3.6|2014-10-28 20:20:00|80.739023103730261|2|4800000245|171|35.168699546082586|0|16|190|-80.847383|29|35.024464|TUNA-CANNED|0.29|1|COS TUNA CHUNK LIGHT|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00048000002457|SEAFOOD-CANNED|G1 GROCERY|-80.739|80.739057375210805|317|4
35.141204|9339c752a779c6b794aef08843068b133100549d|1.59|2014-10-18 18:09:00|80.739023103730261|2|4650073332|171|35.168699574318879|0|16|393|-80.771677|68|35.066546|NFS-AIR FRESHENERS|0.59|1|GLADE AEROSOL PURE VANILLA|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00046500745393|FRESHENERS/DEODORIZERS|G1 GROCERY|-80.739|80.739031129843468|45|1
35.141204|5dd5699884d590fd2cde8b37f31bafd24a49d49f|3.99|2014-10-21 17:27:00|80.739023103730261|2|7203663995|171|35.168699574318879|0|16|342|-80.771677|57|35.066546|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00072036631282|MILK|DAIRY|-80.739|80.739031129843468|45|1
35.141204|a315f823b9ec4282cd3e0906c020365f525cbd60|7.98|2014-10-04 18:32:00|80.739023103730261|2|7203663995|171|35.168699566405451|0|16|342|-80.816172|57|35.059823|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00072036631282|MILK|DAIRY|-80.739|80.739040249992613|66|2
35.141204|453295349d90df715df12170acf809fb95f9799a|7.98|2014-10-11 05:10:00|80.739023103730261|2|7203663995|171|35.16869957992747|0|16|342|-80.78468|57|35.096737|FRESH MILK|1.02|3|HARRIS TEETER FF SKIM MILK|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00072036631282|MILK|DAIRY|-80.739|80.739022531701465|30|2
35.141204|912f7421bbc89fb3a197ba460bd176df8a6f0019|7.98|2014-11-08 17:27:00|80.739023103730261|2|7203663995|171|35.168699585978139|0|16|342|-80.80146|57|35.17739|FRESH MILK|1.02|3|HARRIS TEETER FF SKIM MILK|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00072036631282|MILK|DAIRY|-80.739|80.73900314985741|208|2
35.141204|d9b5adc8c4c755ca6181d6a2675a46947563c6ab|6.98|2015-01-01 08:08:00|1.4091206135396188|2|7203663995|171|0.6133297129150015|0|47|342|-80.739|57|35.141204|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|0.61242566243833529|00072036631282|MILK|DAIRY|-80.739|1.4091613847677018|171|2
35.141204|3db7c59068e3ede7cbea1c6a07afaa6f50f9934e|7.98|2014-11-01 14:50:00|80.739023103730261|2|7203663995|171|35.168699574318879|0|16|342|-80.771677|57|35.066546|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00072036631282|MILK|DAIRY|-80.739|80.739031129843468|45|2
35.141204|62b959691fdc819ebe5e9bfa0574f1cad19414f0|4.9|2014-10-16 15:01:00|80.739023103730261|2|7203663217|171|35.168699580415677|0|16|330|-80.824767|55|35.116751|EGGS|0.45|3|HT GRADE A LARGE EGGS 18 CT|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00072036632173|EGGS FRESH|DAIRY|-80.739|80.739021622112489|294|2
35.141204|1ecb1a68ce714bb1fb4ac77b8b99aa4d979d1654|7.98|2014-11-28 13:17:00|80.739023103730261|2|7203663995|171|35.168699566405451|0|16|342|-80.816172|57|35.059823|FRESH MILK|1.52|3|HARRIS TEETER FF SKIM MILK|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00072036631282|MILK|DAIRY|-80.739|80.739040249992613|66|2
35.141204|9b727c82a0dc973553e0990320269d25ad8104d5|2.03|2014-10-09 18:26:00|80.739023103730261|2||171|35.168699574318879|0|16|522|-80.771677|64|35.066546|FRESH TOMATOES|1.36|4|RED H/H TOMATOES, BULK|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00204799000009|FRESH PRODUCE|PRODUCE|-80.739|80.739031129843468|45|1
35.141204|8f6295b80c228d037d4922574643f6abdbd9e346|2.34|2015-01-27 17:25:00|80.739023103730261|2||171|35.168699585978139|0|16|522|-80.80146|64|35.17739|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00204664000004|FRESH PRODUCE|PRODUCE|-80.739|80.73900314985741|208|1
35.141204|4545df7c9482568eea120c257a4c7aa9615fcaa3|5.29|2014-10-15 20:39:00|80.739023103730261|2|38151918161|171|35.168699574318879|0|16|3530|-80.771677|1045|35.066546|SHAMPOO-MID PRICE|0.0|17|HERBAL ESS SH NAKED VOLUME|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00381519181504|HAIR & SCALP CARE|HBC|-80.739|80.739031129843468|45|1
35.141204|d2e1a83f6bd9fd6e07a63f39ead5ec58d3d4e454|2.77|2014-10-03 16:46:00|80.739023103730261|2|3338353030|171|35.168699585978139|0|16|523|-80.80146|64|35.17739|FRESH POTATOES|0.0|4|RUSSET POTATO 8LB BAG|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00033383530307|FRESH PRODUCE|PRODUCE|-80.739|80.73900314985741|208|1
35.141204|ed7cb532f2ef35168b0dd79576040bd628b82704|4.49|2014-10-19 17:36:00|80.739023103730261|2|2560000226|171|35.168699574318879|0|16|1046|-80.771677|173|35.066546|CAKES|0.0|7|TSTYKAKE PNUT BUTTR KANDYKAKE|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00025600002261|SWEET BAKED GOODS|COMMERCIAL BAKERY|-80.739|80.739031129843468|45|1
35.141204|b93671b6495b1ebbbfaea4662577b9902764a19e|4.19|2015-01-20 18:26:00|80.739023103730261|2|4812110208|171|35.168699574318879|0|16|1037|-80.771677|164|35.066546|ENGLISH MUFFINS|2.1|7|THOMAS ENG MUFFN ORIG 6 PK PP|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00048121102081|BREAKFAST|COMMERCIAL BAKERY|-80.739|80.739031129843468|45|1
35.141204|1af3cebedc5d0e09e20047da529b03c7c84a4044|2.79|2015-01-13 17:01:00|80.739023103730261|2|5150024136|171|35.168699580415677|0|16|125|-80.824767|19|35.116751|PEANUT BUTTER|0.0|1|JIF TO GO 8 PK|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00051500241363|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.739|80.739021622112489|294|1
35.141204|52e599a2463d93bd01bc0db48998890cc051431d|6.38|2014-09-30 19:51:00|80.739023103730261|2|3100090028|171|35.168699580415677|0|16|270|-80.824767|307|35.116751|DESSERTS FROZEN|1.38|5|BER SS TRIPLE CHOC STRATA|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00031000900281|DESSERTS FROZEN|FROZEN|-80.739|80.739021622112489|294|2
35.141204|d3028c0c4b36004b6d053eaf0bd1c98afff3b189|5.26|2014-09-30 20:09:00|80.739023103730261|2|3800039103|171|35.168699580415677|0|16|81|-80.824767|9|35.116751|RTE CEREAL KIDS|0.0|1|KELLOGG SMACKS|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00038000391033|CEREAL|G1 GROCERY|-80.739|80.739021622112489|294|2
35.141204|d20194d63c8d44e5f5a1aa304439419eb52dcf23|3.79|2015-02-01 17:07:00|80.739023103730261|2|4400002854|171|35.168699574318879|0|16|1248|-80.771677|12|35.066546|SANDWICH COOKIES|0.29|1|OREO LEMON TWIST|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00044000031015|COOKIES|G1 GROCERY|-80.739|80.739031129843468|45|1
35.141204|e8ac8adcde89081ebbc17d8109094c57934fb6b6|7.69|2015-01-07 16:52:00|80.739023103730261|2|6233885120|171|35.168699580415677|0|16|393|-80.824767|68|35.116751|NFS-AIR FRESHENERS|3.84|1|AIRWICK CHANGE CANDLE SWT PEA|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00062338883137|FRESHENERS/DEODORIZERS|G1 GROCERY|-80.739|80.739021622112489|294|1
35.141204|2ea05345fd83c128c94cd777d702219ffbaf6c12|1.19|2014-11-23 16:35:00|80.739023103730261|2|4178900701|171|35.168699586081864|0|16|1203|-80.709466|33|35.124987|RAMEN|0.19|1|YAKISOBA NDL TERIYAKI|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00041789007071|SOUP|G1 GROCERY|-80.739|80.739001178142971|157|1
35.141204|33ba1de8ca8673690f7a8b99f9ec5ceac6388281|9.98|2014-10-26 18:01:00|80.739023103730261|2|8265750406|171|35.168699580415677|0|16|31|-80.824767|4|35.116751|NON CARBONATED WATER|2.0|1|(U)DEER PARK WATER 24PK .5LT|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00082657504063|BOTTLED WATER|G1 GROCERY|-80.739|80.739021622112489|294|2
35.141204|4e825ed243164390e80d5793ae865d81abfe8447|9.05|2014-12-30 11:42:00|80.739023103730261|2||171|35.168699549657333|0|16|523|-80.737839|64|35.297134|FRESH POTATOES|1.5|4|COO SWEET POTATOES, BULK|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00204091000004|FRESH PRODUCE|PRODUCE|-80.739|80.739054752532496|258|2
35.141204|63ee5fa5d58b7c440f3e61b85909388c452350a7|2.19|2015-02-14 13:34:00|80.739023103730261|2|3760010743|171|35.168699585093449|0|16|175|-80.825175|27|35.152722|CANNED MEATS|0.69|1|HORMEL CHILI TURKEY BEANS|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00037600107433|PREPARED FOODS-RTS|G1 GROCERY|-80.739|80.739009093941007|160|1
35.141204|5fea737dc188c02370b1cb6b34b78ae412de0974|15.99|2014-11-11 17:54:00|1.4091206135396188|2|87126000465|171|0.6133297129150015|0|47|740|-80.739|87|35.141204|NFS-ROSE BQT|0.0|9|DZ ROSE BQT 3 RED/5 COLOR  ELI|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|0.61242566243833529|00871260004653|FLORAL|FLORAL|-80.739|1.4091613847677018|171|1
35.141204|5824efd94ccdaa083cd3f27e0a15b952b91e8f97|1.77|2014-10-17 16:31:00|80.739023103730261|2|7203698067|171|35.168699574318879|0|16|365|-80.771677|56|35.066546|REFRIGERATED TEAS|0.27|3|HARRIS TEETER DECAF SWEET TEA|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00072036710208|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.739|80.739031129843468|45|1
35.141204|9774232f7f3aa1308cc5e13b91bfaec6d532ae8d|21.92|2014-12-07 15:30:00|80.739023103730261|2|3700013885|171|35.168699574318879|0|16|389|-80.771677|66|35.066546|NFS-LAUNDRY DETERGENTS|1.0|1|TIDE SWEET DREAMS DOWNY 50OZ|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00037000874782|DETERGENTS|G1 GROCERY|-80.739|80.739031129843468|45|4
35.141204|81880dd1f675c2d2d11cd3b267596da885778640|2.0|2014-09-21 13:30:00|80.739023103730261|2|78352032108|171|35.168699574318879|0|16|8598|-80.771677|1792|35.066546|NEWSPAPERS|0.0|18|SUNDAY CHARLOTTE OBSERVER|e95c23cde0c7c30b7a40f3ca6f4b11d4ed00be69|1.8998785999593752|35.169056414731678|00783520321083|NEWSPAPERS|GM|-80.739|80.739031129843468|45|1
35.006282|4e353aa56ef3c26133ff5d6d9f12b4003901f824|5.38|2014-10-13 12:12:00|1.4091206135396188|3|7225001739|60|0.6109748797816256|0|47|1025|-80.562829|162|35.006282|WHITE|1.34|7|NATOWN WHITEWHEAT RTOP BRD|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00072250017398|SLICED BREAD|COMMERCIAL BAKERY|-80.562829|1.4060866207711706|60|2
35.006282|17f1ddbbaf6ba8abde6182fe9ea05aaa4f48574e|6.99|2014-09-17 12:02:00|1.4091206135396188|3||60|0.6109748797816256|0|47|1347|-80.562829|64|35.006282|PUMPKINS|1.99|4|CARVING PUMPKINS, LARGE|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00204737000009|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|1
35.006282|83ef4aedb2238e63974afb12fc4b97b06a34c7b6|2.39|2015-02-27 12:19:00|1.4091206135396188|3|4132100541|60|0.6109748797816256|0|47|184|-80.562829|28|35.006282|SALAD DRESSINGS-LIQUID|0.39|1|WISHBONE DRS VIN ITALIANHOUSE|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00041321006470|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.562829|1.4060866207711706|60|1
35.006282|95f97b87f84a1a767934464c1d30cbb7afb3ca8c|3.89|2014-09-27 15:18:00|1.4091206135396188|3|4400003219|60|0.6109748797816256|0|47|1249|-80.562829|12|35.006282|CHOCOLATE CHIP COOKIES|0.89|1|CHIPS AHOY CHEWY|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00044000032234|COOKIES|G1 GROCERY|-80.562829|1.4060866207711706|60|1
35.006282|9248b8fa2a991b6877c535db888abacde3eff392|3.89|2015-01-17 13:44:00|80.562862110758871|3|4400003219|60|35.053759739563525|0|21|1249|-80.64817|12|35.04711|CHOCOLATE CHIP COOKIES|0.89|1|CHIPS AHOY CHEWY|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|35.054042368968126|00044000032234|COOKIES|G1 GROCERY|-80.562829|80.56283126572356|129|1
35.006282|6ac889c651d643b2438e362b394405d5e6e31154|3.99|2015-02-11 15:25:00|80.562862110758871|3|4400003219|60|35.053759739563525|0|21|1249|-80.64817|12|35.04711|CHOCOLATE CHIP COOKIES|0.99|1|CHIPS AHOY CHEWY|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|35.054042368968126|00044000032234|COOKIES|G1 GROCERY|-80.562829|80.56283126572356|129|1
35.006282|4eff0d4d56e7015c8b166746574f78ae716ce32d|1.79|2014-10-17 11:03:00|1.4091206135396188|3|7339000393|60|0.6109748797816256|0|47|48|-80.562829|7|35.006282|REGISTER GUM|0.4|1|MENTOS RED FRUIT GUM 15CT|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00073390003937|CANDY|G1 GROCERY|-80.562829|1.4060866207711706|60|1
35.006282|1c52ea8647387aaf95b8f9ae6fe7278c9ce9d922|2.0|2014-11-13 11:22:00|1.4091206135396188|3|4300000953|60|0.6109748797816256|0|47|272|-80.562829|307|35.006282|TOPPINGS FROZEN|1.01|5|COOL WHIP WHIPPED TOPPING|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00043000009536|DESSERTS FROZEN|FROZEN|-80.562829|1.4060866207711706|60|1
35.006282|d8158057241afc0f1bd477341513447bd558c64f|7.99|2015-02-12 10:36:00|80.562862110758871|3|4145810534|60|35.053759739563525|0|21|265|-80.64817|307|35.04711|FROZEN PIES|0.0|5|EDWARDS CHOC CREAM W/HERSHEY'S|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|35.054042368968126|00041458105565|DESSERTS FROZEN|FROZEN|-80.562829|80.56283126572356|129|1
35.006282|dec22e250b3ffe777625643f892c5355e0279f9d|1.99|2015-03-05 13:54:00|1.4091206135396188|3|7203688083|60|0.6109748797816256|0|47|526|-80.562829|64|35.006282|FRESH MUSHROOMS|0.0|4|HT WHITE MUSHROOMS, 8 OZ WHOLE|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00072036880833|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|1
35.006282|f62c836b7207185a7e5d3b17c39e12d5a1f1e57a|1.69|2015-01-23 09:56:00|1.4091206135396188|3|7203688003|60|0.6109748797816256|0|47|527|-80.562829|64|35.006282|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00072036880031|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|1
35.006282|75d4f67ee67545447b4bedd75b411d8e9e5c12d7|1.79|2015-02-05 11:22:00|1.4091206135396188|3|7203688032|60|0.6109748797816256|0|47|555|-80.562829|64|35.006282|PACKAGED SALADS|0.0|4|HT SHREDDED ICEBERG LETTUCE|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00072036880321|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|1
35.006282|51abd474ac0573e6436f684a063a10fad23a343e|1.79|2014-09-10 10:44:00|1.4091206135396188|3|7203688032|60|0.6109748797816256|0|47|555|-80.562829|64|35.006282|PACKAGED SALADS|0.0|4|HT SHREDDED ICEBERG LETTUCE|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00072036880321|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|1
35.006282|3bf74bf87ad41ab98433393a8aab99e96f868cde|1.79|2015-01-31 12:33:00|1.4091206135396188|3|7203688032|60|0.6109748797816256|0|47|555|-80.562829|64|35.006282|PACKAGED SALADS|0.29|4|HT SHREDDED ICEBERG LETTUCE|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00072036880321|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|1
35.006282|fc5389be7ee18c23b6c74443b58b06e450afa938|1.79|2014-10-11 11:09:00|1.4091206135396188|3|7203688032|60|0.6109748797816256|0|47|555|-80.562829|64|35.006282|PACKAGED SALADS|0.0|4|HT SHREDDED ICEBERG LETTUCE|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00072036880321|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|1
35.006282|8741b9c29d4780fdf0c4533b32e34099ea0d482b|9.99|2015-02-20 12:26:00|1.4091206135396188|3|7274506839|60|0.6109748797816256|0|47|640|-80.562829|201|35.006282|MARINATED POULTRY|0.0|2|PERDUE PERFECT BNLS BREAST|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00072745068393|POULTRY|MEAT|-80.562829|1.4060866207711706|60|1
35.006282|7d4d98e0d03e768646fe7c993a398f902cab2587|2.79|2014-12-09 11:33:00|1.4091206135396188|3|7878390810|60|0.6109748797816256|0|47|561|-80.562829|64|35.006282|FR PROD ORGANIC PRODUCE|0.79|4|ORG CARROTS, PETITE 12OZ BAG|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00078783908103|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|1
35.006282|776740118530a8e6a03f43fc83115968e6400ffc|1.54|2014-10-19 13:02:00|1.4091206135396188|3||60|0.6109748797816256|0|47|523|-80.562829|64|35.006282|FRESH POTATOES|0.36|4|COO SWEET POTATOES, BULK|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00204091000004|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|1
35.006282|e0914758d54a0d81e3683f2420dcfa3633c50dae|1.27|2015-01-29 12:13:00|1.4091206135396188|3||60|0.6109748797816256|0|47|523|-80.562829|64|35.006282|FRESH POTATOES|0.0|4|COO SWEET POTATOES, BULK|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00204091000004|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|1
35.006282|2b3d52b45cb95fd93dbde33e57407a99faeff33c|1.25|2014-11-09 12:51:00|1.4091206135396188|3||60|0.6109748797816256|0|47|523|-80.562829|64|35.006282|FRESH POTATOES|0.39|4|COO SWEET POTATOES, BULK|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00204091000004|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|1
35.006282|f23e2c422f5e938d491e61b1de11281a7fc7c61f|1.46|2015-01-10 11:16:00|1.4091206135396188|3||60|0.6109748797816256|0|47|523|-80.562829|64|35.006282|FRESH POTATOES|0.0|4|COO SWEET POTATOES, BULK|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00204091000004|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|1
35.006282|f3edd92e50ec0b76e4659a5c116f805df179dcf2|1.68|2014-11-22 10:31:00|1.4091206135396188|3||60|0.6109748797816256|0|47|523|-80.562829|64|35.006282|FRESH POTATOES|1.03|4|COO SWEET POTATOES, BULK|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00204091000004|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|1
35.006282|4521243203e9eacaaf2f6fa193ad1d5904ea0ff5|1.75|2014-09-29 11:27:00|1.4091206135396188|3||60|0.6109748797816256|0|47|523|-80.562829|64|35.006282|FRESH POTATOES|0.4|4|COO SWEET POTATOES, BULK|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00204091000004|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|1
35.006282|fc142be952bcbe41c1e3e029cd8bacc9e3112842|5.38|2014-09-19 11:36:00|1.4091206135396188|3|20337400000|60|0.6109748797816256|0|47|641|-80.562829|137|35.006282|PREMIUM PORK|2.45|2|PORK LOIN CNTER CUT CHOPS BNLS|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00203374000007|PORK|MEAT|-80.562829|1.4060866207711706|60|1
35.006282|eb3c6179f757addd1ad020f35b20e0b1d05ba980|1.67|2014-12-22 09:56:00|1.4091206135396188|3|3120001605|60|0.6109748797816256|0|47|106|-80.562829|16|35.006282|CRANBERRY SAUCE|0.17|1|OS CRANBERRY SC JELLIED|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00031200016058|FRUIT-CAN/JAR|G1 GROCERY|-80.562829|1.4060866207711706|60|1
35.006282|b688ef62567c46b8d8c21c1eca8084a152eea059|3.75|2015-01-03 11:02:00|1.4091206135396188|3|4610000012|60|0.6109748797816256|0|47|318|-80.562829|52|35.006282|SHREDDED/GRATED CHEESE|1.25|3|SARGENTO OTB SHRP CHEDD FINE C|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00046100000663|CHEESE|DAIRY|-80.562829|1.4060866207711706|60|1
35.006282|45b0daacf3ea37074c73f0d06ded48915cee9e90|36.81|2014-11-23 14:33:00|1.4091206135396188|3|20001200000|60|0.6109748797816256|0|47|974|-80.562829|201|35.006282|FRESH TURKEY|10.78|2|BUTTERBALL FRSH HEN TRKY 10-15|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00200012000009|POULTRY|MEAT|-80.562829|1.4060866207711706|60|1
35.006282|3f0e8e30bd3c1604d6c9388d626e662eff447d06|3.35|2014-12-21 10:46:00|80.562862110758871|3|2840005597|60|35.053759739563525|0|21|199|-80.64817|31|35.04711|DIPS & SALSAS|0.35|1|TOSTITOS MILD SALSA|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|35.054042368968126|00028400055970|SNACKS|G1 GROCERY|-80.562829|80.56283126572356|129|1
35.006282|fbbd2a534aefc8e9e1b1c098ffb75462fa68a1c9|1.39|2014-09-28 13:19:00|1.4091206135396188|3|1254661959|60|0.6109748797816256|0|47|48|-80.562829|7|35.006282|REGISTER GUM|0.0|1|TRIDENT TROPICAL TWIST|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00012546619592|CANDY|G1 GROCERY|-80.562829|1.4060866207711706|60|1
35.006282|6c6e6f4ab4bd58566f77a7f99d12b73c5d4a63e4|1.17|2014-10-09 11:50:00|1.4091206135396188|3||60|0.6109748797816256|0|47|523|-80.562829|64|35.006282|FRESH POTATOES|0.0|4|"COO RED POTATO ""A""SIZE, BULK"|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00204073000008|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|1
35.006282|3a6aea77e508bd6ca6a0a7934bbf61dc1d1e5827|1.98|2015-01-30 12:04:00|1.4091206135396188|3||60|0.6109748797816256|0|47|509|-80.562829|64|35.006282|FRESH CITRUS-REMAINING|0.0|4|MINNEOLA TANGELOS|e9f3320ce36c5807a17916fec016e539cc63cf14|3.2805971517077825|0.61242566243833529|00204383000002|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|2
35.096737|495cb84d6d26b86b9603f4a1bd294b1d3c91977b|7.88|2014-12-23 18:02:00|80.782094729586973|2|8265750406|30|35.106046699039943|0|27|31|-80.824767|4|35.116751|NON CARBONATED WATER|0.0|1|(U)DEER PARK WATER 24PK .5LT|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00082657504063|BOTTLED WATER|G1 GROCERY|-80.78468|80.784680307739833|294|4
35.096737|ee47ee62348c0b0fbe2c21a7f7c2c5659f38bc57|10.93|2014-09-25 18:47:00|80.782094729586973|2|8265750406|30|35.106046699043247|0|27|31|-80.806073|4|35.106477|NON CARBONATED WATER|0.0|1|(U)DEER PARK WATER 24PK .5LT|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00082657504063|BOTTLED WATER|G1 GROCERY|-80.78468|80.784680052819638|4|3
35.096737|1968dcb74227be6972ff624ab92480f3a3fb0206|9.98|2014-10-26 20:14:00|80.782094729586973|2|8265750406|30|35.106046699039943|0|27|31|-80.824767|4|35.116751|NON CARBONATED WATER|2.0|1|(U)DEER PARK WATER 24PK .5LT|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00082657504063|BOTTLED WATER|G1 GROCERY|-80.78468|80.784680307739833|294|2
35.096737|170ef2b842e38a93f29cc30bff8862b1904ed6a4|0.99|2014-11-12 14:53:00|80.782094729586973|2|7203695306|30|35.106046699039943|0|27|1895|-80.824767|450|35.116751|TEA|0.13|6|FFM LEMONADE|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00072036953070|BEVERAGES|DELI|-80.78468|80.784680307739833|294|1
35.096737|bfda5d8f8dd7648a17531c51d9a188414b2d9f00|2.99|2015-01-13 21:07:00|80.782094729586973|2|7535511210|30|35.106046699039943|0|27|139|-80.824767|20|35.116751|REMAINING SHELF STABLE JUICES|1.5|1|OLD ORCHARD APPLE CRNBRY 100%|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00075355112104|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.78468|80.784680307739833|294|1
35.096737|2feedb6264f079b0edaba6efcae3bcd28c9e12de|4.699999999999998|2014-12-28 14:30:00|80.782094729586973|2|7248600220|30|35.106046699039943|0|27|11|-80.824767|2|35.116751|MUFFIN MIXES|0.47|1|JIFFY CORN MUFFIN MIX|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00072486002205|BAKING MIXES|G1 GROCERY|-80.78468|80.784680307739833|294|10
35.096737|d02f067974449b152654da2c4e781978661c880a|11.58|2015-01-09 21:53:00|80.782094729586973|2|7247000603|30|35.106046699039943|0|27|1641|-80.824767|377|35.116751|PACKAGED DONUTS|0.0|14|K K 12 CT GLAZED DONUTS PP|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00072470006035|DONUTS|BAKERY|-80.78468|80.784680307739833|294|2
35.096737|ef585d69a449eb30cf7a9d9a9f8da7948aaf4f7d|1.88|2014-11-04 11:32:00|80.782094729586973|2|4133500053|30|35.106046699039943|0|27|184|-80.824767|28|35.116751|SALAD DRESSINGS-LIQUID|0.0|1|KENS DRS HONEY MUSTARD|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00041335000341|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.78468|80.784680307739833|294|1
35.096737|a37782abbc9123e9e97eaceac13538b8ca638df9|3.88|2014-10-11 12:46:00|80.782094729586973|2|4175701101|30|35.106046699039943|0|27|2020|-80.824767|505|35.116751|CHEESE SPECIALTIES|0.0|6|LAUGHING COW LITE SWISS WEDGES|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00041757011062|SPECIALTY CHEESE|DELI|-80.78468|80.784680307739833|294|4
35.096737|20b59e28c647e53799f450428a08f4f8b5b44d9f|11.67|2014-11-23 18:17:00|80.782094729586973|2|3666906138|30|35.106046699039943|0|27|499|-80.824767|110|35.116751|MEATBALLS|4.26|19|COOKED PERFECT HOMESTYLE MTBLS|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00036669061380|FROZEN CASE MEAT|CASE READY MEATS|-80.78468|80.784680307739833|294|3
35.096737|45540d94c35e52f2279f2f8449a45b06d214068c|4.0|2014-12-14 16:33:00|80.782094729586973|2|4000000435|30|35.106046699039943|0|27|47|-80.824767|7|35.116751|REGISTER BARS|0.2|1|(FE)M&M PEANUT CANDY|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00040000000327|CANDY|G1 GROCERY|-80.78468|80.784680307739833|294|4
35.096737|ef6e8ee2c406fde08a9d46828a61d89449be790a|3.25|2015-01-11 12:13:00|80.782094729586973|2|3700007100|30|35.106046699039943|0|27|393|-80.824767|68|35.116751|NFS-AIR FRESHENERS|0.25|1|I/O FEBREZE AE SPICED PEAR|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00037000898689|FRESHENERS/DEODORIZERS|G1 GROCERY|-80.78468|80.784680307739833|294|1
35.096737|ac299bd41cc661e3e2eb5632d251dcf71f084ddc|19.86|2014-12-14 17:10:00|80.782094729586973|2|4720015264|30|35.106046699039943|0|27|312|-80.824767|51|35.116751|BUTTER|0.0|3|CHALLENGE SALTED BUTTER|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00047200152641|BUTTER & MARGARINE|DAIRY|-80.78468|80.784680307739833|294|6
35.096737|41b0c98dedab4743a8b42a604b3711cb4a2f2c7f|11.97|2014-09-28 20:06:00|80.782094729586973|2|4400002854|30|35.106046699039943|0|27|1248|-80.824767|12|35.116751|SANDWICH COOKIES|4.47|1|OREO GOLDEN DOUBLE STUF|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00044000025403|COOKIES|G1 GROCERY|-80.78468|80.784680307739833|294|3
35.096737|ff72aa3285cede43237c5b859268eb384fb27e24|1.1|2015-02-16 09:27:00|80.782094729586973|2|5000000124|30|35.106046699043247|0|27|154|-80.806073|24|35.106477|NFS-CAT FOOD WET|0.0|1|FANCY FEAST SEAFOOD FEAST|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00050000429349|PET FOOD/SUPPLIES|G1 GROCERY|-80.78468|80.784680052819638|4|2
35.096737|6d4030ac0f6bea10fb617a7632b0c6cd87ae35df|6.7|2014-10-28 07:57:00|80.782094729586973|2|7203656080|30|35.106046699039943|0|27|318|-80.824767|52|35.116751|SHREDDED/GRATED CHEESE|1.8499999999999999|3|HT SHRED WISC XTRA SHARP CHED|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00072036705181|CHEESE|DAIRY|-80.78468|80.784680307739833|294|2
35.096737|b5e5b9a39acedb54f7b0ee7e9e268413feb45afc|1.29|2014-12-02 12:18:00|80.782094729586973|2|8379152001|30|35.106046699039943|0|27|1981|-80.824767|480|35.116751|CHIPS|0.0|6|DIRTY POTATO CHIP BBQ|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00083791520049|DRY GOODS|DELI|-80.78468|80.784680307739833|294|1
35.096737|07822afaecac14f8af194007ccc804854bb85ece|7.3|2014-12-13 20:03:00|80.782094729586973|2|7585600110|30|35.106046699039943|0|27|273|-80.824767|43|35.116751|PREMIUM NOVELTIES|0.0|5|KLONDIKE HEATH BAR|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00075856011135|FROZEN NOVELTIES|FROZEN|-80.78468|80.784680307739833|294|2
35.096737|678665515692e5f4b76cf285ddb78fe3e01bb219|5.49|2014-09-13 20:19:00|80.782094729586973|2|4450098196|30|35.106046699039943|0|27|839|-80.824767|102|35.116751|STACK PACKS|0.0|19|HF CLASSIC SMOKED HAM|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00044500981995|LUNCHMEATS|CASE READY MEATS|-80.78468|80.784680307739833|294|1
35.096737|a63f2c92f21beadadba1f7fbb2615f2cd8b7e8cd|2.72|2015-01-21 17:32:00|80.782094729586973|2||30|35.106046699039943|0|27|500|-80.824767|64|35.116751|FRESH APPLES|0.0|4|HONEY CRISP APPLE|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00233283000003|FRESH PRODUCE|PRODUCE|-80.78468|80.784680307739833|294|1
35.096737|c7f7feb4fc19d46db93298ff9a36d13c98b8eec8|2.59|2015-02-12 15:21:00|80.782094729586973|2|7203695296|30|35.106046696329372|0|27|1654|-80.80146|381|35.17739|DESSERT CAKES|0.0|14|RED VELVET CAKE SLICE|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00072036952967|CAKES|BAKERY|-80.78468|80.784688688800259|208|1
35.096737|fb6f329d65161839be437f68d088c70c9e97dc4f|3.94|2014-12-07 21:19:00|80.782094729586973|2|73621195143|30|35.106046699039943|0|27|1687|-80.824767|385|35.116751|THAW & SELL (SWEET GOODS)|0.0|14|MINI CINNAMON ROLLS|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00736211951434|SWEET GOODS|BAKERY|-80.78468|80.784680307739833|294|2
35.096737|237956d46a1e56572cb596d1069b2e1f5787c7e7|5.99|2014-11-16 20:36:00|80.782094729586973|2|73621195143|30|35.106046699039943|0|27|1687|-80.824767|385|35.116751|THAW & SELL (SWEET GOODS)|4.52|14|MINI CINNAMON ROLLS|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00736211951434|SWEET GOODS|BAKERY|-80.78468|80.784680307739833|294|1
35.096737|f97ba20ace62318ed9a28e16d74e5c8a87c221ec|6.49|2014-10-18 17:39:00|80.782094729586973|2|7478091136|30|35.106046699039943|0|27|30|-80.824767|4|35.116751|CARBONATED WATER|0.8|1|PERRIER .5L 6PK PET|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00074780911368|BOTTLED WATER|G1 GROCERY|-80.78468|80.784680307739833|294|1
35.096737|7a1988049444337b77162805204c3ac89ef7edb3|2.99|2015-02-16 22:07:00|80.782094729586973|2|7294560136|30|35.106046696329372|0|27|1026|-80.80146|162|35.17739|WHEAT|0.5|7|S L HONEY WHEAT BREAD|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00072945601369|SLICED BREAD|COMMERCIAL BAKERY|-80.78468|80.784688688800259|208|1
35.096737|bad1d7c5cd163a8827dbd9b5133a67ea49f5e1fb|20.97|2014-11-21 20:48:00|80.782094729586973|2|3913116852|30|35.106046699039943|0|27|254|-80.824767|892|35.116751|PREMIUM PIZZA|5.97|5|BELLATORIA ULTIMATE PEPPERONI|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00039131168525|FROZEN PIZZA|FROZEN|-80.78468|80.784680307739833|294|3
35.096737|6e6932a46c8aaf74e2b986937a51b97103ad29b1|1.6|2014-10-12 22:05:00|80.782094729586973|2|7047000641|30|35.106046699039943|0|27|687|-80.824767|61|35.116751|BLENDED|0.3|3|YOPLAIT T/C KEY LIME PIE|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00070470180823|YOGURT|DAIRY|-80.78468|80.784680307739833|294|2
35.096737|d43ec019781c87ae90c1805110c135b7d9b46076|3.47|2014-12-21 11:41:00|80.782094729586973|2||30|35.106046699039943|0|27|566|-80.824767|64|35.116751|SERVICE BAR|0.24|4|HT 7 LAYER MEXICAN BEAN DIP|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00204506000001|FRESH PRODUCE|PRODUCE|-80.78468|80.784680307739833|294|1
35.096737|8042f292e02d4816436bf0eeb245a5af7f9805c5|9.99|2015-02-08 20:54:00|80.782094729586973|2|30997390801|30|35.106046696329372|0|27|3045|-80.80146|1000|35.17739|BRAND-REVLON|0.0|17|PHOTOREADY 3D VOL MASC BLK/BLK|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00309973908017|COSMETICS|HBC|-80.78468|80.784688688800259|208|1
35.096737|50b1e8f165905360185137e3f1edc0831288ae60|4.0|2014-09-14 18:49:00|1.4091206135396188|2||30|0.612553617356517|0|47|511|-80.78468|64|35.096737|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|0.61242566243833529|00204770000004|FRESH PRODUCE|PRODUCE|-80.78468|1.4099586511700126|30|2
35.096737|9b0b727e9f10f6214e1365935b5ed219529bd88e|4.39|2015-02-03 13:31:00|80.782094729586973|2|4400002796|30|35.106046696329372|0|27|90|-80.80146|13|35.17739|SNACK CRACKERS|2.2|1|RICE THINS  BR SWEET BARBEQUE|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00044000037901|CRACKERS|G1 GROCERY|-80.78468|80.784688688800259|208|1
35.096737|0fe810936393af3b529fcf86878850a02a56c6ec|1.3|2014-10-02 22:11:00|80.782094729586973|2|5000042264|30|35.106046696954287|0|27|154|-80.739|24|35.141204|NFS-CAT FOOD WET|0.2|1|FRISKIES MARINERS CATCH|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00050000425044|PET FOOD/SUPPLIES|G1 GROCERY|-80.78468|80.784687623114351|171|2
35.096737|8b129deaa788deca51cad1e3e16e6b130171e2f8|5.58|2014-10-25 16:23:00|80.782094729586973|2|61611227958|30|35.106046699039943|0|27|581|-80.824767|136|35.116751|FRESH SALSA|0.58|4|WHOLLY GUACAMOLE CLASSIC 8OZ|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00616112279588|OTHER MERCHANDISE|PRODUCE|-80.78468|80.784680307739833|294|2
35.096737|42f1981da563827cf54a3336884f530a63d19d6b|1.35|2015-02-13 21:14:00|80.782094729586973|2||30|35.106046699043247|0|27|500|-80.806073|64|35.106477|FRESH APPLES|0.13|4|GALA APPLES|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00204135000007|FRESH PRODUCE|PRODUCE|-80.78468|80.784680052819638|4|1
35.096737|6325bda0fe897678f96b8ba0a2b934fc74a1640f|1.69|2015-03-04 08:39:00|80.782094729586973|2||30|35.106046699039943|0|27|500|-80.824767|64|35.116751|FRESH APPLES|0.85|4|FUJI APPLES|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00204131000001|FRESH PRODUCE|PRODUCE|-80.78468|80.784680307739833|294|1
35.096737|4fc484952e0d3c819c05660c62acb325c7c9987e|2.98|2014-09-21 15:05:00|80.782094729586973|2|5000000457|30|35.106046699039943|0|27|168|-80.824767|24|35.116751|NFS-CAT TREATS|0.48|1|FF APPETIZER SEA BASS & SHRIMP|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00050000004560|PET FOOD/SUPPLIES|G1 GROCERY|-80.78468|80.784680307739833|294|2
35.096737|f70da15e4ad7ae11e5252ae921c26773b367990e|2.69|2014-10-27 11:24:00|80.782094729586973|2|7203630050|30|35.106046699039943|0|27|184|-80.824767|28|35.116751|SALAD DRESSINGS-LIQUID|0.13|1|HT DRS HONEY DIJON|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00072036300553|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.78468|80.784680307739833|294|1
35.096737|ffc0400e7bc48703b9144c3085905e96ec0da328|2.69|2014-10-30 15:37:00|80.782094729586973|2|7203630050|30|35.106046699039943|0|27|184|-80.824767|28|35.116751|SALAD DRESSINGS-LIQUID|0.19|1|HT DRS HONEY DIJON|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00072036300553|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.78468|80.784680307739833|294|1
35.096737|a8a95c1674fc1e51a9fc41cbc4330cd5480b63f3|2.69|2014-12-29 14:19:00|80.782094729586973|2|7203630050|30|35.106046699039943|0|27|184|-80.824767|28|35.116751|SALAD DRESSINGS-LIQUID|0.17|1|HT DRS HONEY DIJON|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00072036300553|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.78468|80.784680307739833|294|1
35.096737|8ec475124b67857df6ce4f1f04fbf3fef5452bb7|2.49|2015-02-13 17:22:00|80.782094729586973|2|7203630050|30|35.106046696329372|0|27|184|-80.80146|28|35.17739|SALAD DRESSINGS-LIQUID|0.12|1|HT DRS HONEY DIJON|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00072036300553|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.78468|80.784688688800259|208|1
35.096737|a6f38604b2a533e1547b55a73765c9190bce2c44|3.49|2015-02-08 20:52:00|80.782094729586973|2|7203663995|30|35.106046696329372|0|27|342|-80.80146|57|35.17739|FRESH MILK|0.18|3|HARRIS TEETER 2% MILK|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00072036639981|MILK|DAIRY|-80.78468|80.784688688800259|208|1
35.096737|7f139c76928451a115d2ec3f5790be6881dcea11|6.99|2014-09-19 12:25:00|80.782094729586973|2|2301290168|30|35.106046699039943|0|27|1477|-80.824767|485|35.116751|SUSHI HYBRID|0.0|6|CRUNCHY CA ROLL SP BR RICE|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00023012901684|SUSHI|DELI|-80.78468|80.784680307739833|294|1
35.096737|961ac66d8249401fffb778c4cf8c259e614783ed|3.3|2015-01-25 16:23:00|80.782094729586973|2|5000000124|30|35.106046699039943|0|27|154|-80.824767|24|35.116751|NFS-CAT FOOD WET|0.0|1|FANCY FEAST FLAKED FISH&SHRIMP|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00050000428748|PET FOOD/SUPPLIES|G1 GROCERY|-80.78468|80.784680307739833|294|6
35.096737|8fb22d8867f802b5c59ed2c9e20727f3caf7b942|1.89|2015-01-30 19:05:00|80.782094729586973|2|3400000220|30|35.106046696329372|0|27|47|-80.80146|7|35.17739|REGISTER BARS|0.0|1|HERSHY MLK CHOC W/ALMDS KING|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00034000002214|CANDY|G1 GROCERY|-80.78468|80.784688688800259|208|1
35.096737|172c15a13073b8c38fe823c7fff68b61486d16b3|1.0|2014-12-02 11:27:00|80.782094729586973|2|3400000031|30|35.106046699039943|0|27|47|-80.824767|7|35.116751|REGISTER BARS|0.25|1|HERSHEY ALMOND BAR|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00034000002412|CANDY|G1 GROCERY|-80.78468|80.784680307739833|294|1
35.096737|bcffff0b0cbd747e32cedc7a9f70cf670144559a|0.77|2014-10-31 09:11:00|80.782094729586973|2|7203636010|30|35.106046699039943|0|27|30|-80.824767|4|35.116751|CARBONATED WATER|0.07|1|HT SIMPLY CLEAR TANGERINE LIME|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00072036030818|BOTTLED WATER|G1 GROCERY|-80.78468|80.784680307739833|294|1
35.096737|2a4485eefc13fa5a92224bbc3b56f68d6dc11fc4|5.99|2015-02-14 23:37:00|80.782094729586973|2|7203689258|30|35.106046696329372|0|27|563|-80.80146|64|35.17739|FRESH VEGETABLE/FRUIT TRAYS|0.0|4|CHOC STRAWBERRIES 6CT|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00072036892584|FRESH PRODUCE|PRODUCE|-80.78468|80.784688688800259|208|1
35.096737|5a12f62065a93c93e3b0f4351048f285ad94f96b|24.99|2014-09-11 19:53:00|80.782094729586973|2|70052211254|30|35.106046692741202|0|27|7185|-80.810056|1600|35.219587|SOFTSIDE COOLERS|0.0|18|RETRO LNCH BAG GRN PAISLEY|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00700522112549|SEASONAL MERCHANDISE|GM|-80.78468|80.784693240419131|401|2
35.096737|dbbd243cc4680fb25f96c8e32b57a6cb569a4d9c|17.97|2014-11-13 20:09:00|80.782094729586973|2|2840026368|30|35.106046699043247|0|27|205|-80.806073|31|35.106477|REMAINING SNACKS|3.0|1|CHEETOS HALLOWEEN 26 CTN|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00028400263689|SNACKS|G1 GROCERY|-80.78468|80.784680052819638|4|3
35.096737|1ec35bc6fa903bb96be1bd5d018448b910faf6a3|22.99|2014-09-18 14:20:00|80.782094729586973|2|7650137526|30|35.106046699039943|0|27|7182|-80.824767|1600|35.116751|HARDSIDE COOLERS|17.24|18|CLMN 20 CAN PARTY STACKER BLUE|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00076501375268|SEASONAL MERCHANDISE|GM|-80.78468|80.784680307739833|294|1
35.096737|b22360e795acb4ddf9f8b7dbdf51a0d94b3a045f|6.79|2014-10-24 12:48:00|80.782094729586973|2|7800001180|30|35.106046699039943|0|27|55|-80.824767|8|35.116751|REGULAR|3.4|23|CD GINGER ALE 12 PACK|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00078000152166|CARBONATED BEVERAGES|BEVERAGE|-80.78468|80.784680307739833|294|1
35.096737|1e857a5169a6736e81b22c0772dc3c189c8623a0|5.0|2015-02-19 18:07:00|80.782094729586973|2|3890004215|30|35.106046696329372|0|27|115|-80.80146|16|35.17739|REMAINING FRUIT|0.0|1|DOLE MANDARIN ORANGES LS|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00038900042158|FRUIT-CAN/JAR|G1 GROCERY|-80.78468|80.784688688800259|208|4
35.096737|98549625fcbf5a11638a60ed324e8b10c0cca5a9|6.48|2015-02-18 18:00:00|80.782094729586973|2|3890004215|30|35.106046696329372|0|27|115|-80.80146|16|35.17739|REMAINING FRUIT|0.0|1|DOLE MANDARIN ORANGES LS|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00038900042158|FRUIT-CAN/JAR|G1 GROCERY|-80.78468|80.784688688800259|208|4
35.096737|694e37217e7b38e70a9cca67796dc89b86817fd4|6.98|2014-11-06 21:02:00|80.782094729586973|2|2068500089|30|35.106046699043247|0|27|197|-80.806073|31|35.106477|POPPED POPCORN|0.99|1|CAPE COD WHITE CHEDDAR POPCRN|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00020685000898|SNACKS|G1 GROCERY|-80.78468|80.784680052819638|4|2
35.096737|3c06aabdcff44fb843f6e3c68a65fa0f8273d6d1|6.98|2015-02-06 22:01:00|80.782094729586973|2|2068500089|30|35.106046699039943|0|27|197|-80.824767|31|35.116751|POPPED POPCORN|1.98|1|CAPE COD WHITE CHEDDAR POPCRN|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00020685000898|SNACKS|G1 GROCERY|-80.78468|80.784680307739833|294|2
35.096737|3669bae01b9a0c08725760ccf93e69a7f01b6d6f|3.39|2014-12-28 16:04:00|80.782094729586973|2|7203620985|30|35.106046699043247|0|27|130|-80.806073|20|35.106477|CRANBERRY JUICE/DRINKS-SHELF|0.3|1|HT CRANBERRY JUICE COCKTAIL|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00072036209856|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.78468|80.784680052819638|4|1
35.096737|f303cf70a80d7d45a65434010202267c449e6b89|12.99|2014-09-10 15:49:00|80.782094729586973|2|68711011200|30|35.106046699039943|0|27|7209|-80.824767|1600|35.116751|BACK TO SCHOOL|9.74|18|EARBUDS W/INLINE MIC|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00687110111750|SEASONAL MERCHANDISE|GM|-80.78468|80.784680307739833|294|1
35.096737|61ccab8aec279cea4191ce5c013422d146a89445|3.79|2015-01-07 16:33:00|80.782094729586973|2|2100062503|30|35.106046699039943|0|27|318|-80.824767|52|35.116751|SHREDDED/GRATED CHEESE|1.29|3|KRAFT MEXICAN CHED&MONTEREY J|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00021000638970|CHEESE|DAIRY|-80.78468|80.784680307739833|294|1
35.096737|778df1732083a0370c849b9b3d50b26e5880c5b4|2.0|2014-11-28 15:43:00|80.782094729586973|2|20496400000|30|35.106046699039943|0|27|756|-80.824767|87|35.116751|NFS-FLORAL ACCESSORIES|0.0|9|*ACCESSORIES|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00204964000001|FLORAL|FLORAL|-80.78468|80.784680307739833|294|2
35.096737|23f2512eec2d5744f4a534d40e1571dfdbeb8684|1.29|2014-09-25 15:30:00|80.782094729586973|2|1657191030|30|35.106046699039943|0|27|30|-80.824767|4|35.116751|CARBONATED WATER|0.29|1|SPARKLING ICE LEMONADE|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00016571940355|BOTTLED WATER|G1 GROCERY|-80.78468|80.784680307739833|294|1
35.096737|08f40adea4dd8cfe6939d2b7aaf8c4ddaf033557|26.98|2014-12-29 11:19:00|80.782094729586973|2|84029701358|30|35.106046699039943|0|27|7329|-80.824767|1600|35.116751|CHRISTMS PRTY GOOD/DECORIMP|10.12|18|I/O WINE CHARM/STOPPER SET|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00840297013587|SEASONAL MERCHANDISE|GM|-80.78468|80.784680307739833|294|2
35.096737|9b47abc9b3cd840b00390d62cdd6e46924f8ce6d|19.18|2015-02-23 22:59:00|80.782094729586973|2|4460002031|30|35.106046696329372|0|27|730|-80.80146|24|35.17739|NFS-CAT LITTER|0.0|1|FRESH STEP CAT LITTER|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00044600020310|PET FOOD/SUPPLIES|G1 GROCERY|-80.78468|80.784688688800259|208|2
35.096737|3998fac4f69f5d871c03cb7a9fc78f1d4255d14b|3.18|2014-11-07 14:05:00|80.782094729586973|2|4280011400|30|35.106046699039943|0|27|255|-80.824767|892|35.116751|VALUE PIZZA|0.34|5|TOTINO'S PEPPERONI PIZZA|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00042800114006|FROZEN PIZZA|FROZEN|-80.78468|80.784680307739833|294|2
35.096737|657b8a3b8a69144f6b4a5434ef47058d48a2f1f9|2.5|2014-11-09 16:17:00|80.782094729586973|2|4900005537|30|35.106046699043247|0|27|55|-80.806073|8|35.106477|REGULAR|0.26|23|CLASSIC 1.25 LITER BOTTLE|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00049000055375|CARBONATED BEVERAGES|BEVERAGE|-80.78468|80.784680052819638|4|2
35.096737|3a44daa9452c677f161de5c8a3a9454fb692d775|1.25|2014-11-10 22:22:00|80.782094729586973|2|4900005537|30|35.106046699043247|0|27|55|-80.806073|8|35.106477|REGULAR|0.26|23|CLASSIC 1.25 LITER BOTTLE|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00049000055375|CARBONATED BEVERAGES|BEVERAGE|-80.78468|80.784680052819638|4|1
35.096737|e0aac5f610b96109c7d88bb542908cb8f650c2f6|11.99|2014-10-08 12:07:00|80.782094729586973|2|68332701490|30|35.106046699039943|0|27|5479|-80.824767|1502|35.116751|LARGE JAR|8.03|18|GLSS CYLINDER CNDL WH/GARDENIA|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00683327014907|CANDLES|GM|-80.78468|80.784680307739833|294|1
35.096737|1041453eb462acd64fba74d4dd906d45dfc1fce8|1.84|2014-12-17 21:15:00|80.782094729586973|2||30|35.106046699039943|0|27|503|-80.824767|64|35.116751|FRESH GRAPES|0.14|4|GREEN GRAPES, SEEDLESS 12/16|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00204022000004|FRESH PRODUCE|PRODUCE|-80.78468|80.784680307739833|294|1
35.096737|36cb85fbf5ceeb59fdf093ec09ee8002fee98dae|1.35|2015-02-26 18:04:00|80.782094729586973|2||30|35.106046699039943|0|27|565|-80.824767|64|35.116751|REDUCED PRODUCE|0.0|4|PRODUCE REWRAP BY CT|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00204845000007|FRESH PRODUCE|PRODUCE|-80.78468|80.784680307739833|294|2
35.096737|4f0514612dbc40d12052d7affa130d4b97640ea0|13.56|2015-01-21 11:31:00|80.782094729586973|2|1862770327|30|35.106046699039943|0|27|61|-80.824767|9|35.116751|RTE CEREAL ADULT|1.56|1|KASHI GO LEAN PRO FIB CEREL|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00018627703211|CEREAL|G1 GROCERY|-80.78468|80.784680307739833|294|4
35.096737|d324c67e14d6ac5b39de6e254b08544e061fe141|1.69|2014-11-20 14:28:00|80.782094729586973|2|4900000044|30|35.106046699039943|0|27|55|-80.824767|8|35.116751|REGULAR|0.0|23|CB COKE SINGLE 20 OZ.|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00049000000443|CARBONATED BEVERAGES|BEVERAGE|-80.78468|80.784680307739833|294|1
35.096737|896f89083b6cf4064007d10a3b0831dab29b0eb3|1.69|2014-10-10 11:41:00|80.782094729586973|2|4900000044|30|35.106046699039943|0|27|55|-80.824767|8|35.116751|REGULAR|0.0|23|CB COKE SINGLE 20 OZ.|ec5f5b33fe37b0956baef0110b7257cc0a0118d2|0.6432777217770961|35.102887530186244|00049000000443|CARBONATED BEVERAGES|BEVERAGE|-80.78468|80.784680307739833|294|1
35.04711|5c70caa8e1de4ea338eb5aa415b8ba531a72ddef|2.29|2015-01-29 15:28:00|1.4091206135396188|4|7203653023|129|0.6116874628086298|0|47|1273|-80.64817|50|35.04711|BAG VEG NON STEAM|0.29|5|HT GREEN PEAS|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00072036530141|VEGETABLES-FROZEN|FROZEN|-80.64817|1.407576102208115|129|1
35.04711|c5329f35eb316b85a5786ad317ad2cdc98629dfc|3.19|2014-11-20 19:03:00|1.4091206135396188|4|7203655010|129|0.6116874628086298|0|47|317|-80.64817|52|35.04711|CHUNK AND BAR CHEESE|0.0|3|HT EXTRA SHARP CHEDDAR CHEESE|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00072036559951|CHEESE|DAIRY|-80.64817|1.407576102208115|129|1
35.04711|77617f67fec25dec1f0dee3f9c324571df169439|2.89|2014-12-22 13:38:00|1.4091206135396188|4|7203663102|129|0.6116874628086298|0|47|339|-80.64817|57|35.04711|EGGNOGS/DRINKS|0.89|3|I/O HARRIS TEETER EGG NOG|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00072036631022|MILK|DAIRY|-80.64817|1.407576102208115|129|1
35.04711|8ccb948e273e415bb238150542434fe8b54db70f|4.49|2014-12-23 11:40:00|1.4091206135396188|4|3980003283|129|0.6116874628086298|0|47|8481|-80.64817|1769|35.04711|BATTERY-WATCH & CALC|0.0|18|ENERG WATCH BATTERY 2025BP|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00039800032836|BATTERY & FLASHLIGHT|GM|-80.64817|1.407576102208115|129|1
35.04711|b4214bec41c32eedba25893a5cbe8447f78a3739|8.99|2015-01-28 14:01:00|1.4091206135396188|4|4242116191|129|0.6116874628086298|0|47|1855|-80.64817|430|35.04711|BH SALAMI/CHUBBS|3.0|6|BH SUPERIORE SOPRESSATA|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00042421161915|SPECIALTY MEAT|DELI|-80.64817|1.407576102208115|129|1
35.04711|21ad8c82b26d3adf993c1a287f0640d1d22c548b|0.97|2015-01-08 17:26:00|1.4091206135396188|4|7203688002|129|0.6116874628086298|0|47|527|-80.64817|64|35.04711|FRESH CARROTS|0.0|4|HT WHOLE CARROTS 2LB BAG|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00072036880024|FRESH PRODUCE|PRODUCE|-80.64817|1.407576102208115|129|1
35.04711|9df208c6cfb604f6200654bb7e042ec448a0026a|5.35|2014-12-15 17:04:00|1.4091206135396188|4|7203697668|129|0.6116874628086298|0|47|317|-80.64817|52|35.04711|CHUNK AND BAR CHEESE|2.35|3|HT SWISS CHEESE|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00072036980465|CHEESE|DAIRY|-80.64817|1.407576102208115|129|1
35.04711|47bacbc07b4c82fceb3fbfdcfa25b174363709b3|4.99|2014-12-07 10:33:00|1.4091206135396188|4|7203695992|129|0.6116874628086298|0|47|1603|-80.64817|371|35.04711|PRIVATE LABEL BREAD|2.0|14|BAND OF BAKERS PUMPKIN BREAD|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00072036959928|BREAD|BAKERY|-80.64817|1.407576102208115|129|1
35.04711|28c1ac7c7b287848d5b030b086a64c6ac24fc1dd|1.49|2014-12-17 16:25:00|1.4091206135396188|4|2840002819|129|0.6116874628086298|0|47|206|-80.64817|31|35.04711|FRONT END SNACKS|0.0|1|LAYS CLASSIC|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00028400027960|SNACKS|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|819be91f1d11ad083f939120da0597fbe314e2f7|1.49|2015-02-13 15:15:00|1.4091206135396188|4|2840002819|129|0.6116874628086298|0|47|206|-80.64817|31|35.04711|FRONT END SNACKS|0.0|1|LAYS CLASSIC|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00028400027960|SNACKS|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|b13892e4cf05a9a6387bfe44a37ae421266a0b7e|2.29|2015-02-16 12:40:00|1.4091206135396188|4|7203663996|129|0.6116874628086298|0|47|342|-80.64817|57|35.04711|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00072036631299|MILK|DAIRY|-80.64817|1.407576102208115|129|1
35.04711|b17cc141634121497ae90cef963b014107e0b75d|2.58|2015-01-06 16:26:00|1.4091206135396188|4||129|0.6116874628086298|0|47|508|-80.64817|64|35.04711|FRESH GRAPEFRUIT|0.29|4|RED GRAPEFRUIT, FL  LRG|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00204281000005|FRESH PRODUCE|PRODUCE|-80.64817|1.407576102208115|129|2
35.04711|2c10f4d3b1871283e2cc2926687dfc6a8c5fc4f8|9.99|2014-12-20 07:52:00|1.4091206135396188|4|8858600112|129|0.6116874628086298|0|47|9949|-80.64817|886|35.04711|NFS-PREM-MERLOT|0.0|13|RED DIAMOND MERLOT|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00088586001123|PREMIUM ($8-$10.99)|WINE|-80.64817|1.407576102208115|129|1
35.04711|df51b8cadbc98c9f2280228cd2638bfdb86a4749|2.4|2014-11-29 16:45:00|1.4091206135396188|4|2400001738|129|0.6116874628086298|0|47|257|-80.64817|39|35.04711|TOMATOES|0.0|1|DEL MONTE TOMATO CHILI STYLE|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00024000012672|VEGETABLES-CAN/JAR|G1 GROCERY|-80.64817|1.407576102208115|129|2
35.04711|ae6545f0aa96ef0ad779d79197070a95fd89992e|1.47|2015-02-10 17:07:00|80.648225123995502|4|7203625014|129|35.061235468006103|0|30|145|-80.699686|22|35.000049|MILK-CANNED|0.0|1|HT SWEETENED CONDENSED MILK|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|35.078006462436761|00072036250148|PACKAGED MILKS & MODIFIERS|G1 GROCERY|-80.64817|80.648182495760508|249|1
35.04711|9ea3adabaad53d5b0c5f60de700a4832c9e0aae5|2.0|2014-12-29 17:07:00|1.4091206135396188|4||129|0.6116874628086298|0|47|511|-80.64817|64|35.04711|FRESH AVOCADOS|0.75|4|AVOCADOS, HASS XL 36CT|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00204770000004|FRESH PRODUCE|PRODUCE|-80.64817|1.407576102208115|129|1
35.04711|34bd00af7aa3405aa652ce9fda054576c48c9ecd|2.4|2015-01-31 17:47:00|1.4091206135396188|4||129|0.6116874628086298|0|47|523|-80.64817|64|35.04711|FRESH POTATOES|0.0|4|COO RUSSET POTATOES, BULK|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00204072000009|FRESH PRODUCE|PRODUCE|-80.64817|1.407576102208115|129|1
35.04711|5fa9f5dfaa2898cb69ab425e2a170911059b7065|4.49|2014-11-25 15:59:00|1.4091206135396188|4|7203695498|129|0.6116874628086298|0|47|1603|-80.64817|371|35.04711|PRIVATE LABEL BREAD|0.0|14|BAND OF BAKERS RUSSIAN BLACK|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00072036954985|BREAD|BAKERY|-80.64817|1.407576102208115|129|1
35.04711|86874bf6ada52791c55c57e77448d5d4ca2abcc8|1.89|2015-01-18 10:23:00|1.4091206135396188|4|1300079630|129|0.6116874628086298|0|47|69|-80.64817|26|35.04711|CANNED GRAVY|0.0|1|HEINZ GRAVY MUSHROOM HMSTYLE|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00013000798303|PREPARED FOODS-DRY MIXES|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|a80896768c11a9037019171c2508776c4a5f4aa5|3.99|2015-02-22 13:01:00|1.4091206135396188|4|3338324028|129|0.6116874628086298|0|47|504|-80.64817|64|35.04711|FRESH BERRIES|0.99|4|BLACKBERRIES 5.6 OZ|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00881006001099|FRESH PRODUCE|PRODUCE|-80.64817|1.407576102208115|129|1
35.04711|c4a2560626c96fa6395ed1d30b1ea8e6f417edba|7.99|2015-02-19 16:40:00|1.4091206135396188|4|8857333101|129|0.6116874628086298|0|47|458|-80.64817|82|35.04711|CRAFT BEER|0.0|16|SHINER BOCK 6PK|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00088573331011|DOMESTIC BEER|BEER|-80.64817|1.407576102208115|129|1
35.04711|176beccb3dd7e5acd4062fc54ef32db460fade5b|8.99|2015-01-16 15:52:00|1.4091206135396188|4|8857333101|129|0.6116874628086298|0|47|458|-80.64817|82|35.04711|CRAFT BEER|0.0|16|SHINER BOCK 6PK|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00088573331011|DOMESTIC BEER|BEER|-80.64817|1.407576102208115|129|1
35.04711|8f94fcd0bfd638be4af064a8774efea9b5ee7671|8.99|2014-12-08 15:42:00|1.4091206135396188|4|8857333101|129|0.6116874628086298|0|47|458|-80.64817|82|35.04711|CRAFT BEER|0.0|16|SHINER BOCK 6PK|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00088573331011|DOMESTIC BEER|BEER|-80.64817|1.407576102208115|129|1
35.04711|2cbfcffc8e351e33855204631057c0303975227e|8.99|2015-02-09 13:40:00|1.4091206135396188|4|8857333101|129|0.6116874628086298|0|47|458|-80.64817|82|35.04711|CRAFT BEER|0.0|16|SHINER BOCK 6PK|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00088573331011|DOMESTIC BEER|BEER|-80.64817|1.407576102208115|129|1
35.04711|d99e1f058dcbee8a2633c99a191b175e1c1f0370|8.99|2015-01-30 15:15:00|1.4091206135396188|4|8857333101|129|0.6116874628086298|0|47|458|-80.64817|82|35.04711|CRAFT BEER|0.0|16|SHINER BOCK 6PK|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00088573331011|DOMESTIC BEER|BEER|-80.64817|1.407576102208115|129|1
35.04711|707bd7793c9cf2e9cb7bd09d335fca6e004bf761|8.99|2014-12-11 14:55:00|80.648225123995502|4|8857333101|129|35.061235468926334|0|30|458|-80.816172|82|35.059823|CRAFT BEER|0.0|16|SHINER BOCK 6PK|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|35.078006462436761|00088573331011|DOMESTIC BEER|BEER|-80.64817|80.648180832793159|66|1
35.04711|d83cf05756dd499c6e7bdf3312abdfc0e07ff366|0.77|2015-01-20 17:29:00|80.648225123995502|4||129|35.061235467759673|0|30|502|-80.760919|64|35.024332|FRESH BANANAS|0.0|4|BANANAS, YELLOW|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|35.078006462436761|00204011000008|FRESH PRODUCE|PRODUCE|-80.64817|80.648182904778594|343|1
35.04711|0fee21bc93adc9c221fe330770cf9fe59e117c0b|5.99|2014-11-14 17:17:00|1.4091206135396188|4|7756725423|129|0.6116874628086298|0|47|252|-80.64817|45|35.04711|PREMIUM ICE CREAM|1.61|5|BREYERS FRENCH VANILLA I/C|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00077567254382|ICE CREAM|FROZEN|-80.64817|1.407576102208115|129|1
35.04711|aa2abf1982ae9c18dc933f02b508a62b62120762|4.0|2015-02-01 14:03:00|1.4091206135396188|4|89846000211|129|0.6116874628086298|0|47|1165|-80.64817|87|35.04711|NFS-FRESH CONSUMER BUNCH|0.66|9|C 5 ST TULIP BUNCHES|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00898460002111|FLORAL|FLORAL|-80.64817|1.407576102208115|129|1
35.04711|427498577b3d09edaae7f6be5a0eea470dc1a1c4|5.98|2014-12-31 16:15:00|1.4091206135396188|4||129|0.6116874628086298|0|47|528|-80.64817|64|35.04711|FRESH BROCCOLI|0.0|4|BROCCOLINI|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00203277000005|FRESH PRODUCE|PRODUCE|-80.64817|1.407576102208115|129|2
35.04711|b0fc87024e64cdc66995b17553cf7f252a6caf66|3.79|2015-01-31 15:18:00|1.4091206135396188|4|7203688184|129|0.6116874628086298|0|47|555|-80.64817|64|35.04711|PACKAGED SALADS|0.0|4|HTT ASIAN CHOP SALAD KIT|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00072036881847|FRESH PRODUCE|PRODUCE|-80.64817|1.407576102208115|129|1
35.04711|6cac4f81792c998050699817de9789fdef4df959|3.19|2014-12-22 18:07:00|1.4091206135396188|4|2100000730|129|0.6116874628086298|0|47|316|-80.64817|52|35.04711|CREAM CHEESE|0.0|3|PHILLY SOFT CREAM CHEESE|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00021000000142|CHEESE|DAIRY|-80.64817|1.407576102208115|129|1
35.04711|79cb5ce65c3fbdb6b05a2dc463bd7da36c59d4f7|9.99|2014-12-10 15:55:00|1.4091206135396188|4|8143431530|129|0.6116874628086298|0|47|9962|-80.64817|887|35.04711|NFS-PREM-SAUV/FUME'BLANC|0.0|13|CB-NOBILO SAUVIGNON BLANC|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00081434315304|SUPER PREMIUM ($11-$14.99)|WINE|-80.64817|1.407576102208115|129|1
35.04711|979d68964843b0b34d8d43cf8fb42439c5f55c29|0.69|2015-02-03 15:58:00|1.4091206135396188|4||129|0.6116874628086298|0|47|509|-80.64817|64|35.04711|FRESH CITRUS-REMAINING|0.0|4|LEMONS, LARGE|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00204053000004|FRESH PRODUCE|PRODUCE|-80.64817|1.407576102208115|129|1
35.04711|719bd090511f3617aa643b80f13043cf8abac45f|23.92|2014-11-30 11:23:00|1.4091206135396188|4|20201900000|129|0.6116874628086298|0|47|299|-80.64817|49|35.04711|ANGUS BEEF|0.0|2|ANGUS RIBEYE STEAK CUSTOM CUT|ed783c0158bd0e85c2df1de691d9e146f1cae2d7|0.976035983360577|0.61242566243833529|00202019000006|BEEF|MEAT|-80.64817|1.407576102208115|129|2
35.000049|9331f5157ed193ce53245a9d0345f61f55f523dd|2.7|2014-10-14 16:33:00|80.699698036522989|2|4144311023|249|35.025445031998537|0|18|247|-80.760919|39|35.024332|VEGETABLES-FLANKER|0.7|1|M HOLMES SND LIMA BEANS|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00041443119638|VEGETABLES-CAN/JAR|G1 GROCERY|-80.699686|80.699686735047251|343|2
35.000049|42813a4808267ecb2d1c4a8345c2a1c73443a358|5.49|2014-09-10 19:44:00|1.4091206135396188|2|4450020162|249|0.6108660934093487|0|47|847|-80.699686|102|35.000049|NAT/ORG LUNCHMEATS|0.0|19|HF NATURALS SMOKED TURKEY|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00044500201611|LUNCHMEATS|CASE READY MEATS|-80.699686|1.4084752260255726|249|1
35.000049|cccbb9ddb4f0040f72dd96777f02baf54d7b37ff|4.99|2014-10-16 18:48:00|1.4091206135396188|2|3700084603|249|0.6108660934093487|0|47|3530|-80.699686|1045|35.000049|SHAMPOO-MID PRICE|1.0|17|VS SH COLOR PROTECT 25.3 OZ|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00037000846031|HAIR & SCALP CARE|HBC|-80.699686|1.4084752260255726|249|1
35.000049|3b12f8d50f6a7df6a487f556bb4c02aa7ffea9fa|2.59|2014-10-07 22:04:00|1.4091206135396188|2|4369505631|249|0.6108660934093487|0|47|1276|-80.699686|279|35.000049|FROZEN SANDWICHES|0.59|5|LEAN POCKETS SAUSAGE,EGG,CHEES|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00043695062526|FROZEN SANDWICH AND SNACKS|FROZEN|-80.699686|1.4084752260255726|249|1
35.000049|e394423b3166d5b2ac87fb04072b61ab095d6d0c|2.49|2014-12-09 19:04:00|80.699698036522989|2|4369505631|249|35.025445025075619|0|18|1276|-80.758228|279|34.95459|FROZEN SANDWICHES|0.49|5|LEAN POCKETS SAUSAGE,EGG,CHEES|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00043695062526|FROZEN SANDWICH AND SNACKS|FROZEN|-80.699686|80.699708907052567|182|1
35.000049|1ddd60b61ae050c3e4d6da368792ed8f8c8c5149|3.19|2014-11-17 20:43:00|1.4091206135396188|2|4060034500|249|0.6108660934093487|0|47|313|-80.699686|51|35.000049|MARGARINE|1.19|3|ICBINB LIGHT SOFT BOWL|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00040600387187|BUTTER & MARGARINE|DAIRY|-80.699686|1.4084752260255726|249|1
35.000049|0942740f093090198a8d74198e73beba4964e7b5|1.59|2014-10-21 16:23:00|80.699698036522989|2|4650073332|249|35.025445025075619|0|18|393|-80.758228|68|34.95459|NFS-AIR FRESHENERS|0.59|1|GLADE AEROSOL PURE VANILLA|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00046500745393|FRESHENERS/DEODORIZERS|G1 GROCERY|-80.699686|80.699708907052567|182|1
35.000049|0e0f973a95a93d2c2a9d170e211dba7113c37def|6.79|2014-12-28 18:01:00|1.4091206135396188|2|4900002890|249|0.6108660934093487|0|47|54|-80.699686|8|35.000049|DIET|1.8|23|DT SPRITE ZERO 12PK FRIDGEPKCN|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00049000037111|CARBONATED BEVERAGES|BEVERAGE|-80.699686|1.4084752260255726|249|1
35.000049|d15d478480b9a63de73e564e1fea6af1b78d0d95|2.19|2014-11-03 18:39:00|1.4091206135396188|2|5100002549|249|0.6108660934093487|0|47|1221|-80.699686|275|35.000049|PASTA SC VALUE|0.19|1|PREGO SC ALFREDO BACON|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00051000197627|PASTA SAUCES|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|6c2f4b836018fa7c46a515338115b01c1cc7db9e|3.19|2014-11-11 17:48:00|1.4091206135396188|2|5100015339|249|0.6108660934093487|0|47|137|-80.699686|20|35.000049|TOMATO & VEGETABLE JUICE|1.22|1|V8 VFUSION PEACH MANGO|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00051000153418|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|9a1f840702785e4e87fd4909e58c4d096230a75d|2.5|2015-01-20 19:40:00|1.4091206135396188|2|2000019964|249|0.6108660934093487|0|47|1272|-80.699686|50|35.000049|BAG VEG STEAM|0.0|5|GG STEAMERS BROCCOLI FLORETS|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00020000290157|VEGETABLES-FROZEN|FROZEN|-80.699686|1.4084752260255726|249|1
35.000049|1cf5dec9fcaa463a5ee05862439472a70f5c065c|5.69|2014-09-23 17:07:00|1.4091206135396188|2|2220096216|249|0.6108660934093487|0|47|3876|-80.699686|1070|35.000049|SOLID-MALE|2.19|17|GEAR AP FRESH PEAK DEO 2.7|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00022200962131|DEODORANT|HBC|-80.699686|1.4084752260255726|249|1
35.000049|043f263900a871146525a58215b3f94f8a3bac26|2.99|2015-03-09 18:14:00|1.4091206135396188|2|3000004760|249|0.6108660934093487|0|47|60|-80.699686|9|35.000049|HOT CEREAL|1.5|1|QUAKER INST GRITS REAL BUTTER|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00030000037904|CEREAL|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|fece8ffdcbf913ae2bd743e02a2d81aa74ce0456|2.99|2015-02-10 21:07:00|1.4091206135396188|2|3000004760|249|0.6108660934093487|0|47|60|-80.699686|9|35.000049|HOT CEREAL|1.5|1|QUAKER INST GRITS REAL BUTTER|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00030000037904|CEREAL|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|a0943bb72ef206aca4c17d0b7ad47b443790a0b1|4.29|2014-11-15 16:03:00|1.4091206135396188|2|2840015636|249|0.6108660934093487|0|47|204|-80.699686|31|35.000049|TORTILLA CHIPS|1.79|1|DORTIOS NACHO CHEESE|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00028400156363|SNACKS|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|b4cfcdb3b7c3c3044fc1f54008834f93729a316f|7.98|2014-10-14 16:27:00|80.699698036522989|2|7260001894|249|35.025445031998537|0|18|201|-80.760919|31|35.024332|POTATO CHIPS|0.0|1|I/OHERRS CHS BALLS HALLWN 18PK|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00072600018945|SNACKS|G1 GROCERY|-80.699686|80.699686735047251|343|2
35.000049|5fb064873f451349e4e25f757c9950e8d207769a|3.98|2015-01-27 20:20:00|80.699698036522989|2|7940087240|249|35.025445031998537|0|18|726|-80.760919|73|35.024332|NFS-BODY WASHES|0.0|1|SUAVE BW COCOA & SHEA|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00079400602862|PERSONAL SOAP/BATH ADDITIVES|G1 GROCERY|-80.699686|80.699686735047251|343|2
35.000049|50acb74f05229332d4de6d4d267c9a531aab0864|1.99|2015-02-16 16:44:00|80.699698036522989|2|7940087240|249|35.025445025075619|0|18|726|-80.758228|73|34.95459|NFS-BODY WASHES|0.0|1|SUAVE BW COCOA & SHEA|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00079400602862|PERSONAL SOAP/BATH ADDITIVES|G1 GROCERY|-80.699686|80.699708907052567|182|1
35.000049|b89fce5537188d0e3300d2a32ddfc5072ea8669f|3.19|2014-11-02 15:18:00|80.699698036522989|2|7641090137|249|35.025445025075619|0|18|1255|-80.758228|13|34.95459|LUNCH BOX CRACKERS|0.19|1|LANCE TOASTY PEANUT BUTTER 8PK|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00076410901381|CRACKERS|G1 GROCERY|-80.699686|80.699708907052567|182|1
35.000049|3bcd2caf59443a3574ab267613ede69c8c586039|4.99|2014-10-17 14:12:00|80.699698036522989|2|8087804320|249|35.02544503188772|0|18|3601|-80.816172|1050|35.059823|MOUSSE|0.99|17|PANTENE MS FINE VOL TRPL ACT|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00080878043026|HAIR STYLING|HBC|-80.699686|80.699688988521984|66|1
35.000049|18a3ce86c5ce39a0776b391ad31bfcc04dfa7000|3.45|2015-03-03 17:08:00|1.4091206135396188|2|60308421510|249|0.6108660934093487|0|47|3536|-80.699686|1045|35.000049|SHAMPOO-PREMIUM|0.95|17|S/C FRUCTIS BRAZIL SMOOTH SHAM|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00603084433933|HAIR & SCALP CARE|HBC|-80.699686|1.4084752260255726|249|1
35.000049|428693574c59f26b8cf126df639ef72a73656b4f|6.0|2014-12-19 18:19:00|1.4091206135396188|2||249|0.6108660934093487|0|47|512|-80.699686|64|35.000049|FRSH PROD FRSH FRUIT REM|0.0|4|MANGOS|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00204959000009|FRESH PRODUCE|PRODUCE|-80.699686|1.4084752260255726|249|6
35.000049|8c06187a823b9977b3e36c5c4b37f816e51e56a5|2.0|2015-02-25 18:36:00|1.4091206135396188|2||249|0.6108660934093487|0|47|512|-80.699686|64|35.000049|FRSH PROD FRSH FRUIT REM|0.0|4|MANGOS|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00204959000009|FRESH PRODUCE|PRODUCE|-80.699686|1.4084752260255726|249|2
35.000049|cca94901d35d0b77742cd4da33fdd81bccc76e87|3.99|2014-12-02 17:10:00|1.4091206135396188|2|9451441965|249|0.6108660934093487|0|47|389|-80.699686|66|35.000049|NFS-LAUNDRY DETERGENTS|2.0|1|XTRA DETERGENT SENSITVE SCENTS|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00094514428269|DETERGENTS|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|3635282bdb961f0850cf9bb38a83c931a6460a62|5.0|2014-10-02 19:12:00|80.699698036522989|2||249|35.025445031998537|0|18|512|-80.760919|64|35.024332|FRSH PROD FRSH FRUIT REM|0.0|4|MANGOS|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00204959000009|FRESH PRODUCE|PRODUCE|-80.699686|80.699686735047251|343|5
35.000049|8b76bf78222f9f275a3aef07c7da1c10de0e2d1d|2.79|2014-12-19 16:32:00|80.699698036522989|2|76172020560|249|35.025445025075619|0|18|192|-80.758228|30|34.95459|COOKING SPRAYS|0.4|1|MAZOLA BUTTER COOKING SPRAY|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00761720205501|SHORTENING/OIL|G1 GROCERY|-80.699686|80.699708907052567|182|1
35.000049|070b5d97e522865ff85add3d54b1c997a2467d4d|2.79|2014-10-19 19:19:00|1.4091206135396188|2|76172020560|249|0.6108660934093487|0|47|192|-80.699686|30|35.000049|COOKING SPRAYS|0.0|1|MAZOLA BUTTER COOKING SPRAY|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00761720205501|SHORTENING/OIL|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|b9c1623e2f0cb4049f635b6987701c29507cc724|2.99|2014-10-28 16:29:00|80.699698036522989|2|70601011292|249|35.025445031331081|0|18|1219|-80.770346|275|35.052812|PASTA SC CORE|0.0|1|BARILLA SC MARINARA|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00706010112923|PASTA SAUCES|G1 GROCERY|-80.699686|80.69969314690799|40|1
35.000049|7c235d82b327d1c05eeff60d800235362791541d|2.19|2014-09-12 15:46:00|1.4091206135396188|2|3760003895|249|0.6108660934093487|0|47|659|-80.699686|103|35.000049|CHILDRENS LUNCH SNACKS|0.19|19|HORMEL REV BACON CLUB|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00037600207706|LUNCH SNACKS|CASE READY MEATS|-80.699686|1.4084752260255726|249|1
35.000049|5801d694260f59c898d5ae645c244dc39990de75|3.58|2014-11-25 18:49:00|80.699698036522989|2|4100000362|249|35.025445025075619|0|18|213|-80.758228|33|34.95459|SOUP MIXES|0.58|1|LIPTON ONION SOUP & DIP MIX|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00041000003622|SOUP|G1 GROCERY|-80.699686|80.699708907052567|182|2
35.000049|7cac7dfb091b14f47c36da820bb7f27c15676e2d|4.89|2014-10-15 16:51:00|80.699698036522989|2|3700084609|249|35.025445025075619|0|18|3592|-80.758228|1050|34.95459|HAIR STYLING HAIR SPRAY|1.4|17|VS FLEXIBLE HOLD HAIR SPRAY|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00037000846925|HAIR STYLING|HBC|-80.699686|80.699708907052567|182|1
35.000049|c428446f25a6f8e478742498fab827beb24be77d|11.98|2014-10-20 16:02:00|80.699698036522989|2|3700050954|249|35.025445025075619|0|18|1513|-80.758228|66|34.95459|NFS-LAUNDRY DETERGENT PODS|2.0|1|GAIN FLINGS MB 16CT|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00037000867517|DETERGENTS|G1 GROCERY|-80.699686|80.699708907052567|182|2
35.000049|1760f66279e7b7c5c8a66be6cc2bcf6283fe4c15|2.67|2014-09-14 17:07:00|1.4091206135396188|2|7203670830|249|0.6108660934093487|0|47|31|-80.699686|4|35.000049|NON CARBONATED WATER|0.0|1|(U)HT PURIFIED WATER .5L 32 PK|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00072036708304|BOTTLED WATER|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|bd0cc2aa1782e41c117e121dd8f6f4d673c024b1|1.79|2014-09-30 18:20:00|80.699698036522989|2|7239231921|249|35.025445025345761|0|18|209|-80.64817|20|35.04711|POWDERED SOFT DRINKS|0.9|1|HAWIAN SNG TO GO LEMON BRY SQZ|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00072392319244|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.699686|80.699708456151342|129|1
35.000049|a4c2816f790488447baba2c381bde37fcc194264|2.49|2014-11-28 17:51:00|80.699698036522989|2|7203670604|249|35.025445031998537|0|18|50|-80.760919|7|35.024332|PEG CANDY|0.49|1|HTT CHOC COVER RAISINS|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00072036706010|CANDY|G1 GROCERY|-80.699686|80.699686735047251|343|1
35.000049|a5b8692afbb78f8c3cc3ed9587ca0fcdd5c85e58|3.29|2014-10-21 20:57:00|80.699698036522989|2|7550000520|249|35.025445031998537|0|18|76|-80.760919|11|35.024332|MEAT SAUCES|1.65|1|TEXAS PETE CHA! SRIRACHA|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00075500005206|CONDIMENTS|G1 GROCERY|-80.699686|80.699686735047251|343|1
35.000049|61128237026dab3201e1474a6b344c94db35c3e5|4.99|2015-02-24 18:01:00|1.4091206135396188|2|7418228129|249|0.6108660934093487|0|47|726|-80.699686|73|35.000049|NFS-BODY WASHES|1.49|1|SS SEA KISSED BODYWASH|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00074182282660|PERSONAL SOAP/BATH ADDITIVES|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|f3ae78d3529d8aa0e3bff217bab9b4aa43f84fa0|2.85|2014-11-05 19:46:00|1.4091206135396188|2|8390000536|249|0.6108660934093487|0|47|365|-80.699686|56|35.000049|REFRIGERATED TEAS|0.81|3|GOLD PEAK LEMONADE TEA|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00083900006549|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.699686|1.4084752260255726|249|1
35.000049|5e8d35b09e59e90025a643ec8855df2a8a86a413|2.29|2014-11-12 18:31:00|1.4091206135396188|2|7800023046|249|0.6108660934093487|0|47|54|-80.699686|8|35.000049|DIET|1.29|23|CANADA DRY DT G/ALE 2 LITER|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00078000148466|CARBONATED BEVERAGES|BEVERAGE|-80.699686|1.4084752260255726|249|1
35.000049|104d88fcbf297fef71a71d42607946c5ce239569|2.29|2014-12-21 20:05:00|1.4091206135396188|2|7800023046|249|0.6108660934093487|0|47|54|-80.699686|8|35.000049|DIET|1.29|23|CANADA DRY DT G/ALE 2 LITER|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00078000148466|CARBONATED BEVERAGES|BEVERAGE|-80.699686|1.4084752260255726|249|1
35.000049|74057742a010a13294f68ae4cd5e0aafef30af24|3.29|2015-01-07 18:05:00|80.699698036522989|2|2265530301|249|35.02544503188772|0|18|483|-80.816172|100|35.059823|TURKEY BACON|0.5|19|BUTTERBALL TURKEY BACON|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00022655303015|BACON|CASE READY MEATS|-80.699686|80.699688988521984|66|1
35.000049|7875fb5fdd62a8935759065f082eb85d1c29f46a|2.89|2014-11-26 20:56:00|1.4091206135396188|2|3120000293|249|0.6108660934093487|0|47|116|-80.699686|17|35.000049|DRIED CRANBERRIES|1.45|1|OS CRAISIN POMEGRANATE|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00031200002945|FRUIT-DRIED|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|75466f8a99c096d5d50f475435d94c0979127a2f|7.3|2015-02-11 21:23:00|1.4091206135396188|2|3800059663|249|0.6108660934093487|0|47|61|-80.699686|9|35.000049|RTE CEREAL ADULT|1.82|1|KELLOGG RAISIN BRAN CRUNCH|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00038000870101|CEREAL|G1 GROCERY|-80.699686|1.4084752260255726|249|2
35.000049|e81fd84e2717e3ffe7a88296609d2eb37a67ba84|3.99|2014-12-24 17:12:00|80.699698036522989|2|4400002854|249|35.025445025075619|0|18|1248|-80.758228|12|34.95459|SANDWICH COOKIES|1.49|1|OREO LEMON TWIST|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00044000031015|COOKIES|G1 GROCERY|-80.699686|80.699708907052567|182|1
35.000049|da6148686a7c9e302031aecfa295d62cf8948f6e|1.0|2015-02-03 17:26:00|1.4091206135396188|2|4000000435|249|0.6108660934093487|0|47|47|-80.699686|7|35.000049|REGISTER BARS|0.5|1|(FE)M&M PEANUT CANDY|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00040000000327|CANDY|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|734178a90c2832be9051955f16bbcdc1aa197dee|7.98|2014-10-18 11:48:00|80.699698036522989|2|4000015140|249|35.025445031998537|0|18|46|-80.760919|7|35.024332|PKG CHOC|0.98|1|SNICKERS FUN SIZE|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00040000151401|CANDY|G1 GROCERY|-80.699686|80.699686735047251|343|2
35.000049|e320280d5eb174184c80652983f0971a4e2d2ca8|2.49|2015-03-08 18:49:00|1.4091206135396188|2|7203630050|249|0.6108660934093487|0|47|184|-80.699686|28|35.000049|SALAD DRESSINGS-LIQUID|0.81|1|HT DRS VIN BALSAMIC|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00072036981400|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|0f44cc6e29e1c4fd38fc16f7123dd9e7b657cace|7.98|2014-10-03 18:10:00|1.4091206135396188|2|7203688037|249|0.6108660934093487|0|47|581|-80.699686|136|35.000049|FRESH SALSA|0.0|4|HTT 5 PEPPER SALSA|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00072036880376|OTHER MERCHANDISE|PRODUCE|-80.699686|1.4084752260255726|249|2
35.000049|6dead276010c7d7e30b36acdd25649991d6db021|5.49|2015-02-12 07:31:00|80.699698036522989|2|7203695136|249|35.025444992492012|0|18|1687|-80.70901|385|35.17335|THAW & SELL (SWEET GOODS)|0.0|14|FUDGE ICED BROWNIE|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00072036951359|SWEET GOODS|BAKERY|-80.699686|80.699740698393967|174|1
35.000049|d858272904cd6be5f539962344c00c4311318205|2.49|2015-02-11 19:19:00|80.699698036522989|2|60504939530|249|35.02544503189079|0|18|509|-80.8062|64|35.037115|FRESH CITRUS-REMAINING|0.0|4|LEMONS, SMALL 1LB BAG|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00605049395300|FRESH PRODUCE|PRODUCE|-80.699686|80.699688949322621|27|1
35.000049|2f2dbb0d5889442cae9629441cc8ab22f848be37|2.85|2015-01-12 16:37:00|80.699698036522989|2|4133500053|249|35.025444992492012|0|18|184|-80.70901|28|35.17335|SALAD DRESSINGS-LIQUID|1.43|1|KENS DRS LT VIN BLUE CHEESE|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00041335353683|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.699686|80.699740698393967|174|1
35.000049|62c65c0d672f4ce1bd79246e5212b047c9dce6e6|2.79|2014-11-16 18:50:00|1.4091206135396188|2|7203688211|249|0.6108660934093487|0|47|555|-80.699686|64|35.000049|PACKAGED SALADS|0.0|4|HT PREMIUM ROMAINE|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00072036882110|FRESH PRODUCE|PRODUCE|-80.699686|1.4084752260255726|249|1
35.000049|e8ee6de631b0de30d1175aa5c3d87d8e241543f8|4.97|2014-12-07 19:49:00|1.4091206135396188|2||249|0.6108660934093487|0|47|500|-80.699686|64|35.000049|FRESH APPLES|0.0|4|RED DEL APPLE, WA  48|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00233284000002|FRESH PRODUCE|PRODUCE|-80.699686|1.4084752260255726|249|1
35.000049|f8a5528b72b4824af9828a9e83af155bfe2cd208|4.43|2014-11-25 20:48:00|1.4091206135396188|2||249|0.6108660934093487|0|47|500|-80.699686|64|35.000049|FRESH APPLES|0.0|4|RED DEL APPLE, WA  48|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00233284000002|FRESH PRODUCE|PRODUCE|-80.699686|1.4084752260255726|249|1
35.000049|8f29e72c5c4c6a3a118c7d539c2c5d09d33b296f|5.17|2015-01-13 08:24:00|1.4091206135396188|2||249|0.6108660934093487|0|47|500|-80.699686|64|35.000049|FRESH APPLES|0.0|4|RED DEL APPLE, WA  48|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00233284000002|FRESH PRODUCE|PRODUCE|-80.699686|1.4084752260255726|249|1
35.000049|e3ef422ffa2aaf3ebd7af1ed6c29806fc11da670|5.98|2014-12-13 21:23:00|1.4091206135396188|2|4850002063|249|0.6108660934093487|0|47|365|-80.699686|56|35.000049|REFRIGERATED TEAS|3.0|3|PURE LEAF SWEET TEA|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00048500020630|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.699686|1.4084752260255726|249|2
35.000049|7f01019a190b6b3203af60a89eca873dc8da2b68|3.79|2015-02-20 20:29:00|1.4091206135396188|2|4850002013|249|0.6108660934093487|0|47|335|-80.699686|56|35.000049|ORANGE JUICE-REGRIGERATED|0.79|3|TROPICANA PP ORANGE TANGERINE|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00048500306734|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.699686|1.4084752260255726|249|1
35.000049|28030c55440aa4bd21cc6d04a506aa855d00a566|1.79|2014-10-11 15:44:00|1.4091206135396188|2|5100001047|249|0.6108660934093487|0|47|212|-80.699686|33|35.000049|CONDENSED SOUP|0.0|1|CAMP COND BEEFY MUSHROOM|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00051000017673|SOUP|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|4db9d42446fa9c9ae93d211982574e1ce0d02345|8.97|2014-10-08 15:51:00|1.4091206135396188|2|7172000788|249|0.6108660934093487|0|47|52|-80.699686|7|35.000049|PKG NON CHOC|4.5|1|TOOTSIE CARAMEL APPLE POP|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00071720007884|CANDY|G1 GROCERY|-80.699686|1.4084752260255726|249|3
35.000049|99ae28a95e2fd69965a51134653a5739bf9ab656|2.85|2014-11-05 19:48:00|1.4091206135396188|2|8390000536|249|0.6108660934093487|0|47|365|-80.699686|56|35.000049|REFRIGERATED TEAS|0.81|3|GOLD PEAK RASPBERRY TEA|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00049000063332|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.699686|1.4084752260255726|249|1
35.000049|0068260cc7436ac39c6aaaf6c6be20d03bb9930c|3.34|2014-10-11 17:45:00|80.699698036522989|2|7203643010|249|35.025445025075619|0|18|252|-80.758228|45|34.95459|PREMIUM ICE CREAM|0.84|5|HT PREM COOKIES & CREAM IC|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00072036430229|ICE CREAM|FROZEN|-80.699686|80.699708907052567|182|1
35.000049|7274f194968fed8059aa8dcdb6a39303eebc045f|2.29|2015-01-10 22:20:00|80.699698036522989|2|1800000260|249|35.025445025075619|0|18|325|-80.758228|54|34.95459|BISCUITS-REFRIGERATED|1.29|3|GRANDS FLAKY BISCUITS|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00018000002603|DOUGH PRODUCTS|DAIRY|-80.699686|80.699708907052567|182|1
35.000049|43ba6d242cda140c8bcf6e4a1379b0a6c5d86dcf|4.29|2014-09-16 20:20:00|1.4091206135396188|2|2840015938|249|0.6108660934093487|0|47|201|-80.699686|31|35.000049|POTATO CHIPS|1.79|1|XXL RUFFLES CHED SOUR CREAM|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00028400159609|SNACKS|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|f9d2015eed3d645d6278c79708a5498177ecd62d|6.76|2015-01-24 21:31:00|1.4091206135396188|2|2840005509|249|0.6108660934093487|0|47|201|-80.699686|31|35.000049|POTATO CHIPS|0.82|1|LAYS STAX BBQ|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00028400055109|SNACKS|G1 GROCERY|-80.699686|1.4084752260255726|249|4
35.000049|ffc17dc5b0fb87f14ddb8cc618825a45e34feb86|4.0|2014-11-01 17:27:00|80.699698036522989|2|2700038040|249|35.025445031998537|0|18|257|-80.760919|39|35.024332|TOMATOES|2.0100000000000002|1|D HUNTS STARTER CHILI|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00027000392218|VEGETABLES-CAN/JAR|G1 GROCERY|-80.699686|80.699686735047251|343|3
35.000049|3e4476facf0f9687bfc56c08a7a7d40871d63f28|4.89|2014-10-20 20:46:00|80.699698036522989|2|3700086986|249|35.025445030290072|0|18|3586|-80.771677|1050|35.066546|GELS|1.4|17|VS WAVES TEXTURIZNG GELEE|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00037000869863|HAIR STYLING|HBC|-80.699686|80.699697397476299|45|1
35.000049|5e8850aa4313bcb49147ac9104aedb84d4ecb12d|5.38|2015-03-02 21:21:00|1.4091206135396188|2|1450000253|249|0.6108660934093487|0|47|1272|-80.699686|50|35.000049|BAG VEG STEAM|1.35|5|BE STFRSH BROC/CAUL/CARROTS|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00014500011299|VEGETABLES-FROZEN|FROZEN|-80.699686|1.4084752260255726|249|2
35.000049|fb6a8c0a3f0b5db68d418059e391c14c11f6b5c1|1.89|2014-11-21 16:09:00|80.699698036522989|2|3400000220|249|35.025445025075619|0|18|47|-80.758228|7|34.95459|REGISTER BARS|0.55|1|REESE'S PB CUP KING|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00034000004805|CANDY|G1 GROCERY|-80.699686|80.699708907052567|182|1
35.000049|a2a238ca4a20aafb16e120ce8069bbc0ff80fdec|1.79|2014-10-05 16:16:00|1.4091206135396188|2|5000001011|249|0.6108660934093487|0|47|145|-80.699686|22|35.000049|MILK-CANNED|0.0|1|CARNATION EVAPORATED MILK|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00050000010110|PACKAGED MILKS & MODIFIERS|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|20ab85acfb0943bae728e63b19d8d9e947ba2017|2.99|2014-10-20 19:44:00|1.4091206135396188|2|7073400003|249|0.6108660934093487|0|47|230|-80.699686|37|35.000049|HERBAL TEA|0.49|1|CELESTIAL ZINGER TANGERINE|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00070734053184|TEA|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|9714b752a2f885eaca846a59e84ea3b54c16e1a9|1.69|2014-12-05 14:56:00|80.699698036522989|2|4900000044|249|35.025445025075619|0|18|54|-80.758228|8|34.95459|DIET|0.0|23|CB DIET SPRITE ZERO20OZ|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00049000037197|CARBONATED BEVERAGES|BEVERAGE|-80.699686|80.699708907052567|182|1
35.000049|7877f5a9ad70792b3cdf6e86ea485695a4234a78|4.19|2015-01-13 20:37:00|80.699698036522989|2|60308424372|249|35.025445031998537|0|18|3592|-80.760919|1050|35.024332|HAIR STYLING HAIR SPRAY|1.2|17|S/TFRUCT SLEEK&SHINE FLAT IRON|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00603084223893|HAIR STYLING|HBC|-80.699686|80.699686735047251|343|1
35.000049|5c0aa2d9a0d6b6230710a4560ce2f76bdca9c964|2.99|2015-03-03 20:55:00|80.699698036522989|2|7790047132|249|35.025445031998537|0|18|1271|-80.760919|41|35.024332|PROTEIN BREAKFAST|1.5|5|JIMMY DEAN SAUSAGE BRKFST BOWL|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00077900471322|BREAKFAST FOODS FROZEN|FROZEN|-80.699686|80.699686735047251|343|1
35.000049|430e27816edab3652b3ba85d9dd16dde96d9bab4|5.99|2015-03-08 15:30:00|80.699698036522989|2|76401420805|249|35.025445031998537|0|18|356|-80.760919|104|35.024332|GOURMET SAUSAGE|0.0|19|AIDELLS ITALIAN MOZZARELLA|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00764014293529|DINNER SAUSAGE|CASE READY MEATS|-80.699686|80.699686735047251|343|1
35.000049|fc13c8239e0d40274674680e54e6c8c90eed695c|4.23|2015-02-10 17:09:00|1.4091206135396188|2||249|0.6108660934093487|0|47|529|-80.699686|64|35.000049|FRESH ASPARAGUS|1.06|4|GREEN  ASPARAGUS|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00204080000008|FRESH PRODUCE|PRODUCE|-80.699686|1.4084752260255726|249|1
35.000049|0ee77935e5606ac1dbeee56358c2e328be01a03b|4.9|2014-11-02 15:13:00|80.699698036522989|2||249|35.025445031998537|0|18|500|-80.760919|64|35.024332|FRESH APPLES|0.0|4|RED DEL APPLES, WA  72|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00204016000003|FRESH PRODUCE|PRODUCE|-80.699686|80.699686735047251|343|1
35.000049|fc0f0bb4c1f38debee569e04d9e1e47a246f99eb|9.14|2015-03-09 19:36:00|1.4091206135396188|2||249|0.6108660934093487|0|47|503|-80.699686|64|35.000049|FRESH GRAPES|5.24|4|RED GRAPES,SEEDLESS 12/16|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00204023000003|FRESH PRODUCE|PRODUCE|-80.699686|1.4084752260255726|249|1
35.000049|3c95d29a49e1372e4ff48a2497097f484ccbcec9|12.58|2015-01-10 14:26:00|1.4091206135396188|2|38137003342|249|0.6108660934093487|0|47|3237|-80.699686|1020|35.000049|ACNE PRODUCTS|0.0|17|CLN&CLEAR DEEP ACT CLNSG SCRUB|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00381370019367|FACIAL CLEANSER & MOISTURIZER|HBC|-80.699686|1.4084752260255726|249|2
35.000049|04e4f46f2a83cb588b794af3613da53e491d365b|1.94|2014-12-24 18:40:00|1.4091206135396188|2|4300020431|249|0.6108660934093487|0|47|94|-80.699686|14|35.000049|PUDDING MIXES|0.22|1|JELLO INST PUDDING LEMON|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00043000204405|DESSERTS/GELS/SYRUPS|G1 GROCERY|-80.699686|1.4084752260255726|249|2
35.000049|bb62adca159b7c49a7446e6e0fa0b946e7f1156e|1.59|2015-01-07 16:20:00|1.4091206135396188|2|2200000512|249|0.6108660934093487|0|47|48|-80.699686|7|35.000049|REGISTER GUM|0.0|1|(FE) 5 RPM MINT GUM 15 PC|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00022000014719|CANDY|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|d3e38f92d44c67813b9a24dbe4d86d7b00bf8a0a|5.94|2014-09-27 08:36:00|80.699698036522989|2|3400000031|249|35.02544503189079|0|18|47|-80.8062|7|35.037115|REGISTER BARS|0.5|1|HERSHEY MILK CHOC BAR|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00034000002405|CANDY|G1 GROCERY|-80.699686|80.699688949322621|27|6
35.000049|69b7773a51035751d69e3a67b97a1489ffe5fa78|8.99|2014-12-21 19:59:00|1.4091206135396188|2|7069002336|249|0.6108660934093487|0|47|757|-80.699686|3|35.000049|BAKING NUTS|3.0|1|FISHER PECAN HALVES|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00070690023344|BAKING SUPPLIES|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|d929bb9501db0b5c12754ab4d4d5ca2ad7e92c08|1.39|2014-12-11 16:27:00|1.4091206135396188|2|1254667609|249|0.6108660934093487|0|47|48|-80.699686|7|35.000049|REGISTER GUM|0.14|1|TRIDENT WHITE PEPPERMINT|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00012546676090|CANDY|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|92dcbb158eeb3ca3e56cffc1806ef801399d8f1e|3.19|2014-10-10 19:49:00|1.4091206135396188|2|2073509275|249|0.6108660934093487|0|47|365|-80.699686|56|35.000049|REFRIGERATED TEAS|1.19|3|TURKEY HILL PEACH TEA|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|0.61242566243833529|00020735096338|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.699686|1.4084752260255726|249|1
35.000049|5cf89f814fbcf5726f0c49060eec40dd844aa3f7|4.49|2014-10-20 20:13:00|80.699698036522989|2|2840023847|249|35.025445031331081|0|18|201|-80.770346|31|35.052812|POTATO CHIPS|0.5|1|DORITOS MINIS VARIETY 10  CT|edeae3ece521016ca1bd3b1c73100be3baaaaba0|1.754804482370625|35.030887098939942|00028400238472|SNACKS|G1 GROCERY|-80.699686|80.69969314690799|40|1
35.17335|21938ca7d7bdf00e12bc6ef48e113e347ccd4602|2.99|2015-01-03 17:41:00|80.728244613218536|2|3338365583|174|35.278508321469332|0|5|522|-81.027334|64|34.977331|FRESH TOMATOES|0.2|4|SWEET GRAPE TOMATO (PINT)|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00072036880284|FRESH PRODUCE|PRODUCE|-80.70901|80.709457905536979|149|1
35.17335|23b3b78ef48ed0bda037bf3e175cd44cfcca8814|5.99|2014-10-25 16:49:00|80.728244613218536|2|7203688216|174|35.278508321469332|0|5|500|-81.027334|64|34.977331|FRESH APPLES|0.0|4|HT HONEYCRISP APPLE 3LB|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00072036882165|FRESH PRODUCE|PRODUCE|-80.70901|80.709457905536979|149|1
35.17335|2ae28d932e3416859332515821f77ee1a618877a|2.99|2014-09-13 13:01:00|80.728244613218536|2|3338365583|174|35.278508321469332|0|5|522|-81.027334|64|34.977331|FRESH TOMATOES|0.49|4|SWEET GRAPE TOMATO (PINT)|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00072036880284|FRESH PRODUCE|PRODUCE|-80.70901|80.709457905536979|149|1
35.17335|8597488c4e233195c56fee95864a41720026eb67|1.99|2015-01-10 18:20:00|80.728244613218536|2|4800000095|174|35.278508321469332|0|5|190|-81.027334|29|34.977331|TUNA-CANNED|0.49|1|COS TUNA SOLID WHITE ALB|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00048000000958|SEAFOOD-CANNED|G1 GROCERY|-80.70901|80.709457905536979|149|1
35.17335|96676c70d0414e7abbf7a5b1d351b87b8fb34dbf|4.99|2014-12-20 19:13:00|80.728244613218536|2|5000031474|174|35.278508321469332|0|5|144|-81.027334|229|34.977331|CEAMERS-POWDERED|0.0|1|COFFEE MATE SWEET ORIG PWDR|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00050000525171|COCOAS CREAMERS SYRUPS|G1 GROCERY|-80.70901|80.709457905536979|149|1
35.17335|cda007d32b7915b47c4581ce4b832e98c6f5415d|3.89|2014-11-01 16:53:00|80.728244613218536|2|4800009030|174|35.278508321469332|0|5|190|-81.027334|29|34.977331|TUNA-CANNED|0.39|1|C0S TUNA 3PK SOLID WHITE ALB|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00048000090300|SEAFOOD-CANNED|G1 GROCERY|-80.70901|80.709457905536979|149|1
35.17335|1d23be8ead11ecb53f004e45ab7f16c186e48b10|1.17|2014-09-26 19:40:00|80.728244613218536|2|7203690021|174|35.278508321469332|0|5|1033|-81.027334|163|34.977331|HAMBURGER|0.0|7|H T HAMBURGER BUNS|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00072036900210|BUNS/ROLLS|COMMERCIAL BAKERY|-80.70901|80.709457905536979|149|1
35.17335|f65b1e9e56aa730e75d21bc3429646d7944ff04a|1.17|2014-11-29 16:38:00|80.728244613218536|2|7203690021|174|35.278508321469332|0|5|1033|-81.027334|163|34.977331|HAMBURGER|0.0|7|H T HAMBURGER BUNS|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00072036900210|BUNS/ROLLS|COMMERCIAL BAKERY|-80.70901|80.709457905536979|149|1
35.17335|d6be0fe2f2d2fd3b895c9c8463df26f573f82266|1.17|2014-10-18 17:39:00|80.728244613218536|2|7203690021|174|35.278508321469332|0|5|1033|-81.027334|163|34.977331|HAMBURGER|0.0|7|H T HAMBURGER BUNS|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00072036900210|BUNS/ROLLS|COMMERCIAL BAKERY|-80.70901|80.709457905536979|149|1
35.17335|0a412e7b40e79d802844f0476c77699543c4757a|3.69|2014-09-21 19:06:00|80.728244613218536|2|7203670310|174|35.278508321469332|0|5|728|-81.027334|72|34.977331|NFS-PLASTIC FLATWARE|0.0|1|"YH 10"" FLEX NEON STRAWS"|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00072036703101|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.70901|80.709457905536979|149|1
35.17335|d658936d2bd47a23d6fe88d502a4b32e216100c3|5.99|2015-02-14 17:41:00|80.728244613218536|2|76108880157|174|35.278508321469332|0|5|1939|-81.027334|465|34.977331|COLD PREP FOODS SIDES|0.0|6|YUKON GOLD MASHED POTATOES|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00761088801575|COLD PREPARED FOODS|DELI|-80.70901|80.709457905536979|149|1
35.17335|9794e911b0e41819424218fb8b47199e2e98f55c|3.78|2014-10-04 17:47:00|80.728244613218536|2|73639310343|174|35.278508321469332|0|5|247|-81.027334|39|34.977331|VEGETABLES-FLANKER|0.0|1|GLORY SND GREEN BEANS|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00736393709137|VEGETABLES-CAN/JAR|G1 GROCERY|-80.70901|80.709457905536979|149|2
35.17335|63dc41683c070e49b12d73d3ad6708f125d0ca69|1.19|2014-12-27 15:35:00|80.728244613218536|2|88439506101|174|35.278508321469332|0|5|242|-81.027334|39|34.977331|CANNED BEANS|0.6|1|LUCKS BEAN PINTO|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00884395061019|VEGETABLES-CAN/JAR|G1 GROCERY|-80.70901|80.709457905536979|149|1
35.17335|9367b5a67185fa8a60715005c9830b8792d5f71f|3.99|2014-11-15 18:15:00|80.728244613218536|2|7127927100|174|35.278508321469332|0|5|555|-81.027334|64|34.977331|PACKAGED SALADS|0.0|4|F.E. BABY SPINACH|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00071279271002|FRESH PRODUCE|PRODUCE|-80.70901|80.709457905536979|149|1
35.17335|82b61ab6defe537c53fbdeb9d08b8fc153b63f19|3.49|2015-03-07 16:14:00|80.728244613218536|2|3800080681|174|35.278508321469332|0|5|60|-81.027334|9|34.977331|HOT CEREAL|0.0|1|SPEC K NOURISH MAPLE B S CRUNH|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00038000806667|CEREAL|G1 GROCERY|-80.70901|80.709457905536979|149|1
35.17335|2a65bb7eadef373134e0dfbf7954c2af2fdf289e|2.39|2014-12-08 18:50:00|80.728244613218536|2|4127102562|174|35.278508321469332|0|5|341|-81.027334|57|34.977331|CREAMERS|0.0|3|ITNAT'L FF/SF CARM MARSHMALLOW|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00041271022513|MILK|DAIRY|-80.70901|80.709457905536979|149|1
35.17335|55fbadad6a7f4f3a27912387dcdd039f97059a82|4.19|2014-10-11 15:32:00|80.728244613218536|2|4812127620|174|35.278508321469332|0|5|1037|-81.027334|164|34.977331|ENGLISH MUFFINS|2.1|7|THOMAS LITE MULTIGRAIN EM PP|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00048121276201|BREAKFAST|COMMERCIAL BAKERY|-80.70901|80.709457905536979|149|1
35.17335|333aab20051b0257fc41a11f14993d9e26202857|2.98|2015-02-21 16:31:00|80.728244613218536|2|5000000457|174|35.278508321469332|0|5|168|-81.027334|24|34.977331|NFS-CAT TREATS|0.48|1|FF APPETIZER CHICKEN & TUNA|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00050000004683|PET FOOD/SUPPLIES|G1 GROCERY|-80.70901|80.709457905536979|149|2
35.17335|e17ba12abfa60dfa8e8036858d0b0a88592af05f|2.5|2014-11-09 16:11:00|80.728244613218536|2|5000029089|174|35.278508321469332|0|5|154|-81.027334|24|34.977331|NFS-CAT FOOD WET|0.0|1|FF BROTHS TUNA,WHTFSH&ANCHOVIE|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00050000291090|PET FOOD/SUPPLIES|G1 GROCERY|-80.70901|80.709457905536979|149|2
35.17335|1052b1f099c7dbed92b69e2a8f6000fd6e696616|6.98|2015-01-19 14:37:00|80.728244613218536|2|7641090137|174|35.278508321469332|0|5|1255|-81.027334|13|34.977331|LUNCH BOX CRACKERS|1.74|1|LANCE R/F TOASTCHEESE|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00076410523330|CRACKERS|G1 GROCERY|-80.70901|80.709457905536979|149|2
35.17335|f320407768ff43325cec62c39f82a98da6cc3256|4.85|2014-12-23 21:17:00|80.728244613218536|2|7790011553|174|35.278508321469332|0|5|361|-81.027334|105|34.977331|BREAKFAST SAUSAGE|1.51|19|JIMMY DEAN SAGE SAUSAGE|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00077900116339|BREAKFAST SAUSAGE|CASE READY MEATS|-80.70901|80.709457905536979|149|1
35.17335|ccea704cd6cc7be0bc2cf81a7055ed5a64ac9adf|3.59|2015-02-03 17:19:00|80.728244613218536|2|7353000003|174|35.278508321469332|0|5|68|-81.027334|11|34.977331|BARBECUE SAUCES|0.0|1|CAROLINA TREET BBQ SAUCE|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00073530000031|CONDIMENTS|G1 GROCERY|-80.70901|80.709457905536979|149|1
35.17335|68c822b3223c9a934bea0b33a1d0d621fa5b1920|2.99|2014-11-19 19:17:00|80.728244613218536|2|7203663104|174|35.278508321469332|0|5|364|-81.027334|55|34.977331|ORGANIC AND CF EGGS|0.0|3|HTN NEST GRADE A LARGE EGG BRO|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00072036631046|EGGS FRESH|DAIRY|-80.70901|80.709457905536979|149|1
35.17335|1377a7cb98b6afdd804db092c00462bcb69dd73c|3.99|2014-11-07 17:45:00|80.728244613218536|2|7976503272|174|35.278508954234148|0|5|31|-80.654118|4|35.123768|NON CARBONATED WATER|2.0|1|CRYSTAL SPRINGS .5 LT 12 PACK|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00079765032724|BOTTLED WATER|G1 GROCERY|-80.70901|80.709044444921375|473|1
35.17335|bd74e877f33119fb05a2d6d547934a026bb6f1f7|7.29|2015-01-17 16:51:00|80.728244613218536|2||174|35.278508321469332|0|5|503|-81.027334|64|34.977331|FRESH GRAPES|1.04|4|RED GRAPES,SEEDLESS 12/16|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00204023000003|FRESH PRODUCE|PRODUCE|-80.70901|80.709457905536979|149|1
35.17335|7e4badea676340b201c057c0fe50e0f8b8f0e110|10.94|2014-11-10 12:16:00|80.728244613218536|2|2550000367|174|35.278508321469332|0|5|66|-81.027334|10|34.977331|GROUND CAN|0.0|1|FOLGERS SPECIAL ROAST|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00025500900308|COFFEE|G1 GROCERY|-80.70901|80.709457905536979|149|2
35.17335|414579d828012cec556db3368a0692ba1a98930d|3.49|2014-12-24 18:12:00|80.728244613218536|2|2500004786|174|35.278508321469332|0|5|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.5|3|MINUTE MAID LOW ACID|f3d64954a3429e9105f76af02286f11e3cb79828|7.266230047906999|35.296297200616316|00025000047985|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.70901|80.709457905536979|149|1
35.297134|146bf3ffc31b128e9aa3fc062053c4d94e5fac24|2.69|2014-11-11 17:29:00|80.728244613218536|4|2700039023|258|35.307113336561528|0|5|257|-80.66939|39|35.28326|TOMATOES|0.0|1|HUNTS TOMATO SAUCE 29|f488fabfaa44bf761e3a81b1771b166ff662158a|0.6895480667870099|35.296297200616316|00027000390238|VEGETABLES-CAN/JAR|G1 GROCERY|-80.737839|80.737841042540936|46|1
35.297134|294069e0839fa8262f2974b24a1aac1f8e2143bc|4.99|2015-02-16 18:24:00|80.728244613218536|4|4900005235|258|35.307113336561528|0|5|55|-80.66939|8|35.28326|REGULAR|1.0|23|DT DR PEPPER  7.5 OZ 8PK|f488fabfaa44bf761e3a81b1771b166ff662158a|0.6895480667870099|35.296297200616316|00078000009729|CARBONATED BEVERAGES|BEVERAGE|-80.737839|80.737841042540936|46|1
35.297134|006774bcc5048c0e4c5eb50d9fc83ea6114f4d1e|16.17|2015-02-15 11:14:00|80.728244613218536|4|20229500000|258|35.307113336561528|0|5|299|-80.66939|49|35.28326|ANGUS BEEF|0.0|2|ANGUS BEEF EYE OF ROUND ROAST|f488fabfaa44bf761e3a81b1771b166ff662158a|0.6895480667870099|35.296297200616316|00202295000004|BEEF|MEAT|-80.737839|80.737841042540936|46|1
35.43259|a77d763d70ec1896a315ada06340d4dc33649a39|0.97|2015-02-04 21:28:00|1.4057311447477159|4|7203671102|202|0.6184153580092175|0|52|1025|-80.605588|162|35.43259|WHITE|0.0|7|HT OLD FASHIONED BREAD|fc1456ee62e52c903a8b11e08eb708a7104187db|0.4435307800413147|0.6209993146566879|00072036711021|SLICED BREAD|COMMERCIAL BAKERY|-80.605588|1.406832906106031|202|1
35.43259|d7293ff25b33b71abd9e1ac64d7be1df8757b43a|5.34|2015-01-31 18:06:00|1.4057311447477159|4|20165700000|202|0.6184153580092175|0|52|297|-80.605588|49|35.43259|GROUND BEEF|1.19|2|HT GROUND BEEF CHUCK 80% LEAN|fc1456ee62e52c903a8b11e08eb708a7104187db|0.4435307800413147|0.6209993146566879|00201657000003|BEEF|MEAT|-80.605588|1.406832906106031|202|1
35.219587|ddffea148ed5b46ea5006fc085a826893d83ed7f|5.99|2015-02-16 17:23:00|80.810069425230125|4|7756725423|401|35.235071766875151|0|23|252|-80.826724|45|35.195689|PREMIUM ICE CREAM|2.99|5|BREYERS BUTTER PECAN I/C|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00077567254405|ICE CREAM|FROZEN|-80.810056|80.81006214331299|412|1
35.219587|d215a57affada6b76cb479e0182f6e773d0f6d80|1.29|2014-10-29 12:55:00|1.4094857484078087|4|8379152001|401|0.6146977543425921|0|26|1981|-80.810056|480|35.219587|CHIPS|0.0|6|DIRTY POTATO CHIP BBQ|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|0.61471665291522548|00083791520049|DRY GOODS|DELI|-80.810056|1.4104015459209989|401|1
35.219587|b58d13d3d8ef4f6ce9a0ddf2d191f40639ac6a9b|1.29|2014-12-09 12:47:00|80.810069425230125|4|8379152001|401|35.235071766875151|0|23|1981|-80.826724|480|35.195689|CHIPS|0.18|6|DIRTY POTATO CHIP BBQ|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00083791520049|DRY GOODS|DELI|-80.810056|80.81006214331299|412|1
35.219587|db6f4209f3f8927a2682ebdcb50385d94b9cf137|3.59|2014-10-01 14:06:00|1.4094857484078087|4|7641090137|401|0.6146977543425921|0|26|1252|-80.810056|12|35.219587|LUNCH BOX COOKIES|1.09|1|LANCE NEKOT CHOCOLATE FILLING|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|0.61471665291522548|00076410901114|COOKIES|G1 GROCERY|-80.810056|1.4104015459209989|401|1
35.219587|1559976dc109ffe9c601f8dcf84b594ea55cae14|9.75|2014-12-11 14:51:00|1.4094857484078087|4|7203656080|401|0.6146977543425921|0|26|318|-80.810056|52|35.219587|SHREDDED/GRATED CHEESE|0.66|3|HT SHRED WISC XTRA SHARP CHED|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|0.61471665291522548|00072036705181|CHEESE|DAIRY|-80.810056|1.4104015459209989|401|3
35.219587|bca299c6e6b574d1bbcc5ef0b1b34d3a9803d384|4.29|2015-01-04 14:37:00|1.4094857484078087|4|2840016014|401|0.6146977543425921|0|26|201|-80.810056|31|35.219587|POTATO CHIPS|2.15|1|LAYS CLASSIC|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|0.61471665291522548|00028400160148|SNACKS|G1 GROCERY|-80.810056|1.4104015459209989|401|1
35.219587|bc4fc563860e184abca7955cca0ba5cb3df5454b|5.94|2015-01-11 16:35:00|80.810069425230125|4|7203619046|401|35.235071766875151|0|23|122|-80.826724|19|35.195689|HONEY|0.72|1|E  HT PURE HONEY BEAR|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00072036190468|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.810056|80.81006214331299|412|2
35.219587|eaa38f6a0a9bf5a5c0d9ffb84bc1700959676eca|4.0|2015-02-16 17:21:00|80.810069425230125|4|5100000524|401|35.235071766875151|0|23|1201|-80.826724|33|35.195689|RTS CANNED|0.0|1|CHUNKY HR SIRLOIN BURGER|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00051000180346|SOUP|G1 GROCERY|-80.810056|80.81006214331299|412|2
35.219587|206dd10fbef5893ba361a82585f6019ae25ba059|15.86|2015-01-10 16:17:00|80.810069425230125|4|20165700000|401|35.235071766875151|0|23|297|-80.826724|49|35.195689|GROUND BEEF|0.0|2|HT GROUND BEEF CHUCK 80% LEAN|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00201657000003|BEEF|MEAT|-80.810056|80.81006214331299|412|8
35.219587|c2c1454326e3593b543017b437c3dfa1f4cf61c2|4.99|2015-02-22 16:29:00|80.810069425230125|4|7203688077|401|35.235071766875151|0|23|523|-80.826724|64|35.195689|FRESH POTATOES|0.0|4|HT RED POTATO 5LB BAG|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00072036880772|FRESH PRODUCE|PRODUCE|-80.810056|80.81006214331299|412|1
35.219587|92557b7d17fbdd641608e188b8ca7fb7a6f6c6e1|3.79|2015-02-10 14:05:00|1.4094857484078087|4|7203688014|401|0.6146977543425921|0|26|581|-80.810056|136|35.219587|FRESH SALSA|2.06|4|HT FRESH MEDIUM SALSA|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|0.61471665291522548|00072036880222|OTHER MERCHANDISE|PRODUCE|-80.810056|1.4104015459209989|401|1
35.219587|f6c5ad4f5bee90eeedc015ec6b058870f3a47e15|7.49|2015-01-07 17:11:00|80.810069425230125|4|4300079460|401|35.235071766875151|0|23|67|-80.826724|10|35.195689|SOLUBLE INSTANT|0.0|1|MAXWELL HOUSE INSTANT COFFEE|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00043000794609|COFFEE|G1 GROCERY|-80.810056|80.81006214331299|412|1
35.219587|123633bbedecb43e090e903a1c908d8793c1e431|7.49|2015-02-06 16:12:00|80.810069425230125|4|4300079460|401|35.235071766875151|0|23|67|-80.826724|10|35.195689|SOLUBLE INSTANT|0.0|1|MAXWELL HOUSE INSTANT COFFEE|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00043000794609|COFFEE|G1 GROCERY|-80.810056|80.81006214331299|412|1
35.219587|93c5e4e7828695e8e2feb6a3ba084c6b8c069795|7.94|2014-10-21 11:37:00|1.4094857484078087|4|5400011971|401|0.6146977543425921|0|26|427|-80.810056|72|35.219587|NFS-TOILET TISSUE|0.0|1|SCOTT 1000 WHITE 8 ROLL|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|0.61471665291522548|00054000119712|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.810056|1.4104015459209989|401|2
35.219587|c71e9313843b981c72f2a9866c44e26ee8d78229|2.59|2014-12-01 18:41:00|80.810069425230125|4|7203663996|401|35.235071766875151|0|23|342|-80.826724|57|35.195689|FRESH MILK|0.26|3|HARRIS TEETER WHOLE MILK|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00072036639967|MILK|DAIRY|-80.810056|80.81006214331299|412|1
35.219587|706700f4e9d4bf28c46c1f1cb759334ae2fbb378|4.29|2014-12-07 20:04:00|80.810069425230125|4|2840016014|401|35.235071766449451|0|23|201|-80.80146|31|35.17739|POTATO CHIPS|0.29|1|LAYS BBQ|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00028400160131|SNACKS|G1 GROCERY|-80.810056|80.810063582707045|208|1
35.219587|f7aefc3dbee72d74f6f5177b82648e94609c7da2|4.29|2014-11-21 19:58:00|1.4094857484078087|4|2840016014|401|0.6146977543425921|0|26|201|-80.810056|31|35.219587|POTATO CHIPS|2.15|1|LAYS DILL PICKLE|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|0.61471665291522548|00028400160285|SNACKS|G1 GROCERY|-80.810056|1.4104015459209989|401|1
35.219587|033a05a030b36fa44ce9c00f67e2ae7657f05ed1|1.49|2014-10-25 11:57:00|80.810069425230125|4|2840002819|401|35.235071766875151|0|23|206|-80.826724|31|35.195689|FRONT END SNACKS|0.0|1|LAYS CLASSIC|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00028400027960|SNACKS|G1 GROCERY|-80.810056|80.81006214331299|412|1
35.219587|6af1d0483ff4572a2cbda86686000370acea7b69|1.49|2015-01-16 16:20:00|80.810069425230125|4|2840002819|401|35.235071766875151|0|23|206|-80.826724|31|35.195689|FRONT END SNACKS|0.0|1|LAYS CLASSIC|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00028400027960|SNACKS|G1 GROCERY|-80.810056|80.81006214331299|412|1
35.219587|14551ac034c284b6644831f10cbf2592e62064ca|1.49|2015-01-17 19:09:00|80.810069425230125|4|2840002819|401|35.235071766875151|0|23|206|-80.826724|31|35.195689|FRONT END SNACKS|0.0|1|LAYS CLASSIC|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00028400027960|SNACKS|G1 GROCERY|-80.810056|80.81006214331299|412|1
35.219587|fa7672aad4fae977b1da178c157da38804dd0d55|1.49|2014-12-31 14:13:00|80.810069425230125|4|2840002819|401|35.235071766875151|0|23|206|-80.826724|31|35.195689|FRONT END SNACKS|0.0|1|LAYS CLASSIC|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00028400027960|SNACKS|G1 GROCERY|-80.810056|80.81006214331299|412|1
35.219587|3563519caba432108410d4d4ff76ba084c172c5e|3.98|2014-10-14 23:43:00|80.810069425230125|4|4115289616|401|35.235071766449451|0|23|139|-80.80146|20|35.17739|REMAINING SHELF STABLE JUICES|2.0|1|OASIS BREEZE PINK LEMONADE|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00041152896165|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.810056|80.810063582707045|208|2
35.219587|3723f3dd1207dafd1fd90f18d8af7afcbee46c4a|9.44|2015-02-16 17:45:00|80.810069425230125|4|20596200000|401|35.235071766875151|0|23|1821|-80.826724|410|35.195689|BH TURKEY|1.71|6|BOARS HEAD MAPLE HONEY TURKEY|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00205962000000|BH MEAT|DELI|-80.810056|80.81006214331299|412|1
35.219587|b861eea62bee90c1bfff8b4e01c9c5ca8940694b|11.32|2014-10-08 18:02:00|80.810069425230125|4|20596200000|401|35.235071766875151|0|23|1821|-80.826724|410|35.195689|BH TURKEY|0.0|6|BOARS HEAD MAPLE HONEY TURKEY|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00205962000000|BH MEAT|DELI|-80.810056|80.81006214331299|412|1
35.219587|14868e78e1de119b83143d13ebdad02a2b73d8bd|0.99|2014-12-08 08:46:00|80.810069425230125|4|7203695306|401|35.235071766875151|0|23|1895|-80.826724|450|35.195689|TEA|0.0|6|FFM RASP. LEMONADE|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00072036018922|BEVERAGES|DELI|-80.810056|80.81006214331299|412|1
35.219587|678d649dd62d8a920a9a64c2700abb69bfff7893|0.99|2014-12-10 12:36:00|80.810069425230125|4|7203695306|401|35.235071766875151|0|23|1895|-80.826724|450|35.195689|TEA|0.0|6|FFM RASP. LEMONADE|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00072036018922|BEVERAGES|DELI|-80.810056|80.81006214331299|412|1
35.219587|b02e02692562552dcab615d3ce66f7ac1f8e23a5|0.99|2014-12-10 17:12:00|80.810069425230125|4|7203695306|401|35.235071766875151|0|23|1895|-80.826724|450|35.195689|TEA|0.0|6|FFM HALF TEA/LEMONADE|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00072036018878|BEVERAGES|DELI|-80.810056|80.81006214331299|412|1
35.219587|5e4ad3eb43ecf49b691114aa7aedccb9d54230fe|0.99|2015-01-30 11:26:00|80.810069425230125|4|7203695306|401|35.235071766875151|0|23|1895|-80.826724|450|35.195689|TEA|0.0|6|FFM RASP. LEMONADE|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00072036018922|BEVERAGES|DELI|-80.810056|80.81006214331299|412|1
35.219587|1772cf95510b8b2cd361e5b0db697bbd16b65749|0.99|2015-01-09 11:59:00|80.810069425230125|4|7203695306|401|35.235071766875151|0|23|1895|-80.826724|450|35.195689|TEA|0.0|6|FFM RASP. LEMONADE|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00072036018922|BEVERAGES|DELI|-80.810056|80.81006214331299|412|1
35.219587|1209f9ebdf47f303a19c6f771dd64a8da5990a35|0.99|2015-01-07 15:00:00|80.810069425230125|4|7203695306|401|35.235071766875151|0|23|1895|-80.826724|450|35.195689|TEA|0.0|6|FFM RASP. LEMONADE|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00072036018922|BEVERAGES|DELI|-80.810056|80.81006214331299|412|1
35.219587|8ffe33b7367f6067672c24efe52a7abd6d84bf0c|0.99|2015-02-02 11:57:00|80.810069425230125|4|7203695306|401|35.235071766875151|0|23|1895|-80.826724|450|35.195689|TEA|0.0|6|FFM RASP. LEMONADE|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00072036018922|BEVERAGES|DELI|-80.810056|80.81006214331299|412|1
35.219587|457f24ea1037a55f57538391f9f022bf53e90c76|0.99|2015-01-07 11:24:00|80.810069425230125|4|7203695306|401|35.235071766875151|0|23|1895|-80.826724|450|35.195689|TEA|0.0|6|FFM RASP. LEMONADE|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00072036018922|BEVERAGES|DELI|-80.810056|80.81006214331299|412|1
35.219587|15ea7f892de42aeced34e0811555578daab8868c|0.99|2015-01-28 16:12:00|80.810069425230125|4|7203695306|401|35.235071766875151|0|23|1895|-80.826724|450|35.195689|TEA|0.0|6|FFM RASP. LEMONADE|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00072036018922|BEVERAGES|DELI|-80.810056|80.81006214331299|412|1
35.219587|fa78c65cd5dadec94559282b46533a0c1daa1274|0.99|2015-01-17 13:19:00|80.810069425230125|4|7203695306|401|35.235071766875151|0|23|1895|-80.826724|450|35.195689|TEA|0.0|6|FFM RASP. LEMONADE|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00072036018922|BEVERAGES|DELI|-80.810056|80.81006214331299|412|1
35.219587|25ebbad846e86749a874326e96d5714ab7f660e1|0.99|2015-01-06 13:28:00|80.810069425230125|4|7203695306|401|35.235071766875151|0|23|1895|-80.826724|450|35.195689|TEA|0.0|6|FFM RASP. LEMONADE|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00072036018922|BEVERAGES|DELI|-80.810056|80.81006214331299|412|1
35.219587|cf5bf2477f3115ee31eadf1a1d8e7e05c9b1f1cb|0.58|2014-12-14 16:03:00|80.810069425230125|4|4133507899|401|35.235071766875151|0|23|1984|-80.826724|480|35.195689|PC CONDIMENTS|0.0|6|KEN'S CREAMY RANCH DRESSING|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00041335078999|DRY GOODS|DELI|-80.810056|80.81006214331299|412|2
35.219587|2150e960bf2e5368c4a137761d7974b9834f9aff|5.49|2015-01-14 16:03:00|80.810069425230125|4|7144830025|401|35.235071766875151|0|23|2021|-80.826724|505|35.195689|FRESH CHEESE|0.0|6|ALOUETTE CRANBERRY APPLE|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00071448300823|SPECIALTY CHEESE|DELI|-80.810056|80.81006214331299|412|1
35.219587|bfbcb4852f10e7fd2c1eef7e520b554e3a47b498|11.19|2014-10-21 11:38:00|1.4094857484078087|4|5400010060|401|0.6146977543425921|0|26|427|-80.810056|72|35.219587|NFS-TOILET TISSUE|0.0|1|SCOTT 1000 WHITE 12 ROLL|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|0.61471665291522548|00054000100604|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.810056|1.4104015459209989|401|1
35.219587|f976973ff461294114c27184bd064ad33d463840|2.75|2014-12-09 21:49:00|80.810069425230125|4|5100012573|401|35.235071766875151|0|23|137|-80.826724|20|35.195689|TOMATO & VEGETABLE JUICE|0.56|1|V8 SPLASH TROPICAL BLEND|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00051000125736|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.810056|80.81006214331299|412|1
35.219587|88ace529b6ed867654d7f92659b6c3399c1a6c36|11.67|2014-12-27 17:01:00|80.810069425230125|4|20251400000|401|35.235071766875151|0|23|297|-80.826724|49|35.195689|GROUND BEEF|0.0|2|ANGUS GROUND SIRLOIN|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00202514000006|BEEF|MEAT|-80.810056|80.81006214331299|412|10
35.219587|3c6913b268d8f4f91b71da93ef8e520cf68ac69a|2.0|2014-11-09 15:44:00|80.810069425230125|4|78352032108|401|35.235071766875151|0|23|8598|-80.826724|1792|35.195689|NEWSPAPERS|0.0|18|SUNDAY CHARLOTTE OBSERVER|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00783520321083|NEWSPAPERS|GM|-80.810056|80.81006214331299|412|1
35.219587|348d24623c37d2700efe40596f1256895099112d|1.39|2014-10-09 16:08:00|80.810069425230125|4|1254661959|401|35.235071766875151|0|23|48|-80.826724|7|35.195689|REGISTER GUM|0.39|1|TRIDENT TROPICAL TWIST|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012546619592|CANDY|G1 GROCERY|-80.810056|80.81006214331299|412|1
35.219587|2915daac0aef7732330fc92c53afc0b807b0b653|0.75|2014-11-12 16:24:00|80.810069425230125|4||401|35.235071766875151|0|23|1617|-80.826724|373|35.195689|ROLLS BULK|0.0|14|BULK ROLLS|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00072036955555|ROLLS|BAKERY|-80.810056|80.81006214331299|412|1
35.219587|da143a06880ea1dcc63cfec1bf102922173d9e95|0.75|2015-01-01 15:12:00|80.810069425230125|4||401|35.235071766875151|0|23|1617|-80.826724|373|35.195689|ROLLS BULK|0.0|14|BULK ROLLS|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00072036955555|ROLLS|BAKERY|-80.810056|80.81006214331299|412|1
35.219587|c27a97b946e732d126c3204ae3b3fbf35764d166|0.75|2015-01-26 11:56:00|80.810069425230125|4||401|35.235071766875151|0|23|1617|-80.826724|373|35.195689|ROLLS BULK|0.0|14|BULK ROLLS|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00072036955555|ROLLS|BAKERY|-80.810056|80.81006214331299|412|1
35.219587|211241a83c7020e52189b310dbb089075f44dff3|2.19|2014-10-29 12:32:00|1.4094857484078087|4|1200000230|401|0.6146977543425921|0|26|55|-80.810056|8|35.219587|REGULAR|0.69|23|WILD CHERRY PEPSI 2 LTR|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|0.61471665291522548|00012000003110|CARBONATED BEVERAGES|BEVERAGE|-80.810056|1.4104015459209989|401|1
35.219587|f328ab40426f71273f87bbeadb1483cd2bc40a36|3.99|2014-12-16 06:12:00|80.810069425230125|4|77482603060|401|35.235071766449451|0|23|1656|-80.80146|381|35.17739|CUP CAKES|0.5|14|MINI XMAS VANILLA CUPCAKES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00774826030601|CAKES|BAKERY|-80.810056|80.810063582707045|208|1
35.219587|8a7f8a70214ab21620c8a2d6bebe28fd3072b5ae|1.69|2015-01-13 11:40:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|70aee625fb8203900ba6bcb3b2f6a89d70f0dc96|1.69|2014-10-25 14:11:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|c237941a59b64522af750e330c7a9515c3177898|1.69|2014-10-13 21:47:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|058559a3c993b79bb3cb749f612885127eb53c94|1.69|2015-01-16 13:06:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|0401f1e6f6ef504fe710e27cc6faf3284fc8ecd6|1.69|2014-12-21 12:40:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|c01799bd02b3dc7ba98c4b37d6557d5f9787a523|1.69|2014-12-17 17:09:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|f965ae5a25ef9bd951b3391e99254a2e7ca47b9f|1.69|2015-02-20 14:29:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|609fb8d54bdabdffe1e0d1bc15fe15a0034274ed|1.69|2015-02-07 11:05:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|377eb9178631e006232ac8eacedfea56f41f85f7|1.69|2014-11-05 08:40:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|19763c7cbf4c380bed1352e810c3d6086b7e100c|1.69|2014-10-13 17:28:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|96c0170155657dac213f8ce60a73bb4acb0f07b3|1.69|2015-02-04 14:08:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|bdbc246ee54d2e6111e330024e4849dea8620a49|1.69|2015-01-21 11:47:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|cbd246f7585d1580120d276a251ca0e3723639ce|1.69|2015-02-14 11:58:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|2caeb0d6a426cebadda9eba14e436e4b9e0d2b32|1.69|2014-11-12 12:10:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|4a0b91ba5d65e599b1f1abc59aa16f2c356561e7|1.69|2015-01-05 12:15:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|b080b91f8162ec8ee3dd7739e96b2a0dfcd6080e|1.69|2014-11-25 07:31:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|b47b788678131f15dd3c9b7665f4b9d28b1fef34|1.69|2014-12-01 12:35:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|f6788c8e6117674e2786f810f12507e42cfd32f7|1.69|2014-11-21 11:47:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|274d7414c9022c72dfbc5608ff1ef98680acff82|1.69|2015-02-18 12:08:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|58eb03c6aa42a9912be6711503f990de1b896c80|1.69|2014-11-25 14:55:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|a2dc0a4b60fbdda893ecf8b8de6c81f647809f20|1.69|2014-12-09 17:19:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|0f13514c4c9f1dc8895db3845396f230e555f899|1.69|2015-01-28 12:04:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|3ae6e50b4ad3964836f91b2ca1878e54f1dbeb17|1.69|2014-10-24 13:16:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|f05c5ac2ad6ef89312f17fb0cb6bd52c133dd73a|1.69|2014-10-23 09:35:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|5d122a8c1ca470a84461f28a45985d53e7daa780|1.69|2014-10-03 21:39:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|685179f28b3f9a467bc63afe20fe935cdfd379da|1.69|2014-11-02 12:39:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|b4d73267147df2ec9f970c9928e243eb6bc8af9f|1.69|2014-11-23 17:09:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|62c3e70108a77d7d6b7e4407c37866227be9fbe7|1.69|2015-02-09 14:05:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|7fb705a939f58ed728b337b6537724409a51676e|1.69|2014-11-01 13:03:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|256b9db9de6236100a309a0e62f4fa59460c5c8c|1.69|2014-09-30 12:27:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|21aa2281c285b75a0a602e9a7219de77875e9687|1.69|2014-09-30 14:42:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|a88c93af1ba23448c4aa882fc75003841276d7e2|1.69|2015-01-01 12:48:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|307a5abaac9cc293a29c9ede800296e15e123045|1.69|2014-10-02 09:58:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|aa1f1862c710ed7d102d285aa63b46eca9d0370e|1.69|2015-02-27 12:13:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|2d295d3eef6d5ac74a5040ec4dde52991bdc9baa|1.69|2014-12-27 12:27:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|0555522733ee8538b68f44e74ff89e0056021bd2|1.69|2014-11-08 17:11:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|4bc0b32523195500f0c58b776d276f9deab66920|1.69|2015-01-03 17:37:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|ade69c1dd547cea6ddf6e59a889a10a523cbd299|1.69|2014-12-03 12:47:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|821551695ee763fa90960e6faf1fe6ce50e55be5|1.69|2014-11-29 15:47:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|b87b69994ca1c02b53b02d4398d9db4e2df2bca7|1.69|2015-03-01 14:23:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|c34d3d2f392fb393c41d6018d6dd61fdf11573a3|1.69|2014-12-26 11:58:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|fd92b65adf1437692c526ea5087df4b84a945548|1.69|2014-12-15 15:40:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|23e7ecf639a3404f6b35bf6a5ce3cd4486114a93|1.69|2014-12-12 12:42:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|e18bb72baa2b9c94badd37c6d3ff19cc404a2a29|1.69|2015-01-11 14:18:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|d696249adffc8fa3f4d441691f8082484139f1d9|1.69|2015-02-08 13:46:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|d5b561bd91cc3bf801050006daf672045530f610|1.69|2015-02-11 11:40:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|92c42d2fe3e0694601018277eb36254821899639|1.69|2015-01-19 15:56:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|ed8d6ceaadfc8058470b4c60ade5a10e743e3764|1.69|2014-10-25 09:45:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|ee45833087979d23c860a2a2c9ed08aa46c157ab|1.69|2015-03-04 11:59:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|29d5be3a75ac929be5bd2bdeae628ad06f623927|1.69|2014-10-30 10:48:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|7b4eddd36d044bab921250ae22bc2540c5c0d5b2|1.69|2015-01-25 11:20:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|4f9a3a063f6ece7a6f957ce394b0570bffc6f0ef|1.69|2014-11-26 15:06:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|cb8d64d0bcab964b13817edb70ae62ef17f4485b|1.69|2015-03-02 12:01:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|643e4e9864b5959b810f5f71661f7acd653cc012|1.69|2014-12-07 12:32:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|922aaa898404bba570babc4c3a643b8b6cb93635|1.69|2014-10-15 13:36:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|8fc609166639480ad66d446723ff87c7f4f94580|1.69|2014-12-05 12:30:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|8a65b10b8449b22531f6d8a0f59a80bd6d1a6c93|1.69|2015-02-13 11:39:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|0944d79acfac2047d52e5479f9666d0467cb7fca|1.69|2014-09-20 10:31:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|f242b9dd4ea654940ff511c7723d1bee10615e09|1.69|2015-02-15 11:57:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|165e1f92c3c022bc758d647b0ae62803ebf90acd|3.38|2014-10-03 14:36:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|2
35.219587|53745a7475fc756c9c3ae917092ccbdffc336de6|1.69|2014-11-13 12:45:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|769a7fb4ada8f5cb1ad6f27bc1fdd51b500e9afa|1.69|2015-01-14 14:18:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|76530871d828204825be8e71257c8b8accd9deca|1.69|2014-09-12 14:46:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|f5a4bffe956d76e5acb0696d73462bccd4fc3954|9.58|2014-09-20 14:51:00|80.810069425230125|4|1200010041|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|4.8|23|MTN DEW 16 OZ 6 PK|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000100710|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|2
35.219587|4ed9c1b11cafac2fc8a564bf09c8d027ed77bcca|1.69|2015-01-23 16:15:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|cbb5a78058d162f6de769adf09a21b1d4b36c5c2|1.69|2014-11-14 13:23:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|cae7c56a32f259d56f25c67667a68f8d886cc3f5|1.69|2015-01-09 14:59:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|1a6a374a6c6117518f5326a67ac1f738e166510e|1.69|2015-01-03 08:41:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|f846bb9c5bbc6b241e7250a73ddf1a58172210f7|1.69|2015-01-10 12:17:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|957c4d9cb1595ec026a61d97387632e0f9cdd245|1.69|2014-11-30 14:44:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|51d2884a97460c41cc1e3664827bb5b9f5f389fb|1.69|2014-12-24 14:24:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|e4ebdc6180ee8876928d2e88fd658683ce83d8c3|1.69|2015-01-16 19:13:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|dac2c7c13787ce877ac865d910d7d33934f75a5c|1.69|2015-03-04 16:10:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|cad17db2008aa5a634b32948d894387c1b630dc2|1.69|2014-11-03 13:21:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|7c9a8d385726a7170d973e6166ff7657dda2e3d5|1.69|2015-03-09 16:12:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|03fdf69f5b33ebd53137f33b9e08998e20a62b4e|1.69|2014-10-18 10:06:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|3bbab34b7378e151072be223402e397fd1887517|1.69|2014-10-14 14:21:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|ad35c7ec930bcdf1647eb25499262efde4017b26|1.69|2014-12-30 12:19:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|a0a0f1ff49369934637c73563005888606f47aa8|1.69|2015-02-16 14:08:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|6dd6a2014a371f0cb3939709b8a4cfb242d48510|1.69|2014-11-09 13:10:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|f04b956d0647219a09b32346c74c625c8eb860bd|1.69|2015-02-23 11:52:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|6161fc3cbe7594b720f694060cfd83d19f2a2762|1.69|2014-10-07 12:00:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|43b7a198933593901ca80f11a9bd46e6aacbc654|1.69|2015-01-04 14:43:00|1.4094857484078087|4|1200000129|401|0.6146977543425921|0|26|55|-80.810056|8|35.219587|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|0.61471665291522548|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.810056|1.4104015459209989|401|1
35.219587|2fe323251f6d7c68f5784a36b3455bfd5b529736|5.98|2014-09-13 17:33:00|1.4094857484078087|4|5040073955|401|0.6146977543425921|0|26|1034|-80.810056|163|35.219587|HOT DOG|0.0|7|BALLPARK GLDN HOTDOG BUNS 12PK|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|0.61471665291522548|00050400739550|BUNS/ROLLS|COMMERCIAL BAKERY|-80.810056|1.4104015459209989|401|2
35.219587|40689b76d28bcbd0bc99570ff6a22660a573a995|1.69|2014-10-20 14:20:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|54|-80.826724|8|35.195689|DIET|0.0|23|CB DIET MT. DEW 20 OZ  SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001345|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|ba9be0e0297d35a403b786ce59d5826c360f7552|1.69|2014-11-06 12:53:00|80.810069425230125|4|1200000129|401|35.235071766875151|0|23|54|-80.826724|8|35.195689|DIET|0.0|23|CB DIET MT. DEW 20 OZ  SINGLES|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00012000001345|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.81006214331299|412|1
35.219587|83f98e42193cc768ccf4b8e6a5b5bd46385d8932|7.99|2014-12-23 17:12:00|80.810069425230125|4|3526600351|401|35.235071766875151|0|23|584|-80.826724|136|35.195689|TOPPINGS|1.0|4|CHOC PECAN OBSESSION|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00035266003519|OTHER MERCHANDISE|PRODUCE|-80.810056|80.81006214331299|412|1
35.219587|0adc30ed3cd4bd5eb0c9e598fc59f67cb8e824c0|0.99|2015-02-14 16:01:00|80.810069425230125|4|20506500000|401|35.235071766875151|0|23|2020|-80.826724|505|35.195689|CHEESE SPECIALTIES|0.0|6|SPECIALITY CHEESE BY COUNT|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00205065000006|SPECIALTY CHEESE|DELI|-80.810056|80.81006214331299|412|1
35.219587|1aa5da9a255b2798a2bfbf6326f6e333147a355c|1.0|2014-10-02 12:40:00|80.810069425230125|4|78352054321|401|35.235071766875151|0|23|8598|-80.826724|1792|35.195689|NEWSPAPERS|0.0|18|DAILY  CHARLOTTE OBSERVER|fcc73209ea573fa48b9f89d73e259a280697c041|1.0699600528872146|35.240679762029046|00783520543218|NEWSPAPERS|GM|-80.810056|80.81006214331299|412|1
35.06858|09308b33a37cfb977884eb0f2dc4bcfe92bf3b1a|4.99|2014-12-07 12:33:00|1.4091206135396188|1|7023430470|273|0.612062184999033|0|47|1220|-80.7007|275|35.06858|PASTA SC PREMIUM|2.5|1|GINA PASTA SC MARINARA|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00070234304151|PASTA SAUCES|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|6926f09ba12943495bc73940face9e5b12517b73|3.98|2014-10-25 19:54:00|1.4091206135396188|1|4800000095|273|0.612062184999033|0|47|190|-80.7007|29|35.06858|TUNA-CANNED|0.0|1|COS TUNA SOLID WHITE ALB|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00048000000958|SEAFOOD-CANNED|G1 GROCERY|-80.7007|1.4084929236641879|273|2
35.06858|355a2f586598f6dd52fbf2bccf4ddc209285bedf|5.29|2015-01-03 19:54:00|1.4091206135396188|1|4440018400|273|0.612062184999033|0|47|293|-80.7007|48|35.06858|FROZEN SEAFOOD|2.65|5|GORTON'S GRILLED TILAPIA|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00044400186506|FROZEN MEALS|FROZEN|-80.7007|1.4084929236641879|273|1
35.06858|8e8ea9e72701b94cfc04b0bb4b36bf997ebb61f5|1.49|2015-02-17 16:35:00|1.4091206135396188|1|2070901230|273|0.612062184999033|0|47|50|-80.7007|7|35.06858|PEG CANDY|0.0|1|TROLLI BRITE WATERMELON SHARKS|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00041420100826|CANDY|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|142d0eae4b751e18d93df8ba73647debbeda7aaf|5.98|2015-02-07 12:42:00|1.4091206135396188|1|7341013959|273|0.612062184999033|0|47|1031|-80.7007|162|35.06858|ITALIAN|2.0|7|ARNOLD ITALIAN BRD PP|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00073410139592|SLICED BREAD|COMMERCIAL BAKERY|-80.7007|1.4084929236641879|273|2
35.06858|dbc5545e9e60214b3ea87de43cd7b2cb4ee3f42e|3.55|2014-11-07 20:29:00|1.4091206135396188|1|7433610102|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HIGHLAND CREST 2% REDUCE FAT|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00074336101021|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|acac5a83114c1300e9005ea1afab8fdefe8569ac|3.75|2014-09-15 22:00:00|1.4091206135396188|1|7433610102|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HIGHLAND CREST 2% REDUCE FAT|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00074336101021|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|98a0e2b3edccec5082ef1caa22878de323d0e94b|2.99|2015-02-03 16:34:00|1.4091206135396188|1|7433610102|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HIGHLAND CREST 2% REDUCE FAT|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00074336101021|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|50090b9ec575ca621f68e03423bb76fadff098a8|2.99|2014-10-07 17:53:00|1.4091206135396188|1|7341013959|273|0.612062184999033|0|47|1031|-80.7007|162|35.06858|ITALIAN|0.5|7|ARNOLD ITALIAN BRD PP|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00073410139592|SLICED BREAD|COMMERCIAL BAKERY|-80.7007|1.4084929236641879|273|1
35.06858|1e51ab6044f1fa1e0094a7323acacbccf1ee9c95|5.98|2014-09-22 17:09:00|1.4091206135396188|1|7341013959|273|0.612062184999033|0|47|1031|-80.7007|162|35.06858|ITALIAN|1.49|7|ARNOLD ITALIAN BRD PP|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00073410139592|SLICED BREAD|COMMERCIAL BAKERY|-80.7007|1.4084929236641879|273|2
35.06858|83eff26e0d03ce7c9d1329433f43b7deca56b2c7|5.98|2015-02-13 17:21:00|1.4091206135396188|1|7433610102|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HIGHLAND CREST 2% REDUCE FAT|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00074336101021|MILK|DAIRY|-80.7007|1.4084929236641879|273|2
35.06858|6d2d55d8a70c99ed9791136684317b3873189503|2.99|2014-11-04 17:17:00|1.4091206135396188|1|7341013959|273|0.612062184999033|0|47|1031|-80.7007|162|35.06858|ITALIAN|0.5|7|ARNOLD ITALIAN BRD PP|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00073410139592|SLICED BREAD|COMMERCIAL BAKERY|-80.7007|1.4084929236641879|273|1
35.06858|74e7a822dd88ffb17c9517405b6b70335aec3348|3.49|2014-12-29 17:15:00|1.4091206135396188|1|7433610102|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HIGHLAND CREST 2% REDUCE FAT|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00074336101021|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|44e560294edf429c0d43c653c519ed57c195bab7|2.99|2015-03-05 17:30:00|1.4091206135396188|1|7433610102|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HIGHLAND CREST 2% REDUCE FAT|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00074336101021|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|3732c94e268c4f5a81bcd5c91eef8aed2ecfb3c3|5.79|2014-11-23 07:59:00|80.700712769248256|1|7247000603|273|35.077874295458152|0|42|1641|-80.699686|377|35.000049|PACKAGED DONUTS|0.0|14|K K 12 CT GLAZED DONUTS PP|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|35.088667338853092|00072470006035|DONUTS|BAKERY|-80.7007|80.700708062916888|249|1
35.06858|fd7f78782586dcf178475fe4cfffaacd0bec923a|5.98|2015-02-17 14:00:00|1.4091206135396188|1|7433610102|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HIGHLAND CREST 2% REDUCE FAT|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00074336101021|MILK|DAIRY|-80.7007|1.4084929236641879|273|2
35.06858|a3ddfb3bf8be9c011774af53734ef345d44a5e1f|2.99|2014-09-17 17:40:00|1.4091206135396188|1|7341013959|273|0.612062184999033|0|47|1031|-80.7007|162|35.06858|ITALIAN|1.5|7|ARNOLD ITALIAN BRD PP|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00073410139592|SLICED BREAD|COMMERCIAL BAKERY|-80.7007|1.4084929236641879|273|1
35.06858|ceda73b9faba66d43e6a1bf242d122acb0962fa7|5.98|2015-02-23 17:36:00|1.4091206135396188|1|7433610102|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HIGHLAND CREST 2% REDUCE FAT|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00074336101021|MILK|DAIRY|-80.7007|1.4084929236641879|273|2
35.06858|3f24ca0d9b25ce32563f2d8348ab9a5b3c435250|3.75|2014-09-21 16:29:00|1.4091206135396188|1|7433610102|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HIGHLAND CREST 2% REDUCE FAT|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00074336101021|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|7b2bb3e5ec839692af4e4ed32be649f904361d98|2.99|2014-10-10 17:41:00|1.4091206135396188|1|7341013959|273|0.612062184999033|0|47|1031|-80.7007|162|35.06858|ITALIAN|0.5|7|ARNOLD ITALIAN BRD PP|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00073410139592|SLICED BREAD|COMMERCIAL BAKERY|-80.7007|1.4084929236641879|273|1
35.06858|701d98ae74ea1c6e22056bbd654b247716257e7b|9.99|2014-12-23 20:53:00|1.4091206135396188|1|7203661033|273|0.612062184999033|0|47|666|-80.7007|145|35.06858|PACKAGED COOKED|2.0|12|HT COOKED SHRIMP RING 10OZ|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036610331|SHRIMP|SEAFOOD|-80.7007|1.4084929236641879|273|1
35.06858|181baa3a29d064e85a7df99c9c09b4ebd21daf49|3.0|2014-09-14 19:47:00|1.4091206135396188|1|7203655029|273|0.612062184999033|0|47|331|-80.7007|52|35.06858|NATURAL SLICED|1.0|3|HT MOZZARELLA SLICES|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036550293|CHEESE|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|e20f029eb8e2de8f0d234e34639193158b171a41|12.99|2014-09-27 13:47:00|1.4091206135396188|1|7203695587|273|0.612062184999033|0|47|1707|-80.7007|387|35.06858|MESSAGE|3.0|14|12 INCH MESSAGE COOKIE|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036955876|COOKIES|BAKERY|-80.7007|1.4084929236641879|273|1
35.06858|c6361d7dfaf9f5a143d77e43a58ec6e7160f45e5|1.79|2015-03-08 12:55:00|1.4091206135396188|1||273|0.612062184999033|0|47|535|-80.7007|64|35.06858|FRESH GREENS|0.0|4|SPINACH, BUNCH (RPC)|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00204090000005|FRESH PRODUCE|PRODUCE|-80.7007|1.4084929236641879|273|1
35.06858|56cf7562542293450686e61637ddd99640607908|1.99|2015-01-12 21:23:00|1.4091206135396188|1|74236500454|273|0.612062184999033|0|47|1441|-80.7007|274|35.06858|MAC AND CHEESE|0.74|1|HORIZON CLASSIC MAC AND CHEESE|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00742365004544|PREP FOODS DINNERS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|b6cdf12e7aab148a35cd4b64c7b7ef846094b4d9|3.98|2014-11-09 13:22:00|1.4091206135396188|1|74236500454|273|0.612062184999033|0|47|1441|-80.7007|274|35.06858|MAC AND CHEESE|1.98|1|HORIZON CLASSIC MAC AND CHEESE|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00742365004544|PREP FOODS DINNERS|G1 GROCERY|-80.7007|1.4084929236641879|273|2
35.06858|e437bb8bb82bb5cb13fc8bc139f07462324e964d|6.99|2014-10-20 17:40:00|1.4091206135396188|1|68243020025|273|0.612062184999033|0|47|31|-80.7007|4|35.06858|NON CARBONATED WATER|0.0|1|VOSS WATER PET 6PK|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00682430200252|BOTTLED WATER|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|43844aa6b1a19c063680367697eb716bd9708506|11.98|2014-12-13 14:37:00|80.700712769248256|1|4116740002|273|35.077874297799774|0|42|4436|-80.64817|1210|35.04711|DIARRHEA REMEDY-LIQUID|0.0|17|KAOPECTATE REGULAR 40002|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|35.088667338853092|00041167400029|STOMACH REMEDIES|HBC|-80.7007|80.700700160737696|129|2
35.06858|fe0c8700d55650672f58ffbd5feae3b61c130480|5.99|2014-11-16 14:58:00|1.4091206135396188|1|4116740002|273|0.612062184999033|0|47|4436|-80.7007|1210|35.06858|DIARRHEA REMEDY-LIQUID|0.0|17|KAOPECTATE REGULAR 40002|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00041167400029|STOMACH REMEDIES|HBC|-80.7007|1.4084929236641879|273|1
35.06858|c934d5d2b1c9b8bbd7feb84b6c08355de6528192|4.49|2014-12-24 13:25:00|1.4091206135396188|1|4180071500|273|0.612062184999033|0|47|131|-80.7007|20|35.06858|GRAPE JUICE-SHELF|2.25|1|WELCH'S SPARKLING WHITE GRAPE|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00041800715008|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|c04bf656405ec6d585345cf75708f1e5e6c1e7ad|1.39|2014-10-04 16:51:00|1.4091206135396188|1|3710003578|273|0.612062184999033|0|47|245|-80.7007|39|35.06858|VEGETABLES-CORE|0.39|1|LIBBY WK CORN|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00037100036622|VEGETABLES-CAN/JAR|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|a675f8a820bfaf1e11faa283e955bdb5255c5650|3.55|2015-01-18 17:52:00|1.4091206135396188|1|3620001401|273|0.612062184999033|0|47|1221|-80.7007|275|35.06858|PASTA SC VALUE|1.05|1|RAGU SC 45 OWS TRADITIONAL|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00036200014011|PASTA SAUCES|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|faea833e8a785097338bb0f62faff700a5a1c804|0.99|2014-10-19 21:26:00|1.4091206135396188|1|5210009860|273|0.612062184999033|0|47|75|-80.7007|34|35.06858|GRAVY MIXES|0.0|1|E  MC BROWN GRAVY MIX|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00052100098609|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|68dcaf60b7e2ddcc32419d1dc8e4af2363ebc3fa|1.27|2014-11-01 17:59:00|1.4091206135396188|1|7203624010|273|0.612062184999033|0|47|150|-80.7007|23|35.06858|NOODLES/DUMPLINGS-DRY|0.0|1|HT NOODLE EGG WIDE|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036240101|PASTA|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|e0c130039e4520b6bdddb5ace224d275bd210a79|1.67|2015-02-16 17:09:00|1.4091206135396188|1|7203613031|273|0.612062184999033|0|47|716|-80.7007|15|35.06858|SELF-RISING|0.0|1|HARRIS TEETER S/RISING FLOUR|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036130310|FLOUR|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|95ee8078fc4db41edf6bb215c0a2877c31aae177|0.67|2014-11-12 16:23:00|80.700712769248256|1|7203629030|273|35.077874297799774|0|42|179|-80.64817|27|35.04711|CANNED PASTA|0.0|1|HT SPAGHETTI RINGS|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|35.088667338853092|00072036290359|PREPARED FOODS-RTS|G1 GROCERY|-80.7007|80.700700160737696|129|1
35.06858|854dca6c20a6265ecdaab59e18688e8e8bd7f9bd|3.99|2015-01-15 16:57:00|1.4091206135396188|1|7835470843|273|0.612062184999033|0|47|317|-80.7007|52|35.06858|CHUNK AND BAR CHEESE|1.49|3|CABOT MONTEREY JACK|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00078354702185|CHEESE|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|6b71cd3b6db48fb67118adf823d15fff332edf9a|2.99|2015-02-07 15:47:00|1.4091206135396188|1|7203670381|273|0.612062184999033|0|47|5558|-80.7007|1508|35.06858|LAUNDRY SUPPLIES|1.0|18|(JHK)(PPL) YH W/M SPR BTL 24OZ|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036703811|LAUNDRY/IRONING/VACUUM|GM|-80.7007|1.4084929236641879|273|1
35.06858|a95cd3b7541c38282c3d1454f708020cd867f73c|2.59|2014-12-19 10:42:00|1.4091206135396188|1|7203670440|273|0.612062184999033|0|47|729|-80.7007|69|35.06858|NFS-SCOUR PAD/STEEL WOOL|0.0|1|YH HVY DUTY SCOURING PADS 3CT|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036704405|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|84bc99f91d8ac6fee9a7c98714b85cf591510d3c|2.39|2014-10-17 17:39:00|80.700712769248256|1|7203670014|273|35.077874297800669|0|42|4816|-80.732725|1235|35.082768|FIRST AID ADHESIVE BANDG|0.89|17|HT PLASTIC STRIP BANDAGE-70014|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|35.088667338853092|00072036700148|FIRST AID|HBC|-80.7007|80.700700032126576|147|1
35.06858|80f4b129444351dd06a4125f6c2bcf19575065bb|2.99|2014-12-22 13:06:00|1.4091206135396188|1|7203620074|273|0.612062184999033|0|47|128|-80.7007|20|35.06858|APPLE JUICE-SHELF|0.99|1|HT APPLE JUICE NATURAL|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036200747|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|937df9f7b6a9e9fe0daf8178a340f5b8abe40cff|2.79|2015-02-21 17:29:00|1.4091206135396188|1|7203698295|273|0.612062184999033|0|47|81|-80.7007|9|35.06858|RTE CEREAL KIDS|0.32|1|HT CER COCOA PEANUT BUTTER|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036170101|CEREAL|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|f3e63af40b9b29730e4143699c3499e4315f7908|1.39|2015-02-25 18:22:00|1.4091206135396188|1|7203608016|273|0.612062184999033|0|47|70|-80.7007|11|35.06858|KETCHUP|0.39|1|HT KETCHUP 24|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036080165|CONDIMENTS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|a5c5a09588d069d4c2d31be5f6f5d537f986102a|2.49|2015-03-08 16:00:00|1.4091206135396188|1|7203609056|273|0.612062184999033|0|47|1253|-80.7007|12|35.06858|ALL OTHER COOKIES|0.0|1|HT VANILLA WAFERS|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036090560|COOKIES|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|5998b3d7a3e29a08b5980aa43958a067aecca1b3|1.39|2014-12-31 13:59:00|1.4091206135396188|1|7203602056|273|0.612062184999033|0|47|78|-80.7007|11|35.06858|MUSTARD|0.7|1|HT MUSTARD YELLOW 14 OZ|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036020567|CONDIMENTS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|e1b4e264fcc92ec0de5223c6885317bc9dbf6ee6|2.79|2014-09-29 20:52:00|1.4091206135396188|1|7203698295|273|0.612062184999033|0|47|81|-80.7007|9|35.06858|RTE CEREAL KIDS|1.29|1|HT CER COCOA PEANUT BUTTER|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036170101|CEREAL|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|690543a19610af258b2114b1b8f0380cae37a445|1.54|2015-02-05 17:52:00|1.4091206135396188|1|7203632360|273|0.612062184999033|0|47|1441|-80.7007|274|35.06858|MAC AND CHEESE|0.0|1|HT DIN MAC CHEESE|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036323606|PREP FOODS DINNERS|G1 GROCERY|-80.7007|1.4084929236641879|273|2
35.06858|91081f21a9abe0265cca1a6b2762283498071772|4.29|2015-01-23 22:02:00|1.4091206135396188|1|2840015938|273|0.612062184999033|0|47|201|-80.7007|31|35.06858|POTATO CHIPS|1.79|1|RUFFLES ULTIMATE BCN CHED SKIN|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00028400208949|SNACKS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|80bdfe2d9b62972d9e75b6abc8025fe3d13c5c6a|3.29|2014-10-21 18:11:00|1.4091206135396188|1|2840011895|273|0.612062184999033|0|47|204|-80.7007|31|35.06858|TORTILLA CHIPS|0.79|1|TOSTITOS CANTINA TRADITIONAL|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00028400118958|SNACKS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|1d00de98f1b5d075285117a0a2555eed8e22efbe|2.19|2015-02-27 21:50:00|1.4091206135396188|1|7225003106|273|0.612062184999033|0|47|1031|-80.7007|162|35.06858|ITALIAN|0.69|7|SPOLETTO ITALIAN BREAD|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072250031066|SLICED BREAD|COMMERCIAL BAKERY|-80.7007|1.4084929236641879|273|1
35.06858|4185235950eb13b124b511a58ff2a7e743d19b02|2.39|2014-12-24 14:14:00|1.4091206135396188|1|7203695175|273|0.612062184999033|0|47|1607|-80.7007|371|35.06858|FROZEN DOUGH (BREAD)|0.0|14|FRESH LRG FRENCH BREAD|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036951755|BREAD|BAKERY|-80.7007|1.4084929236641879|273|1
35.06858|5e07f56d40d2ed750986b0de12627f1743acc019|3.49|2014-12-04 16:53:00|1.4091206135396188|1|2840023981|273|0.612062184999033|0|47|203|-80.7007|31|35.06858|CHEESE SNACKS|0.0|1|CHEETOS JUMBO PUFFS|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00028400239875|SNACKS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|4d4a4ad2af8de8f6dc2c57f61e90ceab607cb174|2.89|2014-09-26 17:34:00|1.4091206135396188|1|2100065894|273|0.612062184999033|0|47|1441|-80.7007|274|35.06858|MAC AND CHEESE|0.0|1|KRAFT DIN MAC CHS FAMILY|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00021000658947|PREP FOODS DINNERS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|eaa33ce8e0c28b031f0482799215ba5c2cccb802|3.33|2015-01-05 20:31:00|1.4091206135396188|1|7203643010|273|0.612062184999033|0|47|252|-80.7007|45|35.06858|PREMIUM ICE CREAM|0.0|5|HT SMTH & CRMY COOKIE DOUGH IC|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036981714|ICE CREAM|FROZEN|-80.7007|1.4084929236641879|273|1
35.06858|aa18935ae737541a1605507fcb53ddfea4b72296|0.97|2014-11-18 21:04:00|1.4091206135396188|1|7203671102|273|0.612062184999033|0|47|1025|-80.7007|162|35.06858|WHITE|0.0|7|HT OLD FASHIONED BREAD|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036711021|SLICED BREAD|COMMERCIAL BAKERY|-80.7007|1.4084929236641879|273|1
35.06858|7f7d0538cad96601f7c43499695e4f0f092d0ae9|0.97|2014-10-30 19:00:00|1.4091206135396188|1|7203671102|273|0.612062184999033|0|47|1025|-80.7007|162|35.06858|WHITE|0.0|7|HT OLD FASHIONED BREAD|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036711021|SLICED BREAD|COMMERCIAL BAKERY|-80.7007|1.4084929236641879|273|1
35.06858|c8ee2635a03dad481dd3911a8ebd3dd9144fb3fa|1.17|2014-11-29 17:11:00|1.4091206135396188|1|7203690021|273|0.612062184999033|0|47|1033|-80.7007|163|35.06858|HAMBURGER|0.0|7|H T HAMBURGER BUNS|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036900210|BUNS/ROLLS|COMMERCIAL BAKERY|-80.7007|1.4084929236641879|273|1
35.06858|bd77fbbda2511b3ea79a58c8805f3b31800f4a2c|0.97|2014-09-16 18:46:00|1.4091206135396188|1|7203671102|273|0.612062184999033|0|47|1025|-80.7007|162|35.06858|WHITE|0.0|7|HT OLD FASHIONED BREAD|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036711021|SLICED BREAD|COMMERCIAL BAKERY|-80.7007|1.4084929236641879|273|1
35.06858|f1710c21c2dd53b3817427d95872136cc11c8f45|1.37|2015-02-08 12:42:00|80.700712769248256|1|7203690021|273|35.077874295458152|0|42|1033|-80.699686|163|35.000049|HAMBURGER|0.0|7|H T HAMBURGER BUNS|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|35.088667338853092|00072036900210|BUNS/ROLLS|COMMERCIAL BAKERY|-80.7007|80.700708062916888|249|1
35.06858|92f38916a59fe013fdf7519a556c1a2f8f8b98e4|0.97|2015-01-02 16:46:00|1.4091206135396188|1|7203671102|273|0.612062184999033|0|47|1025|-80.7007|162|35.06858|WHITE|0.0|7|HT OLD FASHIONED BREAD|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036711021|SLICED BREAD|COMMERCIAL BAKERY|-80.7007|1.4084929236641879|273|1
35.06858|507deb2b1e6ab8fb06c18c38d721273b50524f70|2.89|2014-12-09 18:17:00|1.4091206135396188|1|7203695922|273|0.612062184999033|0|47|1625|-80.7007|373|35.06858|FROZEN DOUGH (ROLLS)|0.0|14|FRESH WHITE SUB ROLLS 4 CT.|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036959225|ROLLS|BAKERY|-80.7007|1.4084929236641879|273|1
35.06858|87e77d6b6f7500d956dbe2ee6564159a6ee0b817|2.29|2014-11-14 17:39:00|1.4091206135396188|1|7800023046|273|0.612062184999033|0|47|55|-80.7007|8|35.06858|REGULAR|1.29|23|CHEERWINE 2 LTR NR|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00070925000300|CARBONATED BEVERAGES|BEVERAGE|-80.7007|1.4084929236641879|273|1
35.06858|d088923fe7300dec1c74cdf1830cbdad28e15d71|2.29|2014-09-12 17:47:00|80.700712769248256|1|7800023046|273|35.077874297799774|0|42|55|-80.64817|8|35.04711|REGULAR|0.79|23|CHEERWINE 2 LTR NR|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|35.088667338853092|00070925000300|CARBONATED BEVERAGES|BEVERAGE|-80.7007|80.700700160737696|129|1
35.06858|042befa8c3b9c55945aae725863b9f8a430b38a0|7.99|2014-10-11 18:00:00|1.4091206135396188|1|7203629093|273|0.612062184999033|0|47|152|-80.7007|24|35.06858|NFS-CAT FOOD DRY|0.0|1|HT YOURPET ADULT CAT FOOD|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036290939|PET FOOD/SUPPLIES|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|e54b912b1131dc6189d043519803a77912732f12|1.29|2015-01-17 13:12:00|1.4091206135396188|1|5100002524|273|0.612062184999033|0|47|179|-80.7007|27|35.06858|CANNED PASTA|0.29|1|SPAGHETTIOS ORIGINAL|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00051000025241|PREPARED FOODS-RTS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|14cb5f7f2494e933b7d37aab2f0aaece87c098be|1.99|2014-11-08 07:42:00|1.4091206135396188|1|5100017520|273|0.612062184999033|0|47|1201|-80.7007|33|35.06858|RTS CANNED|0.49|1|CAM HOMESTYLE HR CHIC BRN RICE|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00051000169044|SOUP|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|f8302e9e1258619805d8eb5928b6292e050c118b|1.29|2014-12-11 17:03:00|1.4091206135396188|1|5100002524|273|0.612062184999033|0|47|179|-80.7007|27|35.06858|CANNED PASTA|0.29|1|SPAGHETTIOS CHEESY PIZZA|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00051000213990|PREPARED FOODS-RTS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|67f7f06224ec7cc7db2021400c52c5045833244d|0.79|2014-12-27 21:51:00|1.4091206135396188|1|7294075709|273|0.612062184999033|0|47|257|-80.7007|39|35.06858|TOMATOES|0.12|1|TUTTOROSSO TOMATO PASTE 6 OZ.|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072940757092|VEGETABLES-CAN/JAR|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|1fd829dcce02906ec509f2362a242739f8996700|9.98|2015-01-24 15:55:00|1.4091206135396188|1|8265750406|273|0.612062184999033|0|47|31|-80.7007|4|35.06858|NON CARBONATED WATER|2.98|1|(U)DEER PARK WATER 24PK .5LT|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00082657504063|BOTTLED WATER|G1 GROCERY|-80.7007|1.4084929236641879|273|2
35.06858|2e5701412e57b005132c0c28d2aefd78e75246fc|0.99|2014-09-12 17:46:00|80.700712769248256|1|7780200651|273|35.077874297799774|0|42|3055|-80.64817|1000|35.04711|BRAND-WET N WILD|0.0|17|C655 WET WILD CHARCOAL EYELINE|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|35.088667338853092|00077802006554|COSMETICS|HBC|-80.7007|80.700700160737696|129|1
35.06858|1fb7bedee3a54865d29dfcde432d77df78e9f788|0.59|2015-01-26 17:23:00|1.4091206135396188|1|7978454482|273|0.612062184999033|0|47|6524|-80.7007|1564|35.06858|ACTIVITY PAPER|0.0|18|POSTER BOARD WHITE 4 PLY 22X28|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00079784544826|SCHOOL & OFFICE SUPPLY|GM|-80.7007|1.4084929236641879|273|1
35.06858|ca8b5ebab08aed295f6e141190edfe30c08bf4b1|5.49|2014-12-05 13:48:00|80.700712769248256|1|827411111|273|35.077874297799774|0|42|55|-80.64817|8|35.04711|REGULAR|1.5|23|VIRGILS CREAM SODA|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|35.088667338853092|00090341543212|CARBONATED BEVERAGES|BEVERAGE|-80.7007|80.700700160737696|129|1
35.06858|f3f4d67765a291a4011840d736a160ca2e5aabf1|1.34|2014-10-01 18:02:00|1.4091206135396188|1|3100010101|273|0.612062184999033|0|47|1279|-80.7007|48|35.06858|SINGLE SERVE FLAVOR|0.0|5|BANQUET BEEF POT PIE|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00031000101022|FROZEN MEALS|FROZEN|-80.7007|1.4084929236641879|273|2
35.06858|74d9ec87c6c57e35bdb2f7f762678ae7524d0f41|0.67|2015-03-09 17:09:00|1.4091206135396188|1|3100010101|273|0.612062184999033|0|47|1279|-80.7007|48|35.06858|SINGLE SERVE FLAVOR|0.0|5|BANQUET BEEF POT PIE|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00031000101022|FROZEN MEALS|FROZEN|-80.7007|1.4084929236641879|273|1
35.06858|28a6d8ad8cf5a96da981c669b671aabb35037fb3|6.98|2014-12-28 13:00:00|1.4091206135396188|1|2840024053|273|0.612062184999033|0|47|198|-80.7007|31|35.06858|CORN CHIPS|0.0|1|FRITOS REGULAR|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00028400240536|SNACKS|G1 GROCERY|-80.7007|1.4084929236641879|273|2
35.06858|1985996edea4854659eb53341c5511bed63caade|4.99|2015-01-31 16:01:00|1.4091206135396188|1|2840015297|273|0.612062184999033|0|47|204|-80.7007|31|35.06858|TORTILLA CHIPS|1.0|1|DORITOS NACHO CHEES PARTY SIZE|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00028400152976|SNACKS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|6d5738c18247e96d05755a9944e665bbfbd43be2|0.74|2015-01-09 07:57:00|1.4091206135396188|1||273|0.612062184999033|0|47|500|-80.7007|64|35.06858|FRESH APPLES|0.0|4|RED DEL APPLE, WA  48|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00233284000002|FRESH PRODUCE|PRODUCE|-80.7007|1.4084929236641879|273|1
35.06858|f1ace35c2b071aeacef19530160652a184df77d1|3.99|2015-01-25 16:09:00|1.4091206135396188|1|7910090202|273|0.612062184999033|0|47|155|-80.7007|24|35.06858|NFS-DOG TREATS|0.71|1|MILK-BONE DOG BSCUTS-MEDIUM|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00079100514106|PET FOOD/SUPPLIES|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|0751ac56d87c1840336d57fa166133ecc320baf3|1.89|2014-11-03 19:13:00|1.4091206135396188|1|1200062036|273|0.612062184999033|0|47|1214|-80.7007|272|35.06858|AUTHENTIC HISPANIC|0.0|1|PEPSI-MEXICAN|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00012000620362|HISPANIC PREP. FOODS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|b9ba7eb4ae476ab60ad59b1fea59b11eb5a7079c|2.69|2014-12-02 19:43:00|80.700712769248256|1|7102501597|273|35.077874295458152|0|42|1025|-80.699686|162|35.000049|WHITE|0.7|7|BUNNY OLD FASHIONED BREAD|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|35.088667338853092|00071025015973|SLICED BREAD|COMMERCIAL BAKERY|-80.7007|80.700708062916888|249|1
35.06858|d0107ad40bae3ec739f837d4eb522c6400110fd6|2.19|2014-11-09 17:22:00|1.4091206135396188|1|1200000496|273|0.612062184999033|0|47|54|-80.7007|8|35.06858|DIET|0.69|23|DIET WILD CHERRY PEPSI 2 LITER|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00012000003417|CARBONATED BEVERAGES|BEVERAGE|-80.7007|1.4084929236641879|273|1
35.06858|e5de0f06a7ad5c0ca3be0dbaa4a664db518193f9|3.79|2014-12-20 14:01:00|1.4091206135396188|1|7910051352|273|0.612062184999033|0|47|155|-80.7007|24|35.06858|NFS-DOG TREATS|0.0|1|MILK BONE DOG BISCUITS MEDIUM|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00079100513529|PET FOOD/SUPPLIES|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|e1cec71b1aac83508815d1810b703991764c22dd|2.99|2015-01-08 18:00:00|1.4091206135396188|1|7433610102|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HIGHLAND CREST WHOLE MILK|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00074336879203|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|9e2af1df14ca8546e7be1bdf7a299839374696da|6.99|2014-11-10 12:49:00|80.700712769248256|1|7468210906|273|35.077874297799774|0|42|128|-80.64817|20|35.04711|APPLE JUICE-SHELF|1.0|1|I/O KNUDSEN CIDER 96 OZ|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|35.088667338853092|00074682109061|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.7007|80.700700160737696|129|1
35.06858|a27fddf90eebecd78c77ad11b08d2a6567bc3886|2.49|2015-01-11 21:30:00|1.4091206135396188|1|4369505631|273|0.612062184999033|0|47|1276|-80.7007|279|35.06858|FROZEN SANDWICHES|0.49|5|HOT PKT CHICKEN MELT|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00043695071085|FROZEN SANDWICH AND SNACKS|FROZEN|-80.7007|1.4084929236641879|273|1
35.06858|9f61f68c28d53d61842ba005e8938aef16a6eb44|8.79|2015-01-25 17:42:00|1.4091206135396188|1|4133382501|273|0.612062184999033|0|47|8433|-80.7007|1769|35.06858|ALKALINE AA|0.0|18|(JHK) (FE) DU CPPRTOP  AA 8PK|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00041333825014|BATTERY & FLASHLIGHT|GM|-80.7007|1.4084929236641879|273|1
35.06858|4bb8867ac43849042089948c047d606d6aec9e50|1.0|2015-01-12 17:18:00|1.4091206135396188|1|4000000435|273|0.612062184999033|0|47|47|-80.7007|7|35.06858|REGISTER BARS|0.0|1|(FE)3-MUSKETEER BARS|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00040000422082|CANDY|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|c56f67039bbb52417b64fd3a2ef3a2cc1121f850|3.19|2014-11-22 12:02:00|1.4091206135396188|1|3900008568|273|0.612062184999033|0|47|175|-80.7007|27|35.06858|CANNED MEATS|0.0|1|LIBBYS CORNED BEEF HASH|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00039000085687|PREPARED FOODS-RTS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|1c8aa005f50ccc9a48e8afa4f22c38859f1bd264|10.5|2015-01-02 21:25:00|1.4091206135396188|1|7203698425|273|0.612062184999033|0|47|254|-80.7007|892|35.06858|PREMIUM PIZZA|1.5|5|HT THIN CRUST PEPP/SAUS PIZZA|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036984265|FROZEN PIZZA|FROZEN|-80.7007|1.4084929236641879|273|3
35.06858|10b53ea62fa1152b17ef1e629efce35ae11e936f|8.78|2014-12-05 17:02:00|1.4091206135396188|1|4400002747|273|0.612062184999033|0|47|91|-80.7007|13|35.06858|SPRAYED BUTTER CRACKERS|0.91|1|RITZ REDUCED FAT|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00044000031183|CRACKERS|G1 GROCERY|-80.7007|1.4084929236641879|273|2
35.06858|bcc6289a060595005c499dbd09a1619de4b8f17e|2.79|2015-02-20 21:45:00|1.4091206135396188|1|4227200070|273|0.612062184999033|0|47|1277|-80.7007|279|35.06858|FROZEN SNACKS|0.0|5|AMY'S BEAN & RICE BURRITO N-D|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00042272000708|FROZEN SANDWICH AND SNACKS|FROZEN|-80.7007|1.4084929236641879|273|1
35.06858|bfbb83e3a5aa78a012fa4ec83623cae7a34721f7|3.39|2014-09-20 07:17:00|1.4091206135396188|1|7203698705|273|0.612062184999033|0|47|4317|-80.7007|1205|35.06858|IBUPROFEN|1.42|17|HT IBUPROFEN TABLETS BROWN|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036987051|PAIN RELIEF|HBC|-80.7007|1.4084929236641879|273|1
35.06858|f2245e08cd4a63b00d3517eb029bf81039423c31|2.99|2015-01-21 16:12:00|1.4091206135396188|1|3700000309|273|0.612062184999033|0|47|4072|-80.7007|1080|35.06858|TOOTHPASTE-CAVITY|0.49|17|CREST REG ANTCAVITY TPASTE GEL|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00037000003120|ORAL HYGIENE|HBC|-80.7007|1.4084929236641879|273|1
35.06858|298b5694683ec17bfcdeb10a67e296d26c704e6c|0.87|2014-10-31 07:33:00|80.700712769248256|1|7203610114|273|35.077874297799774|0|42|55|-80.64817|8|35.04711|REGULAR|0.0|23|HT ROOT BEER 2 LITER|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|35.088667338853092|00072036110251|CARBONATED BEVERAGES|BEVERAGE|-80.7007|80.700700160737696|129|1
35.06858|c61845b0fc2bd42314e20eb765716db1260289c6|0.87|2015-02-11 17:16:00|1.4091206135396188|1|7203610114|273|0.612062184999033|0|47|55|-80.7007|8|35.06858|REGULAR|0.0|23|HT COLA 2 LITER|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036101143|CARBONATED BEVERAGES|BEVERAGE|-80.7007|1.4084929236641879|273|1
35.06858|bb4aac9aba2b8968bf41acd084887da0227250dd|6.58|2014-11-21 16:07:00|1.4091206135396188|1|1600027527|273|0.612062184999033|0|47|74|-80.7007|9|35.06858|RTE CEREAL ALL FAMILY|1.58|1|GM CHEERIOS HONEY NUT 12.25OZ|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00016000275270|CEREAL|G1 GROCERY|-80.7007|1.4084929236641879|273|2
35.06858|3fb4eda0383936211721dfc2a9ab2a0fb182f768|6.98|2015-02-20 17:42:00|1.4091206135396188|1|3760011544|273|0.612062184999033|0|47|175|-80.7007|27|35.06858|CANNED MEATS|0.0|1|SPAM 12 OZ|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00037600138727|PREPARED FOODS-RTS|G1 GROCERY|-80.7007|1.4084929236641879|273|2
35.06858|57fee180827471449245b22c9cf2293fd37ed8b5|1.39|2015-02-20 21:42:00|1.4091206135396188|1|4100002253|273|0.612062184999033|0|47|1439|-80.7007|274|35.06858|DRY DINNERS|0.0|1|KNORR PASTA PARMESAN|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00041000022555|PREP FOODS DINNERS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|ef52cf859217faf05540b13eec7493aef98d0687|7.9|2014-12-14 15:31:00|1.4091206135396188|1|7203663995|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|1.98|3|HARRIS TEETER 2% MILK|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036639981|MILK|DAIRY|-80.7007|1.4084929236641879|273|2
35.06858|7aa5faa9d688d28bc2dcd345015222a33dec072d|0.99|2014-09-10 13:50:00|80.700712769248256|1|7203695306|273|35.077874297799774|0|42|1895|-80.64817|450|35.04711|TEA|0.0|6|FFM SWEET TEA|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|35.088667338853092|00072036953063|BEVERAGES|DELI|-80.7007|80.700700160737696|129|1
35.06858|f550ef45eaea6b7e68351b36a875c1614b7c207a|0.99|2014-10-29 17:24:00|1.4091206135396188|1|1708289774|273|0.612062184999033|0|47|206|-80.7007|31|35.06858|FRONT END SNACKS|0.0|1|J LINKS CLSC BEEF STKS PP $.99|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00017082897749|SNACKS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|d6b7602df81dac7d136f6f34be848857525f1ed9|0.99|2014-10-11 14:16:00|1.4091206135396188|1|1708289774|273|0.612062184999033|0|47|206|-80.7007|31|35.06858|FRONT END SNACKS|0.0|1|J LINKS CLSC BEEF STKS PP $.99|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00017082897749|SNACKS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|1b638bf62dbb7655fd6114228e3efb37e557c502|5.49|2015-01-23 14:24:00|1.4091206135396188|1|827411111|273|0.612062184999033|0|47|55|-80.7007|8|35.06858|REGULAR|0.0|23|VIRGILS BLACK CHERRY CREAM|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00090341231157|CARBONATED BEVERAGES|BEVERAGE|-80.7007|1.4084929236641879|273|1
35.06858|f3e1c93869c6c5919928c5c64452965429baa0c1|1.89|2014-09-15 17:28:00|1.4091206135396188|1|3400000220|273|0.612062184999033|0|47|47|-80.7007|7|35.06858|REGISTER BARS|0.0|1|REESE'S PB CUP KING|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00034000004805|CANDY|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|76b116dbe329a56aebf1b9ea435832832a049fce|4.58|2014-12-17 19:08:00|1.4091206135396188|1|1900008501|273|0.612062184999033|0|47|50|-80.7007|7|35.06858|PEG CANDY|0.0|1|LIFESAVERS FIVE FLAVOR BAG|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00019000085016|CANDY|G1 GROCERY|-80.7007|1.4084929236641879|273|2
35.06858|81a8d3722359d1f9ba40f98a43e90b019a48885b|2.69|2014-11-05 21:34:00|1.4091206135396188|1|7373100415|273|0.612062184999033|0|47|495|-80.7007|108|35.06858|NON REFRIGERATED|0.19|19|MISSION SOFT TACO 10 CT|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00073731004159|TORTILLAS|CASE READY MEATS|-80.7007|1.4084929236641879|273|1
35.06858|f4cc0818a31ffed7aee27b5fe8d4967596085c85|4.39|2014-10-14 21:44:00|1.4091206135396188|1|7433610006|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HUNTER 2%  MILK GALLON|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00074336100222|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|f04528d4c9ed0c4b5f7f09990cea2a7e75959464|1.69|2014-10-30 19:01:00|1.4091206135396188|1|1200000129|273|0.612062184999033|0|47|55|-80.7007|8|35.06858|REGULAR|0.0|23|CB DR PEPPER 20 OZ NR SINGLE|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00078000082401|CARBONATED BEVERAGES|BEVERAGE|-80.7007|1.4084929236641879|273|1
35.06858|4a80b53c89db076583856d09a2d2c8c3d1063e87|1.69|2015-01-30 17:25:00|1.4091206135396188|1|1200000129|273|0.612062184999033|0|47|55|-80.7007|8|35.06858|REGULAR|0.0|23|CB DR PEPPER 20 OZ NR SINGLE|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00078000082401|CARBONATED BEVERAGES|BEVERAGE|-80.7007|1.4084929236641879|273|1
35.06858|95883f56fa12dc73298ee7995b5490670258aa82|2.19|2015-01-06 18:31:00|1.4091206135396188|1|7800008246|273|0.612062184999033|0|47|54|-80.7007|8|35.06858|DIET|0.2|23|DIET DR PEPPER 2 LITER|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00078000083460|CARBONATED BEVERAGES|BEVERAGE|-80.7007|1.4084929236641879|273|1
35.06858|a7d008cccb3343dce90cd090b331c30878da8b83|2.19|2014-11-30 20:06:00|1.4091206135396188|1|1200000496|273|0.612062184999033|0|47|54|-80.7007|8|35.06858|DIET|0.69|23|DIET PEPSI 2 LTR NR|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00012000002311|CARBONATED BEVERAGES|BEVERAGE|-80.7007|1.4084929236641879|273|1
35.06858|62379bc7272b2f8914e011b7c931f08406d8997a|3.39|2014-12-05 08:25:00|1.4091206135396188|1|1312000286|273|0.612062184999033|0|47|1471|-80.7007|278|35.06858|HASH BROWN POTATOES|0.5|5|ORE-IDA SOUTH STYLE HASH BRWN|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00013120003929|FROZEN POTATO|FROZEN|-80.7007|1.4084929236641879|273|1
35.06858|2e8766be3d41738d812e1a7a757893fdf8db1961|1.89|2014-10-31 18:10:00|1.4091206135396188|1|2700038811|273|0.612062184999033|0|47|257|-80.7007|39|35.06858|TOMATOES|0.0|1|HUNTS TOMATO PASTE 12 OZ.|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00027000388112|VEGETABLES-CAN/JAR|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|a679fa5789bfa57a05c8129e8b286de13580f0d0|2.19|2015-03-03 15:36:00|1.4091206135396188|1|1200000230|273|0.612062184999033|0|47|55|-80.7007|8|35.06858|REGULAR|1.2|23|DR WHAM 2 LTR|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00071854000546|CARBONATED BEVERAGES|BEVERAGE|-80.7007|1.4084929236641879|273|1
35.06858|50eddc40f754582a2effb2d4d618e7eb9529dac7|2.19|2015-01-27 16:51:00|1.4091206135396188|1|1200000230|273|0.612062184999033|0|47|55|-80.7007|8|35.06858|REGULAR|1.2|23|DR WHAM 2 LTR|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00071854000546|CARBONATED BEVERAGES|BEVERAGE|-80.7007|1.4084929236641879|273|1
35.06858|ae566205f2f42ba1377243cd838f96a835e56e1a|2.19|2015-01-06 21:30:00|1.4091206135396188|1|7203670293|273|0.612062184999033|0|47|423|-80.7007|72|35.06858|NFS-DISPOSE PLATES/BOWLS|0.3|1|YH FOAM BOWLS 12 OZ|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036702937|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|a39c46ad636cc758f380dff25c83abef070e4e83|6.79|2014-11-06 16:31:00|1.4091206135396188|1|7064003404|273|0.612062184999033|0|47|252|-80.7007|45|35.06858|PREMIUM ICE CREAM|2.81|5|B BUNNY PREM PNUT BUTTER PANIC|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00070640034086|ICE CREAM|FROZEN|-80.7007|1.4084929236641879|273|1
35.06858|a7d2f0edb5f077e4aa029b7ba30187fbd656f559|3.55|2014-11-05 18:33:00|1.4091206135396188|1|7433610102|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HIGHLAND CREST 2% REDUCE FAT|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00074336101021|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|4a29b8c4d6baf6fc43bdf7edeadaef22a103c6ff|2.19|2014-10-16 18:31:00|1.4091206135396188|1|1200000230|273|0.612062184999033|0|47|55|-80.7007|8|35.06858|REGULAR|0.2|23|DR PEPPER 2 LITER|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00078000082463|CARBONATED BEVERAGES|BEVERAGE|-80.7007|1.4084929236641879|273|1
35.06858|804f7ae9be7b22f9fb56cd65ac63fbf48f0249df|3.19|2014-10-03 06:22:00|1.4091206135396188|1|8265741157|273|0.612062184999033|0|47|31|-80.7007|4|35.06858|NON CARBONATED WATER|0.69|1|DEER PARK SPR WATER HALF PINT|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00082657411576|BOTTLED WATER|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|d795908d864efa77764793777acbb3c35232b5af|3.55|2014-10-23 18:32:00|1.4091206135396188|1|7433610102|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HIGHLAND CREST 2% REDUCE FAT|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00074336101021|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|ac816ad9dfd4f66c82202fe1a299bac14469ef2d|4.79|2014-11-26 12:12:00|80.700712769248256|1|1200010041|273|35.077874297799774|0|42|54|-80.64817|8|35.04711|DIET|2.39|23|DIET PEPSI COLA 16OZ NR|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|35.088667338853092|00012000100413|CARBONATED BEVERAGES|BEVERAGE|-80.7007|80.700700160737696|129|1
35.06858|a1aad52d28eded449e472da64b4660b3c9939714|9.58|2015-01-07 17:23:00|1.4091206135396188|1|1200010041|273|0.612062184999033|0|47|54|-80.7007|8|35.06858|DIET|2.4|23|DIET PEPSI COLA 16OZ NR|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00012000100413|CARBONATED BEVERAGES|BEVERAGE|-80.7007|1.4084929236641879|273|2
35.06858|863de8af5d1879e10a7a9fdfb83ad9934bc017fa|1.69|2015-01-08 22:21:00|80.700712769248256|1|1200000129|273|35.077874297799774|0|42|55|-80.64817|8|35.04711|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|35.088667338853092|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.7007|80.700700160737696|129|1
35.06858|9d7b1bdf71cd2ba0a133209123404093c5829c89|9.58|2015-01-15 17:40:00|1.4091206135396188|1|1200010041|273|0.612062184999033|0|47|54|-80.7007|8|35.06858|DIET|2.39|23|DIET PEPSI COLA 16OZ NR|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00012000100413|CARBONATED BEVERAGES|BEVERAGE|-80.7007|1.4084929236641879|273|2
35.06858|3647419f0870bbc3653c043cbd343c459b9b4f9a|9.58|2015-02-04 17:14:00|1.4091206135396188|1|1200010041|273|0.612062184999033|0|47|54|-80.7007|8|35.06858|DIET|2.39|23|DIET PEPSI COLA 16OZ NR|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00012000100413|CARBONATED BEVERAGES|BEVERAGE|-80.7007|1.4084929236641879|273|2
35.06858|7971ce11be5d0a98f373f081c7d9760f97f5e571|5.98|2014-12-17 19:10:00|1.4091206135396188|1|1117962067|273|0.612062184999033|0|47|7407|-80.7007|1600|35.06858|CHRISTMAS PARTY GOODS/DECOR|1.0|18|I/O RED/GM PDOT CELLO BAGS|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00011179620678|SEASONAL MERCHANDISE|GM|-80.7007|1.4084929236641879|273|2
35.06858|4a7bb7ddf3b53cdbb796fdd812f5c0b72f26ed3f|4.89|2014-09-27 14:37:00|1.4091206135396188|1|30149003908|273|0.612062184999033|0|47|4418|-80.7007|1210|35.06858|ANTINAUSEA REMEDY-LIQUID|0.9|17|PEPTO-BISMOL LIQUID  -03908|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00301490039083|STOMACH REMEDIES|HBC|-80.7007|1.4084929236641879|273|1
35.06858|046f405c46d18cf08f2dbc40e525a6f5146ebeb4|5.99|2014-12-17 21:43:00|1.4091206135396188|1|7756725423|273|0.612062184999033|0|47|275|-80.7007|45|35.06858|SUPER PREMIUM ICE CREAM|2.99|5|BREYERS BLASTS M&MS|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00077567300072|ICE CREAM|FROZEN|-80.7007|1.4084929236641879|273|1
35.06858|f30adc17bcda4db6e4b9bc103f4f3d58fe739eec|7.98|2014-10-23 21:08:00|1.4091206135396188|1|7279600271|273|0.612062184999033|0|47|55|-80.7007|8|35.06858|REGULAR|1.98|23|IBC CREAM SODA 6PK|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072796990001|CARBONATED BEVERAGES|BEVERAGE|-80.7007|1.4084929236641879|273|2
35.06858|442f9b1f04f0b6382b39956d7fa17dd4117453ba|11.99|2015-02-05 13:27:00|1.4091206135396188|1|7726006273|273|0.612062184999033|0|47|727|-80.7007|7|35.06858|SEASONAL CANDY-SINGLE FAC|3.0|1|I/O(V15)RS PECAN DELIGHT HEART|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00077260062734|CANDY|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|706b7ff52c9aca526f3b33491566516178308b31|2.27|2014-12-31 14:35:00|1.4091206135396188|1|7203656065|273|0.612062184999033|0|47|315|-80.7007|52|35.06858|CHEESE-PROCESSED-SLICED|0.0|3|HT SINGLE WRAP CHEESE|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|0.61242566243833529|00072036560650|CHEESE|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|d3d38aa8087874f04a5805fc82beb2f185a94a99|12.76|2014-11-06 08:05:00|80.700712769248256|1|2520000109|273|35.077874295458152|0|42|236|-80.699686|38|35.000049|DRY BEANS|0.0|1|HURST SOUP MIX CAJUN 15 BEANS|fd8b6c9ae459387db92dfe347eb96b528b999b30|0.6422135331034634|35.088667338853092|00025200001145|RICE GRAINS AND BEANS|G1 GROCERY|-80.7007|80.700708062916888|249|4
35.103409|44114d690189d8880e437b60f26dce2ad0f1bf16|2.0|2014-11-23 14:40:00|1.4132775322775095|4|4300000953|88|0.6126700657242101|0|58|272|-80.992182|307|35.103409|TOPPINGS FROZEN|1.01|5|COOL WHIP WHIPPED TOPPING|fe0b3ff9e82c459b51e7b5d07108b224a7f2607f|0.8776114689600995|0.61177642288969325|00043000009536|DESSERTS FROZEN|FROZEN|-80.992182|1.413580244274486|88|1
35.103409|65d8d25830502ac34aa1e6b78e82d3c8eaeeaf7d|2.19|2014-12-07 15:42:00|1.4132775322775095|4|4900005010|88|0.6126700657242101|0|58|55|-80.992182|8|35.103409|REGULAR|0.69|23|D FUZE ICE TEA LEMON 2 LITER|fe0b3ff9e82c459b51e7b5d07108b224a7f2607f|0.8776114689600995|0.61177642288969325|00080793808571|CARBONATED BEVERAGES|BEVERAGE|-80.992182|1.413580244274486|88|1
35.103409|42bb68677062882f720b5480e01234d2368a635f|8.19|2015-02-17 17:42:00|1.4132775322775095|4|5150004817|88|0.6126700657242101|0|58|1270|-80.992182|41|35.103409|SWEET BREAKFAST|0.0|5|SMUCKER PB&GRAPE UNCRUSTABLES|fe0b3ff9e82c459b51e7b5d07108b224a7f2607f|0.8776114689600995|0.61177642288969325|00051500048177|BREAKFAST FOODS FROZEN|FROZEN|-80.992182|1.413580244274486|88|1
35.103409|188d8dbb38aba53f4c70d0dc8b8e3e6b3e013213|8.19|2015-02-25 20:47:00|1.4132775322775095|4|5150004817|88|0.6126700657242101|0|58|1270|-80.992182|41|35.103409|SWEET BREAKFAST|0.0|5|SMUCKER PB&GRAPE UNCRUSTABLES|fe0b3ff9e82c459b51e7b5d07108b224a7f2607f|0.8776114689600995|0.61177642288969325|00051500048177|BREAKFAST FOODS FROZEN|FROZEN|-80.992182|1.413580244274486|88|1
35.103409|a58360cc53948cb02377b947475d73578c18e1e7|2.0|2014-10-31 18:23:00|1.4132775322775095|4|2840000210|88|0.6126700657242101|0|58|204|-80.992182|31|35.103409|TORTILLA CHIPS|0.0|1|SANTITAS BLENDED CORN|fe0b3ff9e82c459b51e7b5d07108b224a7f2607f|0.8776114689600995|0.61177642288969325|00028400002110|SNACKS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|818d425045392a219b66e28909e815b09dce4f2c|1.69|2015-03-08 21:47:00|1.4132775322775095|4|7203688003|88|0.6126700657242101|0|58|527|-80.992182|64|35.103409|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|fe0b3ff9e82c459b51e7b5d07108b224a7f2607f|0.8776114689600995|0.61177642288969325|00072036880031|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|1
35.103409|a935fd4a9cd91a384ebeba756ee6c21b81f28dee|8.99|2014-09-22 20:32:00|1.4132775322775095|4|31254742592|88|0.6126700657242101|0|58|4039|-80.992182|1080|35.103409|ORAL RINSE WHITENING|0.0|17|LISTERINE WHT/RESTOR FLOU RNSE|fe0b3ff9e82c459b51e7b5d07108b224a7f2607f|0.8776114689600995|0.61177642288969325|00312547425926|ORAL HYGIENE|HBC|-80.992182|1.413580244274486|88|1
35.103409|90424bfab7b2beb30f17b6a2282d7db53f25fd7f|1.79|2014-09-11 17:42:00|1.4132775322775095|4|7339000393|88|0.6126700657242101|0|58|48|-80.992182|7|35.103409|REGISTER GUM|0.5|1|MENTOS FRESH MINT GUM 15CT|fe0b3ff9e82c459b51e7b5d07108b224a7f2607f|0.8776114689600995|0.61177642288969325|00073390013936|CANDY|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|9aea448dc32b9083e9d59871ea609f23ce963f67|0.94|2015-02-06 20:32:00|1.4132775322775095|4|1310077027|88|0.6126700657242101|0|58|426|-80.992182|72|35.103409|NFS-PAPER TOWELS|0.0|1|SPA PAPER TOWEL|fe0b3ff9e82c459b51e7b5d07108b224a7f2607f|0.8776114689600995|0.61177642288969325|00013100770278|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|fce89d4f7d87fee652cfd234c20b807a95d9ce8f|3.58|2014-09-13 20:40:00|1.4132775322775095|4|2430004101|88|0.6126700657242101|0|58|1044|-80.992182|173|35.103409|SW BAKD GOOD SNACK CAKES|0.29|7|LD HONEY BUNS|fe0b3ff9e82c459b51e7b5d07108b224a7f2607f|0.8776114689600995|0.61177642288969325|00024300041020|SWEET BAKED GOODS|COMMERCIAL BAKERY|-80.992182|1.413580244274486|88|2
35.103409|ab072678fcc0b245910c39d07cf13fb87aae970d|4.29|2014-10-27 20:32:00|1.4132775322775095|4|1090000015|88|0.6126700657242101|0|58|440|-80.992182|76|35.103409|NFS-ALUMINUM FOIL|1.29|1|REYNOLDS FOIL HEAVY DUTY 50 FT|fe0b3ff9e82c459b51e7b5d07108b224a7f2607f|0.8776114689600995|0.61177642288969325|00010900000215|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|1309cf9fc15e7634907ff784e9d404d1ac137cc6|2.67|2014-10-26 18:44:00|1.4132775322775095|4|7064000461|88|0.6126700657242101|0|58|275|-80.992182|45|35.103409|SUPER PREMIUM ICE CREAM|0.34|5|B BUNNY PERSONL PNUT BTR PANIC|fe0b3ff9e82c459b51e7b5d07108b224a7f2607f|0.8776114689600995|0.61177642288969325|00070640004638|ICE CREAM|FROZEN|-80.992182|1.413580244274486|88|2
35.333742|0c2d26000f86e26ed25b655ef9aeed8376086888|3.55|2014-11-27 07:29:00|80.780380710856576|4|7433610102|472|35.370498620627068|0|48|342|-80.764523|57|35.341927|FRESH MILK|0.0|3|HIGHLAND CREST 2% REDUCE FAT|0ab57bd802d6bfb89c0f7801010291abc6abbefb|2.5397938437587544|35.351085445956379|00074336101021|MILK|DAIRY|-80.814133|80.814146996411907|220|1
35.116638|9cc8bc6087e59585f720476ad5f4e61af2dfcbff|9.98|2015-02-04 18:19:00|80.856688219393845|4|7203688080|204|35.134105651841615|0|15|523|-80.699686|64|35.000049|FRESH POTATOES|2.49|4|HT YUKON GOLD 5 LB BAG|0ad59eeb4dc3a7e24e7a01350db474e915028845|1.2069727108377397|35.134355925261694|00072036880802|FRESH PRODUCE|PRODUCE|-80.85753|80.857540698893658|249|2
35.116638|cf2e9ddcc902200e82c6e1badaec113050eb2898|2.71|2014-12-23 19:07:00|80.856688219393845|4||204|35.134105651841615|0|15|522|-80.699686|64|35.000049|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|0ad59eeb4dc3a7e24e7a01350db474e915028845|1.2069727108377397|35.134355925261694|00204664000004|FRESH PRODUCE|PRODUCE|-80.85753|80.857540698893658|249|1
35.116638|da2838e8d50d79a3c347769ef5c4bc4a6e10ec76|0.51|2014-11-01 19:45:00|80.856688219393845|4||204|35.134105651841615|0|15|522|-80.699686|64|35.000049|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|0ad59eeb4dc3a7e24e7a01350db474e915028845|1.2069727108377397|35.134355925261694|00204664000004|FRESH PRODUCE|PRODUCE|-80.85753|80.857540698893658|249|1
35.116638|4684780f2dc10dc3a9702e96a136b077c2f67c4c|4.99|2014-10-25 15:19:00|80.856688219393845|4|7023430470|204|35.134105651841615|0|15|1220|-80.699686|275|35.000049|PASTA SC PREMIUM|0.0|1|GINA PASTA SC VODKA|0ad59eeb4dc3a7e24e7a01350db474e915028845|1.2069727108377397|35.134355925261694|00070234304502|PASTA SAUCES|G1 GROCERY|-80.85753|80.857540698893658|249|1
35.116638|ede930afeea73424283b478bd9e1cb7d16a3bbaa|4.69|2014-10-16 21:49:00|80.856688219393845|4|4900002468|204|35.134105651841615|0|15|54|-80.699686|8|35.000049|DIET|0.0|23|COKE ZERO .5L 6PK PET|0ad59eeb4dc3a7e24e7a01350db474e915028845|1.2069727108377397|35.134355925261694|00049000045840|CARBONATED BEVERAGES|BEVERAGE|-80.85753|80.857540698893658|249|1
35.116638|acd4447b3d9cc973fd62cb2e721e869e239431be|1.99|2014-10-12 10:57:00|80.856688219393845|4|4069503007|204|35.134105651841615|0|15|555|-80.699686|64|35.000049|PACKAGED SALADS|0.0|4|ROMIANE HEARTS|0ad59eeb4dc3a7e24e7a01350db474e915028845|1.2069727108377397|35.134355925261694|00033383651620|FRESH PRODUCE|PRODUCE|-80.85753|80.857540698893658|249|1
35.116638|9f908a64085e292d6f82ee43dad42fa1fbcb27e9|1.29|2014-11-15 14:15:00|80.856688219393845|4|7152416007|204|35.134105651841615|0|15|1214|-80.699686|272|35.000049|AUTHENTIC HISPANIC|0.0|1|LA PREF GREEN CHILE DICED|0ad59eeb4dc3a7e24e7a01350db474e915028845|1.2069727108377397|35.134355925261694|00071524160075|HISPANIC PREP. FOODS|G1 GROCERY|-80.85753|80.857540698893658|249|1
35.116638|7e6b13a87d4de993ca9a675c1c4c35ea491b6bfd|0.99|2014-10-11 12:00:00|80.856688219393845|4|7203698291|204|35.134105651841615|0|15|245|-80.699686|39|35.000049|VEGETABLES-CORE|0.22|1|HT CORN WK GOLDEN|0ad59eeb4dc3a7e24e7a01350db474e915028845|1.2069727108377397|35.134355925261694|00072036411815|VEGETABLES-CAN/JAR|G1 GROCERY|-80.85753|80.857540698893658|249|1
35.116638|43183c9f2ed3fe19670623d4962d29f9143db5d2|6.1|2014-11-15 14:30:00|80.856688219393845|4|20895100000|204|35.134105651841615|0|15|977|-80.699686|201|35.000049|FRESH HT CHICKEN|0.0|2|HT FRESH CHICKEN THIGHS|0ad59eeb4dc3a7e24e7a01350db474e915028845|1.2069727108377397|35.134355925261694|00208951000005|POULTRY|MEAT|-80.85753|80.857540698893658|249|1
35.116638|ddcf1d30e1b078c9a1f04704b763297bec64ed56|2.0|2015-01-24 18:32:00|80.856688219393845|4|2500004748|204|35.134105651841615|0|15|338|-80.699686|56|35.000049|OTHER FRUIT JUICES|0.0|3|MINUTE MAID LEMONADE|0ad59eeb4dc3a7e24e7a01350db474e915028845|1.2069727108377397|35.134355925261694|00025000047480|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.85753|80.857540698893658|249|1
35.116638|be4f9c28e6415b664df0f4113d3a75cac37ac370|1.68|2014-11-09 17:22:00|80.856688219393845|4|20401600000|204|35.134105651841615|0|15|500|-80.699686|64|35.000049|FRESH APPLES|0.0|4|RED DEL APPLES  72|0ad59eeb4dc3a7e24e7a01350db474e915028845|1.2069727108377397|35.134355925261694|00891658001163|FRESH PRODUCE|PRODUCE|-80.85753|80.857540698893658|249|1
35.116638|52ef70ab5491aa3698537bd0a240ee73a35c8dbc|2.19|2015-02-15 15:52:00|80.856688219393845|4|76857300210|204|35.134105651841615|0|15|544|-80.699686|64|35.000049|FRESH PRODUCE FRSH HERBS|0.0|4|PKG FRESH MINT|0ad59eeb4dc3a7e24e7a01350db474e915028845|1.2069727108377397|35.134355925261694|00768573001106|FRESH PRODUCE|PRODUCE|-80.85753|80.857540698893658|249|1
35.116638|38fc47ac72ae8e3a50719327e68dc1852c562976|4.49|2014-11-18 20:31:00|80.856688219393845|4|4000041331|204|35.134105651841615|0|15|727|-80.699686|7|35.000049|SEASONAL CANDY-SINGLE FAC|0.5|1|I/O(C14)DOVE AST CHOC CHRISTMS|0ad59eeb4dc3a7e24e7a01350db474e915028845|1.2069727108377397|35.134355925261694|00040000413318|CANDY|G1 GROCERY|-80.85753|80.857540698893658|249|1
35.116638|b9a9875363e99b53574f21f326de85d33252006b|3.69|2014-11-19 19:10:00|80.856688219393845|4|78142117010|204|35.134105651841615|0|15|1609|-80.699686|371|35.000049|TAKE & BAKE BREAD|0.7|14|LB TAKE/BAKE RUST CIABATT ROLL|0ad59eeb4dc3a7e24e7a01350db474e915028845|1.2069727108377397|35.134355925261694|00781421170076|BREAD|BAKERY|-80.85753|80.857540698893658|249|1
35.116638|b2c9ae6276cc2604ff4fe96573aadd7a5fff6bea|1.5|2014-10-18 10:33:00|80.856688219393845|4||204|35.134105651841615|0|15|1617|-80.699686|373|35.000049|ROLLS BULK|0.0|14|BULK ROLLS|0ad59eeb4dc3a7e24e7a01350db474e915028845|1.2069727108377397|35.134355925261694|00072036955555|ROLLS|BAKERY|-80.85753|80.857540698893658|249|2
35.116638|b490952281fecd95dc1d28fbb28a82411367a410|7.38|2014-12-31 17:38:00|80.856688219393845|4|4300095051|204|35.134105651841615|0|15|209|-80.699686|20|35.000049|POWDERED SOFT DRINKS|0.69|1|CRYSTAL LT GRN TEA PCH MANGO|0ad59eeb4dc3a7e24e7a01350db474e915028845|1.2069727108377397|35.134355925261694|00043000028858|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.85753|80.857540698893658|249|2
35.116638|7ee9e7b6868f114f65b31755d27c99a804b7540f|1.72|2014-12-24 16:22:00|80.856688219393845|4||204|35.134105651841615|0|15|500|-80.699686|64|35.000049|FRESH APPLES|0.0|4|RED DEL APPLE, WA  48|0ad59eeb4dc3a7e24e7a01350db474e915028845|1.2069727108377397|35.134355925261694|00233284000002|FRESH PRODUCE|PRODUCE|-80.85753|80.857540698893658|249|1
35.116638|2e44938108ad311d20f43a60178443fbf6465b26|4.99|2015-01-11 12:36:00|80.856688219393845|4|2840008313|204|35.134105651841615|0|15|204|-80.699686|31|35.000049|TORTILLA CHIPS|1.0|1|TOSTITOS RSTC FAMILY SIZE|0ad59eeb4dc3a7e24e7a01350db474e915028845|1.2069727108377397|35.134355925261694|00028400083133|SNACKS|G1 GROCERY|-80.85753|80.857540698893658|249|1
35.195689|8ceee2a2a55ed514c277de5032953dce6fb13c1b|7.98|2014-12-03 12:42:00|1.4094857484078087|1|3338324028|412|0.6142806555579505|0|26|504|-80.826724|64|35.195689|FRESH BERRIES|4.64|4|BLACKBERRIES 5.6 OZ|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00761635202602|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|2
35.195689|de3537eaead7369a2cd16c93cc54a8ba309ef605|4.29|2014-10-22 14:40:00|1.4094857484078087|1|70875800101|412|0.6142806555579505|0|26|8|-80.826724|2|35.195689|BROWNIE MIXES|0.0|1|NO PUDGE FF ORIGINAL BROWNIE|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00708758001019|BAKING MIXES|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|afe98c59e898ba50af0f85f442be443c8a0911f3|4.29|2015-01-26 13:30:00|1.4094857484078087|1|70875800101|412|0.6142806555579505|0|26|8|-80.826724|2|35.195689|BROWNIE MIXES|0.0|1|NO PUDGE FF ORIGINAL BROWNIE|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00708758001019|BAKING MIXES|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|7e19b95a2f648b5fffce81898e857eb76c047246|2.2|2014-10-19 17:38:00|1.4094857484078087|1|20631400000|412|0.6142806555579505|0|26|1825|-80.826724|410|35.195689|BH SALAMI|0.0|6|BH SLICED HARD SALAMI|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00205938000003|BH MEAT|DELI|-80.826724|1.4106924574007214|412|1
35.195689|46612f2c1ee50c073a3c5810513c9bbcf1f5a5b3|1.4|2014-12-24 14:34:00|1.4094857484078087|1||412|0.6142806555579505|0|26|524|-80.826724|64|35.195689|FRESH PROD FRESH ONIONS|0.0|4|COO SHALLOTS, BULK|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00204662000006|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|1
35.195689|246cf4ef5bb07e08283c2af1bbb6abb674fdc3dc|0.75|2015-01-25 15:30:00|1.4094857484078087|1||412|0.6142806555579505|0|26|502|-80.826724|64|35.195689|FRESH BANANAS|0.0|4|REWRAP BANANAS BY POUND|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00204186000001|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|1
35.195689|6bb2c8d94a6ab9c7fe6702418d8a7bb78f69a632|1.89|2014-11-26 09:00:00|1.4094857484078087|1|4010000928|412|0.6142806555579505|1|26|29|-80.826724|3|35.195689|REMAINING BAKING SUPPLIES|0.0|1|FLEISCHMAN YEAST PACKETS|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00040100009282|BAKING SUPPLIES|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|bfe281ed5c95d1d24afc61371936aa79a9c9ed70|1.79|2015-03-07 10:26:00|1.4094857484078087|1|5200013446|412|0.6142806555579505|0|26|171|-80.826724|20|35.195689|ISOTONIC DRINKS|0.54|1|GATORADE CHEWS FRUITPUNCH|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00052000134469|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|eda8ed886a8490901014385c4659c4bd98b3c147|3.38|2014-12-05 11:01:00|80.828402574597021|1|4430010632|412|35.205805381648155|0|8|1212|-80.85013|272|35.175855|HISP BEANS/PEPPERS|0.0|1|ROSARITA REFRIED BEANS FF TRAD|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|35.209978091326001|00044300106222|HISPANIC PREP. FOODS|G1 GROCERY|-80.826724|80.826727865697862|218|2
35.195689|450a96c6015452a1adbc9fab431ebdf6faad8efc|5.49|2015-03-05 14:05:00|1.4094857484078087|1|6827443227|412|0.6142806555579505|0|26|31|-80.826724|4|35.195689|NON CARBONATED WATER|1.5|1|NESTLE WATER 24PK 8 OZ|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00068274432279|BOTTLED WATER|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|a16843e026b587361ec03ded68319f25d9648438|5.59|2015-03-01 16:15:00|1.4094857484078087|1|5210003025|412|0.6142806555579505|0|26|220|-80.826724|34|35.195689|PEPPER|0.0|1|MC COARSE GROUND PEPPER|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00052100071268|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|74bceac324d3cb80553a496de0928f048bd93e44|6.99|2014-10-17 09:22:00|1.4094857484078087|1|7580587487|412|0.6142806555579505|0|26|2019|-80.826724|505|35.195689|PRESSED COOKED CHEESE|3.5|6|STELLA ROMANO WEDGE|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00075805874873|SPECIALTY CHEESE|DELI|-80.826724|1.4106924574007214|412|1
35.195689|71c2644464f41482c6be0e4a10a4f95d2e6bc628|5.99|2014-09-26 12:59:00|1.4094857484078087|1|7580582046|412|0.6142806555579505|0|26|2021|-80.826724|505|35.195689|FRESH CHEESE|2.0|6|STELLA BLUE CHEESE CRUMBLES|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00075805820467|SPECIALTY CHEESE|DELI|-80.826724|1.4106924574007214|412|1
35.195689|06a89412e949a15ae77a6e7e37c3de91d929fd2c|3.49|2014-12-11 09:27:00|1.4094857484078087|1|7203670903|412|0.6142806555579505|0|26|214|-80.826724|33|35.195689|BROTH|0.49|1|HT RED SODIUM CHICK BROTH 48OZ|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00072036709042|SOUP|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|711b8511ef1f355076ed511847603561ac0a9513|2.89|2015-02-23 19:38:00|1.4094857484078087|1|7203695917|412|0.6142806555579505|0|26|1625|-80.826724|373|35.195689|FROZEN DOUGH (ROLLS)|0.0|14|FRESH CHICAGO ROLL|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00072036959171|ROLLS|BAKERY|-80.826724|1.4106924574007214|412|1
35.195689|7bf64cdc8c089ad3d1ecf1a52f33acc9c5a22b9d|6.19|2014-12-20 16:25:00|1.4094857484078087|1|2800021560|412|0.6142806555579505|0|26|16|-80.826724|3|35.195689|BAKING CHOCOLATE/CHIPS/MORSELS|0.6|1|NESTLE SEMISWEET MORSELS|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00028000215606|BAKING SUPPLIES|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|7a20a5afec397f209832b303686dd7ab85e6a33b|11.07|2014-11-12 14:13:00|1.4094857484078087|1|1630015353|412|0.6142806555579505|0|26|139|-80.826724|20|35.195689|REMAINING SHELF STABLE JUICES|0.0|1|DD UNSWEET GRAPEFRT JUICE 6PK|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00016300153537|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.826724|1.4106924574007214|412|3
35.195689|73cecba204580fc07e074367f16bb3ea77320b95|2.75|2014-12-14 15:56:00|1.4094857484078087|1|2800021010|412|0.6142806555579505|1|26|16|-80.826724|3|35.195689|BAKING CHOCOLATE/CHIPS/MORSELS|0.25|1|NESTLE TOLL HOUSE CHOC CHUNK|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00028000210205|BAKING SUPPLIES|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|464f39f37cc53ad764ac8513b48c566ca251fc27|3.19|2015-01-17 16:21:00|1.4094857484078087|1|2800021010|412|0.6142806555579505|0|26|16|-80.826724|3|35.195689|BAKING CHOCOLATE/CHIPS/MORSELS|0.0|1|NESTLE SEMISWEET MORSELS|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00028000215804|BAKING SUPPLIES|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|e3bc04aefb0854859f375d1bef8e4fc061134c35|12.38|2014-12-18 10:00:00|80.828402574597021|1|2800021560|412|35.205805381648155|0|8|16|-80.85013|3|35.175855|BAKING CHOCOLATE/CHIPS/MORSELS|1.2|1|NESTLE SEMISWEET MORSELS|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|35.209978091326001|00028000215606|BAKING SUPPLIES|G1 GROCERY|-80.826724|80.826727865697862|218|2
35.195689|1f21d87a0ac172aa5318edf30972d8b23fcc1f66|12.0|2014-12-09 18:42:00|1.4094857484078087|1|66440177739|412|0.6142806555579505|0|26|1165|-80.826724|87|35.195689|NFS-FRESH CONSUMER BUNCH|0.0|9|BUNCH- JUMBO SUNFLOWER 3 ST|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00664401777390|FLORAL|FLORAL|-80.826724|1.4106924574007214|412|3
35.195689|e2688ca9298c8b0e76ed361277cd09d68c97e477|5.89|2015-01-13 14:46:00|1.4094857484078087|1|30081073088|412|0.6142806555579505|1|26|4844|-80.826724|1235|35.195689|FIRST AID TREATMENT|0.0|17|(JHK) NEOSPORIN ORIG OINTMENT|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00300810730884|FIRST AID|HBC|-80.826724|1.4106924574007214|412|1
35.195689|2d55e5c959adc1f3deb9d63b096f2c58effa96a6|4.99|2015-02-09 12:36:00|1.4094857484078087|1|71575620002|412|0.6142806555579505|0|26|504|-80.826724|64|35.195689|FRESH BERRIES|1.49|4|STRAWBERRIES 1LB CLAM|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00715756200023|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|1
35.195689|2d07038773beec174842a2a535b55db99990b762|12.0|2014-12-24 14:52:00|80.828402574597021|1|66440177739|412|35.205805381648155|0|8|1165|-80.85013|87|35.175855|NFS-FRESH CONSUMER BUNCH|0.0|9|BUNCH- JUMBO SUNFLOWER 3 ST|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|35.209978091326001|00664401777390|FLORAL|FLORAL|-80.826724|80.826727865697862|218|3
35.195689|8bacd2604388e8a53e7bd6180570d527cf37f5bf|4.49|2014-11-06 11:40:00|80.828402574597021|1|76770700167|412|35.205805382140767|0|8|312|-80.844274|51|35.204336|BUTTER|0.9|3|KERRYGOLD SPREADABLE BUTTER|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|35.209978091326001|00767707001678|BUTTER & MARGARINE|DAIRY|-80.826724|80.826724129369339|61|1
35.195689|295c8e127208f0a4f080a993afef58fe4be928dc|4.49|2015-01-04 20:26:00|80.828402574597021|1|88491201426|412|35.205805381648155|0|8|74|-80.85013|9|35.175855|RTE CEREAL ALL FAMILY|0.0|1|POST HNY BUNCHES FAM ALMOND|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|35.209978091326001|00884912014276|CEREAL|G1 GROCERY|-80.826724|80.826727865697862|218|1
35.195689|b1a7c8791eb9983c0a4232d727b7d1828ee9707e|3.99|2014-11-22 08:38:00|1.4094857484078087|1|81793900034|412|0.6142806555579505|0|26|722|-80.826724|73|35.195689|NFS-HAND SOAPS|0.0|1|METHOD FOAM SOAP LEMON MINT|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00817939011621|PERSONAL SOAP/BATH ADDITIVES|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|aaf3f8e421f626d681f9d304eab90083fc4d523b|10.49|2015-02-15 19:43:00|1.4094857484078087|1|79849310320|412|0.6142806555579505|0|26|36|-80.826724|10|35.195689|PREMIUM GROUND|4.5|1|CARIBOU COFFEE MORNING BLEND|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00798493103673|COFFEE|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|7deecf4019c09ce2861ec19eddc1b60a2ba5f6b1|3.49|2015-01-19 10:18:00|1.4094857484078087|1|88491201424|412|0.6142806555579505|0|26|74|-80.826724|9|35.195689|RTE CEREAL ALL FAMILY|0.0|1|POST HNY BUNCHES VANLLA|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00884912017864|CEREAL|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|02e0a7f9495bc94ce165e994b070801acf9acdbc|3.89|2014-10-05 15:35:00|1.4094857484078087|1|2120059846|412|0.6142806555579505|1|26|729|-80.826724|69|35.195689|NFS-SCOUR PAD/STEEL WOOL|0.0|1|SCOTCHBRITE HEAVY DUTY SPG 3PK|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00021200572357|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|b6e4eb54ba6131329ea3302a7bb76fa1a080fc40|5.69|2015-02-25 09:50:00|1.4094857484078087|1|1708287631|412|0.6142806555579505|0|26|215|-80.826724|31|35.195689|JERKY SNACKS|0.0|1|JACK LINK'S ORIGINAL JERKY|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00017082007872|SNACKS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|83fedf56ecba0c1da88b570f1783ce552aeeeaa4|3.89|2014-09-17 15:28:00|1.4094857484078087|1|2120059846|412|0.6142806555579505|1|26|729|-80.826724|69|35.195689|NFS-SCOUR PAD/STEEL WOOL|0.0|1|SCOTCHBRITE HEAVY DUTY SPG 3PK|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00021200572357|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|fcc70d71c9294e3efad5eb9b027b128aa6997cb3|4.29|2014-09-10 12:40:00|1.4094857484078087|1|7797508215|412|0.6142806555579505|0|26|202|-80.826724|31|35.195689|PRETZELS|0.3|1|SOH 100 CAL MINI PRETZ LUNCH P|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00077975082157|SNACKS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|e04c35f4649af320ae2ff74c2b83338ed9b6e31d|1.97|2014-10-08 14:35:00|1.4094857484078087|1|7203698240|412|0.6142806555579505|1|26|442|-80.826724|76|35.195689|NFS-COOKING-STORAGE BAGS|0.0|1|YH RESEALABLE SANDWICH BAGS|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00072036982407|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|e8eaf52bceb6b41be24a1aef406fbb7c9284ebc0|2.79|2014-11-30 17:17:00|1.4094857484078087|1|7225001130|412|0.6142806555579505|0|26|1033|-80.826724|163|35.195689|HAMBURGER|0.0|7|MERITA 8PK HAMBURGER BUNS|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00072250011303|BUNS/ROLLS|COMMERCIAL BAKERY|-80.826724|1.4106924574007214|412|1
35.195689|15f3c35dd5cffa2af6ecab2f3de48b89f1df7d21|8.97|2015-02-01 15:16:00|1.4094857484078087|1|7214011020|412|0.6142806555579505|0|26|3202|-80.826724|1015|35.195689|HAND & BODY THERAPEUTIC|0.0|17|EUCERIN SMTHING ESS BDY LOTION|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00072140634827|HAND & BODY LOTION/SUN CARE|HBC|-80.826724|1.4106924574007214|412|1
35.195689|116405c7b43eacc36d80b50d0f16d3b502d52273|2.49|2015-01-05 16:51:00|1.4094857484078087|1|7373107000|412|0.6142806555579505|1|26|495|-80.826724|108|35.195689|NON REFRIGERATED|0.0|19|MISSION FAJITA 8 CT|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00073731070000|TORTILLAS|CASE READY MEATS|-80.826724|1.4106924574007214|412|1
35.195689|1fc8c3ad09a4ccae07374337789ba5062d685331|1.89|2015-02-16 15:01:00|1.4094857484078087|1|7680828008|412|0.6142806555579505|0|26|149|-80.826724|23|35.195689|WHSE PASTA CORE|0.39|1|BARILLA PASTA ANGEL HAIR|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00076808501063|PASTA|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|17035a52e9ae0b37cf521369d7e3e03087c46172|14.98|2014-12-07 15:27:00|1.4094857484078087|1|7490836026|412|0.6142806555579505|0|26|1220|-80.826724|275|35.195689|PASTA SC PREMIUM|3.75|1|DELGROSSO SC TOM BASIL|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00074908360306|PASTA SAUCES|G1 GROCERY|-80.826724|1.4106924574007214|412|2
35.195689|6392d1885b2b92415ccf8f5e409a6477d7187d4f|2.99|2015-01-11 15:11:00|1.4094857484078087|1|7203698384|412|0.6142806555579505|0|26|690|-80.826724|61|35.195689|ORGANIC|0.0|3|HTO ORGANIC VANILLA YOGURT|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00072036983848|YOGURT|DAIRY|-80.826724|1.4106924574007214|412|1
35.195689|e69998c2893d3e304d2055c62847bee482503a73|8.97|2015-03-04 16:55:00|1.4094857484078087|1|7203698384|412|0.6142806555579505|1|26|690|-80.826724|61|35.195689|ORGANIC|1.47|3|HTO ORGANIC VANILLA YOGURT|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00072036983848|YOGURT|DAIRY|-80.826724|1.4106924574007214|412|3
35.195689|f1a8edfdb4884c440c17d20bfa2ea2ed315f7b88|1.49|2015-02-06 10:55:00|1.4094857484078087|1|7203670302|412|0.6142806555579505|0|26|728|-80.826724|72|35.195689|NFS-PLASTIC FLATWARE|0.0|1|YH OCCASIONS FS FORKS|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00072036703019|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|37912ba2890a900074839a387aaa90aa1b81db50|1.69|2015-02-03 13:33:00|80.828402574597021|1|7203688003|412|35.205805381648155|0|8|527|-80.85013|64|35.175855|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|35.209978091326001|00072036880031|FRESH PRODUCE|PRODUCE|-80.826724|80.826727865697862|218|1
35.195689|7ce94f35f9a6a99240a6014df7825a487cf794cc|7.49|2014-09-29 15:03:00|80.828402574597021|1|7490836026|412|35.2058053811622|0|8|1220|-80.825175|275|35.152722|PASTA SC PREMIUM|1.5|1|DELGROSSO SC MARINARA|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|35.209978091326001|00074908360269|PASTA SAUCES|G1 GROCERY|-80.826724|80.826729446921846|160|1
35.195689|d5133907a2d89fa2155ff71fcad086fbd22641f2|10.47|2015-03-02 19:32:00|80.828402574597021|1|8087800218|412|35.205805381648155|0|8|3548|-80.85013|1045|35.175855|HAIR CARE SHPOO 2 IN 1'S|0.47|17|PANTENE SHAM 2N1 CLASSIC CLEAN|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|35.209978091326001|00080878004065|HAIR & SCALP CARE|HBC|-80.826724|80.826727865697862|218|3
35.195689|c21d6fa1128ae3b925fad9893a7d59e85e1b3dc0|6.98|2015-02-08 17:12:00|1.4094857484078087|1|20455000000|412|0.6142806555579505|0|26|542|-80.826724|64|35.195689|FRESH VEGETABLES REMAIN|0.0|4|BRUSSEL SPROUTS 1LB (RPC)|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00094922577160|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|2
35.195689|63acc84c1a0cd98f4e96de10d7f7da836329b2b1|6.98|2015-01-28 11:33:00|1.4094857484078087|1|20455000000|412|0.6142806555579505|0|26|542|-80.826724|64|35.195689|FRESH VEGETABLES REMAIN|0.0|4|BRUSSEL SPROUTS 1LB (RPC)|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00094922577160|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|2
35.195689|fd7464b6e72683f8203cd9db9145140f1b8a505a|3.49|2015-03-03 12:42:00|1.4094857484078087|1|20455000000|412|0.6142806555579505|0|26|542|-80.826724|64|35.195689|FRESH VEGETABLES REMAIN|0.0|4|BRUSSEL SPROUTS 1LB (RPC)|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00094922577160|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|1
35.195689|6862fbc5e817f8885f2c492213e9fbfbcf2c210f|3.49|2015-01-20 16:48:00|1.4094857484078087|1|20455000000|412|0.6142806555579505|0|26|542|-80.826724|64|35.195689|FRESH VEGETABLES REMAIN|0.0|4|BRUSSEL SPROUTS 1LB (RPC)|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00094922577160|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|1
35.195689|d937885fd39b1af4b7e08bcb6566504d3eeed4a5|5.29|2014-11-01 15:55:00|1.4094857484078087|1|85103500301|412|0.6142806555579505|0|26|244|-80.826724|43|35.195689|BETTER-FOR-YOU NOVELTIES|0.0|5|YASSO YOG MINT CHOCOLATE BARS|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00851035003234|FROZEN NOVELTIES|FROZEN|-80.826724|1.4106924574007214|412|1
35.195689|f86440a5917372e794f1e2f8699dfc2117f8e5ff|4.0|2015-01-15 08:29:00|1.4094857484078087|1|84115200734|412|0.6142806555579505|0|26|1165|-80.826724|87|35.195689|NFS-FRESH CONSUMER BUNCH|0.66|9|BUNCH- 3/$12 NOVELTY POMS|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00841152007345|FLORAL|FLORAL|-80.826724|1.4106924574007214|412|1
35.195689|9898a9ab0eaa5de069ce9d32bd0c91ca878a5789|7.75|2014-11-16 16:15:00|1.4094857484078087|1|1258760034|412|0.6142806555579505|0|26|443|-80.826724|76|35.195689|NFS-GARBAGE BAGS|0.4|1|GLAD FF ODOR SHIELD TALL KTCH|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00012587703205|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|d090ae968001548456ab9c6178ff8da363e1eb70|3.95|2015-02-20 16:14:00|1.4094857484078087|1|1410007467|412|0.6142806555579505|0|26|1025|-80.826724|162|35.195689|WHITE|0.0|7|PEP FH SOURDOUGH WP BRD PP|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00014100074670|SLICED BREAD|COMMERCIAL BAKERY|-80.826724|1.4106924574007214|412|1
35.195689|d478ec777009298f2b2feed1f5a2737592d804e9|8.89|2015-02-09 16:37:00|1.4094857484078087|1|1410009655|412|0.6142806555579505|0|26|87|-80.826724|13|35.195689|CHEESE CRACKERS|1.9|1|PF BULK GOLDFISH CHEDDAR|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00014100096559|CRACKERS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|99310e15cc45acf0a5fa50e747403e25eefdae81|23.49|2015-02-02 11:07:00|80.828402574597021|1|1901461081|412|35.2058053811622|0|8|156|-80.825175|24|35.152722|NFS-DOG FOOD-DRY|0.0|1|IAMS DOG CHUNKS DRY|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|35.209978091326001|00019014610815|PET FOOD/SUPPLIES|G1 GROCERY|-80.826724|80.826729446921846|160|1
35.195689|2daca5bd56c82e2460e0586663de0551478e9ac3|3.29|2014-09-23 18:43:00|1.4094857484078087|1|7287827570|412|0.6142806555579505|0|26|1211|-80.826724|272|35.195689|HISP SALSA/DIPS|0.0|1|HERDEZ SALSA CASERA MILD|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00072878275514|HISPANIC PREP. FOODS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|51139cd7cc97ec484b38f4c456585090bf7bf917|6.99|2014-10-10 14:58:00|1.4094857484078087|1|7580587490|412|0.6142806555579505|0|26|2018|-80.826724|505|35.195689|PRESSED CHEESE|3.5|6|STELLA FONTINELLA WEDGE|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00075805874903|SPECIALTY CHEESE|DELI|-80.826724|1.4106924574007214|412|1
35.195689|38014c8843f065580edf01d31cc58827fd365195|3.89|2014-10-03 13:24:00|1.4094857484078087|1|7910094203|412|0.6142806555579505|0|26|155|-80.826724|24|35.195689|NFS-DOG TREATS|0.0|1|MILKBONE GRAVY BONES|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00079100942039|PET FOOD/SUPPLIES|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|07505c6716e81fd125d2b84b4fbc7ba01f1722e5|3.99|2014-10-14 14:10:00|80.828402574597021|1|71514151464|412|35.2058053811622|0|8|364|-80.825175|55|35.152722|ORGANIC AND CF EGGS|0.4|3|EGGLAND'S BEST CAGE FREE LARGE|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|35.209978091326001|00715141514643|EGGS FRESH|DAIRY|-80.826724|80.826729446921846|160|1
35.195689|b19bb94de4177a8dd8c4cd08af432c81611892fa|3.99|2015-03-08 20:36:00|1.4094857484078087|1|30041060686|412|0.6142806555579505|0|26|4056|-80.826724|1080|35.195689|TOOTH BRUSH-PREMIUM|1.0|17|ORAL B INDICATOR TWIN SOFT #17|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00300410606862|ORAL HYGIENE|HBC|-80.826724|1.4106924574007214|412|1
35.195689|19ad180e1eac3de8cd1f962a2f40e2f20ce49eb9|3.49|2014-09-14 16:08:00|1.4094857484078087|1|3800001611|412|0.6142806555579505|0|26|61|-80.826724|9|35.195689|RTE CEREAL ADULT|0.0|1|KELLOGG SPECIAL K 12 OZ BOX|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00038000016110|CEREAL|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|d8109d42e0c7a5bfbdcd64be016cb13550c2e252|14.49|2014-11-14 15:32:00|1.4094857484078087|1|3700088211|412|0.6142806555579505|1|26|426|-80.826724|72|35.195689|NFS-PAPER TOWELS|0.0|1|BOUNTY TOWEL 8 GIANT SAS|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00037000882114|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|fa04473b015991a22f016a5ca4461648f695e855|6.98|2014-11-10 12:49:00|1.4094857484078087|1|3800001611|412|0.6142806555579505|0|26|61|-80.826724|9|35.195689|RTE CEREAL ADULT|0.99|1|KELLOGG SPECIAL K 12 OZ BOX|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00038000016110|CEREAL|G1 GROCERY|-80.826724|1.4106924574007214|412|2
35.195689|9b88104901b18c6d8885f3b9d81c21e8e8cda263|14.49|2014-10-27 14:58:00|1.4094857484078087|1|3700088211|412|0.6142806555579505|1|26|426|-80.826724|72|35.195689|NFS-PAPER TOWELS|4.5|1|BOUNTY TOWEL 8 GIANT SAS|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00037000882114|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|840f2177903773d2425c8a7f8da73a91f2e32e98|4.5|2014-12-14 19:14:00|1.4094857484078087|1|1380017219|412|0.6142806555579505|0|26|1278|-80.826724|48|35.195689|SINGLE SERVE NUTRITIONAL|0.0|5|LC MACARONI CHEESE|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00013800188052|FROZEN MEALS|FROZEN|-80.826724|1.4106924574007214|412|2
35.195689|dbba42318d545494679b28db3faf29c925a758bb|6.79|2014-11-17 17:13:00|1.4094857484078087|1|2500005434|412|0.6142806555579505|0|26|335|-80.826724|56|35.195689|ORANGE JUICE-REGRIGERATED|0.8|3|SIMPLY ORANGE ORIGINAL|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00025000054334|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.826724|1.4106924574007214|412|1
35.195689|aaf7e08091d56488d47a40fcafc179baa8d9ab05|11.19|2014-12-08 15:25:00|1.4094857484078087|1|30041667803|412|0.6142806555579505|0|26|4062|-80.826724|1080|35.195689|TOOTH BRUSH-BATTERY|1.2|17|ORAL B PULSAR 40 SOFT TWIN PK|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00300416678030|ORAL HYGIENE|HBC|-80.826724|1.4106924574007214|412|1
35.195689|e9e635ef384920254945121241406cf00819d461|7.99|2014-11-16 09:56:00|1.4094857484078087|1|64786510001|412|0.6142806555579505|0|26|4195|-80.826724|1200|35.195689|COUGH & COLD REMEDY-ADULT|0.0|17|(FE)(JHK)AIRBORNE REG  ORANGE|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00647865100010|COUGH/COLD/SINUS|HBC|-80.826724|1.4106924574007214|412|1
35.195689|b1b49db586a5976095e9cdf51e5b408e3ffd36c0|7.98|2014-11-19 12:15:00|80.828402574597021|1|20405400000|412|35.2058053811622|0|8|504|-80.825175|64|35.152722|FRESH BERRIES|3.98|4|RED RASPBERRIES 6 OZ|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|35.209978091326001|00715756100019|FRESH PRODUCE|PRODUCE|-80.826724|80.826729446921846|160|2
35.195689|e1daaf362fc10da24007cdc05200291a7a982598|4.0|2015-02-14 08:32:00|80.828402574597021|1|84115200732|412|35.205805381648155|0|8|1165|-80.85013|87|35.175855|NFS-FRESH CONSUMER BUNCH|0.0|9|BUNCH- 3/$12 DAISY BUNCHES|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|35.209978091326001|00841152007321|FLORAL|FLORAL|-80.826724|80.826727865697862|218|1
35.195689|21999c68253820a65af67b0beee23fc71bef1052|3.58|2014-12-17 08:17:00|1.4094857484078087|1|5200033875|412|0.6142806555579505|0|26|171|-80.826724|20|35.195689|ISOTONIC DRINKS|0.9|1|GATORADE G2 GLACIER FREEZE|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00052000320152|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.826724|1.4106924574007214|412|2
35.195689|344f3e8c327660d0704e839050d0b00deb926e98|1.79|2014-12-22 21:45:00|1.4094857484078087|1|5200033875|412|0.6142806555579505|0|26|171|-80.826724|20|35.195689|ISOTONIC DRINKS|0.89|1|GATORADE G2 GLACIER FREEZE|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00052000320152|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|9e507595482f0f92472e8fe0ace44be2077e3ab0|3.58|2014-12-10 13:32:00|80.828402574597021|1|5200033875|412|35.205805381648155|0|8|171|-80.85013|20|35.175855|ISOTONIC DRINKS|0.89|1|GATORADE G2 GLACIER FREEZE|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|35.209978091326001|00052000320152|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.826724|80.826727865697862|218|2
35.195689|901131d680d6bed0ad67e41988007cc8c8d460bb|3.58|2014-12-12 10:59:00|80.828402574597021|1|5200033875|412|35.205805381648155|0|8|171|-80.85013|20|35.175855|ISOTONIC DRINKS|0.9|1|GATORADE G2 GLACIER FREEZE|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|35.209978091326001|00052000320152|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.826724|80.826727865697862|218|2
35.195689|7718125e6cea5ee837fcac9a2098a6d97f79881f|3.79|2015-02-14 17:08:00|1.4094857484078087|1|4950800600|412|0.6142806555579505|0|26|1981|-80.826724|480|35.195689|CHIPS|0.0|6|MINI CHEDDAR PRETZEL CRISPS|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00049508002178|DRY GOODS|DELI|-80.826724|1.4106924574007214|412|1
35.195689|dfeeaacb8fa86d068f921880c6988b1edff868e3|6.99|2015-02-19 16:36:00|1.4094857484078087|1|67729499901|412|0.6142806555579505|0|26|1220|-80.826724|275|35.195689|PASTA SC PREMIUM|2.0|1|MONTE BENE SC TOMATO BASIL|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00677294999022|PASTA SAUCES|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|b42eaa81415c90ed23d38e47f2bad03965f9675f|3.99|2015-02-22 17:52:00|1.4094857484078087|1|4157005982|412|0.6142806555579505|0|26|1148|-80.826724|21|35.195689|ALMONDS|0.0|1|BLUE DIAMOND ALM SALT/VINEGAR|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00041570053386|NUTS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|ec9fe4bf08746bd71c5b2c5131b5f699fdc4aa8a|2.69|2015-01-30 09:16:00|1.4094857484078087|1|5150020441|412|0.6142806555579505|0|26|103|-80.826724|15|35.195689|REMAINING FLOUR|0.0|1|PILLSBURY BEST FLOUR-UNBLEACHD|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00051500222416|FLOUR|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|c43b782a83ad374e4346eae26aaf1bd18bef9a3a|1.69|2014-09-28 12:49:00|1.4094857484078087|1|4900000044|412|0.6142806555579505|0|26|55|-80.826724|8|35.195689|REGULAR|0.0|23|CB COKE SINGLE 20 OZ.|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00049000000443|CARBONATED BEVERAGES|BEVERAGE|-80.826724|1.4106924574007214|412|1
35.195689|aae8fb81b1fe6b3c9d0c6f661dc24f09c59101bc|4.29|2014-12-06 17:54:00|1.4094857484078087|1|4900005235|412|0.6142806555579505|0|26|55|-80.826724|8|35.195689|REGULAR|0.79|23|SPRITE 7.5 OZ CAN|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00049000052374|CARBONATED BEVERAGES|BEVERAGE|-80.826724|1.4106924574007214|412|1
35.195689|6518ee6bd1799c07b70fe0fd85fb6404ea4d7614|4.49|2014-09-15 16:47:00|1.4094857484078087|1|2100000900|412|0.6142806555579505|0|26|317|-80.826724|52|35.195689|CHUNK AND BAR CHEESE|0.0|3|CRACKER BARREL EX SHARP CHED C|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00021000005239|CHEESE|DAIRY|-80.826724|1.4106924574007214|412|1
35.195689|f9a3bda61ce286f89f1de82e5acfa92dc167353a|3.49|2014-11-12 14:10:00|1.4094857484078087|1|7203695248|412|0.6142806555579505|0|26|1611|-80.826724|371|35.195689|PITA'S AND FLAT BREADS|0.0|14|FFM WHEAT PITA POCKET|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00072036952516|BREAD|BAKERY|-80.826724|1.4106924574007214|412|1
35.195689|625ef5dfeb981694c6d5cd19a85961e251c8a962|6.27|2015-02-21 18:27:00|1.4094857484078087|1|7203676359|412|0.6142806555579505|0|26|345|-80.826724|57|35.195689|ORGANIC MILK|0.0|3|HTO ORGANIC FF SKIM GAL|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00072036763624|MILK|DAIRY|-80.826724|1.4106924574007214|412|1
35.195689|40f9a636633130bc942fbc442be8ba0c8efda95e|2.99|2014-11-25 09:05:00|1.4094857484078087|1|7203698444|412|0.6142806555579505|0|26|266|-80.826724|307|35.195689|SHELLS AND PIE CRUSTS|0.99|5|HT PIE CRUSTS DEEP DISH|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00072036984449|DESSERTS FROZEN|FROZEN|-80.826724|1.4106924574007214|412|1
35.195689|3a8244974fc38fad588111d234eec3e83fe220cb|4.58|2015-01-29 10:10:00|1.4094857484078087|1|4800122129|412|0.6142806555579505|0|26|213|-80.826724|33|35.195689|SOUP MIXES|0.0|1|EKNORR SOUP MIX VEGETABLE|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00048001221291|SOUP|G1 GROCERY|-80.826724|1.4106924574007214|412|2
35.195689|bc1197ec479d0f111f6ae913b558df059e79186e|5.69|2014-09-20 08:08:00|1.4094857484078087|1|7756725423|412|0.6142806555579505|0|26|252|-80.826724|45|35.195689|PREMIUM ICE CREAM|2.85|5|BREYERS FRENCH VANILLA I/C|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00077567254382|ICE CREAM|FROZEN|-80.826724|1.4106924574007214|412|1
35.195689|1e87d988d562a864f6717516dcfd0de71f4b3f59|1.54|2015-03-02 16:19:00|1.4094857484078087|1|7203641991|412|0.6142806555579505|0|26|1212|-80.826724|272|35.195689|HISP BEANS/PEPPERS|0.0|1|HT BEANS REFRIED FAT FREE|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00072036419910|HISPANIC PREP. FOODS|G1 GROCERY|-80.826724|1.4106924574007214|412|2
35.195689|374a08e45a2855d3e3214764f52fc30d984fb97c|6.99|2014-10-01 16:49:00|1.4094857484078087|1|5161116589|412|0.6142806555579505|0|26|845|-80.826724|100|35.195689|NATURAL/ORGANIC BACON|0.0|19|COLEMAN UNCURED NATURAL BACON|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00051611165893|BACON|CASE READY MEATS|-80.826724|1.4106924574007214|412|1
35.195689|dff24a71954467e5787bb9fff1b09399dae4e511|6.99|2015-03-07 18:55:00|1.4094857484078087|1|5161116589|412|0.6142806555579505|0|26|845|-80.826724|100|35.195689|NATURAL/ORGANIC BACON|1.0|19|COLEMAN UNCURED NATURAL BACON|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00051611165893|BACON|CASE READY MEATS|-80.826724|1.4106924574007214|412|1
35.195689|64e1837cfefea20180b5018baf83e9faa6c9c24b|7.49|2014-09-12 13:39:00|80.828402574597021|1|4667716751|412|35.2058053811622|0|8|6153|-80.825175|1546|35.152722|BULB-REFLECTORS|0.0|18|PHILIPS 45W R30 I/D FLOOD|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|35.209978091326001|00046677167516|LIGHT BULBS/ELECTRICAL|GM|-80.826724|80.826729446921846|160|1
35.195689|638c2832ef969dc2340518a790a03b0203bb6973|9.19|2014-11-02 17:53:00|1.4094857484078087|1|90000035402|412|0.6142806555579505|0|26|427|-80.826724|72|35.195689|NFS-TOILET TISSUE|2.2|1|NORTHERN ULT SOFT/STRONG 12DR|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00042000963657|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|beb4548a349434c17a5342c9cbe761c9c930f6e2|9.98|2015-01-07 09:39:00|1.4094857484078087|1|71575620002|412|0.6142806555579505|0|26|504|-80.826724|64|35.195689|FRESH BERRIES|2.49|4|STRAWBERRIES 1LB CLAM|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00812049005102|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|2
35.195689|4a8dea5c816ea9166884eb737fa1d08723df3180|3.49|2014-11-03 18:53:00|1.4094857484078087|1|2500004786|412|0.6142806555579505|0|26|335|-80.826724|56|35.195689|ORANGE JUICE-REGRIGERATED|0.5|3|MINUTE MAID PULP FREE|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00025000047893|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.826724|1.4106924574007214|412|1
35.195689|c0e792793e0aae25a23ed302a084bac62378bf61|6.98|2015-01-10 08:34:00|1.4094857484078087|1|2500004786|412|0.6142806555579505|0|26|335|-80.826724|56|35.195689|ORANGE JUICE-REGRIGERATED|1.0|3|MINUTE MAID PULP FREE|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00025000047893|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.826724|1.4106924574007214|412|2
35.195689|2d70555c70a6e0a12dcb8409dcc4efe9564cf839|3.49|2014-09-22 10:06:00|1.4094857484078087|1|2500004786|412|0.6142806555579505|0|26|335|-80.826724|56|35.195689|ORANGE JUICE-REGRIGERATED|0.5|3|MINUTE MAID PULP FREE|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00025000047893|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.826724|1.4106924574007214|412|1
35.195689|49ac8b6b0afa1c50eb1da19d28eb01258915963a|28.56|2015-02-28 07:30:00|1.4094857484078087|1|20496000000|412|0.6142806555579505|0|26|755|-80.826724|87|35.195689|NFS-BALLOONS|0.0|9|*BALLOONS|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00204960000005|FLORAL|FLORAL|-80.826724|1.4106924574007214|412|1
35.195689|0d0e4d3722e06516f76396f5f786c92b26c5e292|14.28|2015-02-07 10:25:00|1.4094857484078087|1|20496000000|412|0.6142806555579505|0|26|755|-80.826724|87|35.195689|NFS-BALLOONS|0.0|9|*BALLOONS|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00204960000005|FLORAL|FLORAL|-80.826724|1.4106924574007214|412|1
35.195689|462d6a8d5a4b6b2666a977fc071bb95bcdda871b|7.14|2015-02-27 10:21:00|1.4094857484078087|1|20496000000|412|0.6142806555579505|0|26|755|-80.826724|87|35.195689|NFS-BALLOONS|0.0|9|*BALLOONS|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00204960000005|FLORAL|FLORAL|-80.826724|1.4106924574007214|412|1
35.195689|8d0a1ae97ffe769530cbbf4394d378ea1789e774|1.69|2014-12-21 16:10:00|1.4094857484078087|1|4600083251|412|0.6142806555579505|0|26|1212|-80.826724|272|35.195689|HISP BEANS/PEPPERS|0.0|1|OEP CHILIES GREEN CHOPPED|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00046000832517|HISPANIC PREP. FOODS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|1f06f0961c6887b9ef9f43cdd901b1b1bddf656c|4.99|2015-01-10 16:35:00|1.4094857484078087|1|7410880050|412|0.6142806555579505|0|26|3671|-80.826724|1060|35.195689|HAIR BRUSH|0.0|17|CONAIR PRO NYLON BRUSH|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00074108800527|HAIR CARE ACCESSORIES|HBC|-80.826724|1.4106924574007214|412|1
35.195689|784814f1891586f4dfdf1fa066b99805537534a9|2.99|2014-11-05 14:47:00|1.4094857484078087|1|7203698315|412|0.6142806555579505|0|26|425|-80.826724|72|35.195689|NFS-PAPER NAPKINS|0.99|1|YH ANTIBAC WIPES CITRUS SCENT|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00072036983145|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|902ffa5860d07c5721ef278545573f20af88c990|7.35|2015-01-13 18:52:00|1.4094857484078087|1|4470002268|412|0.6142806555579505|0|26|481|-80.826724|100|35.195689|CENTER CUT BACON|3.68|19|OSCAR MAYER CTR SLICED BACON|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00044700022689|BACON|CASE READY MEATS|-80.826724|1.4106924574007214|412|1
35.195689|a0558b65b2f0c6327914ddb9ac98aecf16617c71|0.69|2015-03-09 13:38:00|1.4094857484078087|1||412|0.6142806555579505|0|26|509|-80.826724|64|35.195689|FRESH CITRUS-REMAINING|0.09|4|LEMONS, LARGE|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00204053000004|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|1
35.195689|484d7c52ed7a4cef4d10342853f43cd6e4f6056b|1.67|2014-11-26 17:25:00|80.828402574597021|1|3120001605|412|35.205805382112153|0|8|106|-80.80146|16|35.17739|CRANBERRY SAUCE|0.17|1|OS CRANBERRY SC JELLIED|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|35.209978091326001|00031200016058|FRUIT-CAN/JAR|G1 GROCERY|-80.826724|80.826724940034225|208|1
35.195689|7278aec25ecf1184a94555261adf5934bb9c29b0|2.03|2014-10-21 19:40:00|1.4094857484078087|1||412|0.6142806555579505|0|26|528|-80.826724|64|35.195689|FRESH BROCCOLI|0.0|4|COO BROCCOLI CROWNS (RPC)|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00204549000006|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|1
35.195689|4b5f2e47f09f11e3c03106c15549be6cd900c11a|2.19|2015-02-10 16:22:00|1.4094857484078087|1|5150076040|412|0.6142806555579505|0|26|24|-80.826724|3|35.195689|FROSTING-READY-TO-SPREAD|0.4|1|PILLSBURY VANILLA FROSTING|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00051500760802|BAKING SUPPLIES|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|549524b95b292c07e8924e5ef9ef934188c917d4|2.79|2015-03-05 08:16:00|1.4094857484078087|1|5000069386|412|0.6142806555579505|0|26|341|-80.826724|57|35.195689|CREAMERS|0.45|3|COFFE-MATE NAT BLISS VANILLA|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00050000693863|MILK|DAIRY|-80.826724|1.4106924574007214|412|1
35.195689|3d7938ebed8ef3d149e4c11d662262d4e1b6918c|2.79|2015-02-24 09:30:00|1.4094857484078087|1|5000069386|412|0.6142806555579505|0|26|341|-80.826724|57|35.195689|CREAMERS|0.0|3|COFFE-MATE NAT BLISS VANILLA|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00050000693863|MILK|DAIRY|-80.826724|1.4106924574007214|412|1
35.195689|026715df80aae59b58253e7d71a8c789d64788f8|2.79|2015-02-20 09:11:00|1.4094857484078087|1|5000069386|412|0.6142806555579505|0|26|341|-80.826724|57|35.195689|CREAMERS|0.0|3|COFFE-MATE NAT BLISS VANILLA|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00050000693863|MILK|DAIRY|-80.826724|1.4106924574007214|412|1
35.195689|be0450fa97bb175fcdafcc4d9c982b3a03ccb46b|5.59|2014-10-22 14:50:00|1.4094857484078087|1|20631400000|412|0.6142806555579505|0|26|1825|-80.826724|410|35.195689|BH SALAMI|0.0|6|BOARS HEAD HARD SALAMI|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00206314000006|BH MEAT|DELI|-80.826724|1.4106924574007214|412|1
35.195689|07c1a1392a7699115beda8023a41e838e6c3f447|5.6|2014-10-13 19:04:00|1.4094857484078087|1|20598400000|412|0.6142806555579505|0|26|1822|-80.826724|410|35.195689|BH CHICKEN|1.27|6|BOARS HEAD EVERROAST CKN BRST|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00205984000002|BH MEAT|DELI|-80.826724|1.4106924574007214|412|1
35.195689|8c533c784e4d82e964a92abc1bba9f196e33c88d|2.79|2014-11-04 14:29:00|1.4094857484078087|1|4667716948|412|0.6142806555579505|0|26|6123|-80.826724|1546|35.195689|BULB-3 WAYS|0.0|18|PHILIPS 50/100W LONG LIFE 3 WA|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00046677169480|LIGHT BULBS/ELECTRICAL|GM|-80.826724|1.4106924574007214|412|1
35.195689|f61db944743b792abd0edbf5ffecc21fad5ba516|13.25|2015-03-08 19:07:00|1.4094857484078087|1|3700088211|412|0.6142806555579505|0|26|426|-80.826724|72|35.195689|NFS-PAPER TOWELS|1.26|1|BOUNTY TOWEL 8 GIANT WHITE|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00037000882138|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|83a4470428dd274024b4dbba9d3ee0c4b12d730b|2.11|2014-11-16 15:07:00|1.4094857484078087|1||412|0.6142806555579505|0|26|562|-80.826724|64|35.195689|FRESH CUT FRUIT|0.0|4|HONEYDEW CHUNKS (IN-STORE)|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00204343000004|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|1
35.195689|878d9f5a455820a9040ba09b5a5fe411e2137a4b|1.67|2015-02-12 12:41:00|1.4094857484078087|1|7203657050|412|0.6142806555579505|0|26|687|-80.826724|61|35.195689|BLENDED|0.0|3|HT VANILLA NONFAT YOGURT|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00072036570512|YOGURT|DAIRY|-80.826724|1.4106924574007214|412|1
35.195689|e93100ba8ced3759eadc2eb53689990a3ce7d650|1.69|2014-10-06 19:11:00|80.828402574597021|1|1700009270|412|35.205805381648155|0|8|722|-80.85013|73|35.175855|NFS-HAND SOAPS|0.0|1|DIAL LIQ GOLD HAND SOAP|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|35.209978091326001|00017000091532|PERSONAL SOAP/BATH ADDITIVES|G1 GROCERY|-80.826724|80.826727865697862|218|1
35.195689|944ea05b289947c53faaad4018042e6399369926|2.67|2015-02-28 19:59:00|1.4094857484078087|1|7064000461|412|0.6142806555579505|0|26|275|-80.826724|45|35.195689|SUPER PREMIUM ICE CREAM|0.0|5|B BUNNY PERSONALS COOKIE DOUGH|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00070640004645|ICE CREAM|FROZEN|-80.826724|1.4106924574007214|412|2
35.195689|f9261d515c649abaa1a33b7975a5b20ce347a8ec|3.58|2014-11-17 17:23:00|1.4094857484078087|1|5100001047|412|0.6142806555579505|0|26|212|-80.826724|33|35.195689|CONDENSED SOUP|0.54|1|CAMP COND LIGHT CHICKEN GUMBO|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00051000010810|SOUP|G1 GROCERY|-80.826724|1.4106924574007214|412|2
35.195689|9639263baea468bfa55ba36c4e3796f78f3511ce|3.38|2014-10-02 08:17:00|1.4094857484078087|1|5200033875|412|0.6142806555579505|0|26|171|-80.826724|20|35.195689|ISOTONIC DRINKS|0.44|1|GATORADE G2 FRUIT PUNCH|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00052000321982|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.826724|1.4106924574007214|412|2
35.195689|c9c3d996d3071a03bcde4ffb7eeb6a1b6fb9f380|1.69|2014-11-23 16:37:00|1.4094857484078087|1|7680828073|412|0.6142806555579505|0|26|149|-80.826724|23|35.195689|WHSE PASTA CORE|0.31|1|BARILLA PASTA MEDIUM SHELLS|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00076808517989|PASTA|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|16d044f8f8d8f2a21a17e8ba4ca122d7a235357a|7.16|2014-12-17 15:13:00|1.4094857484078087|1|5000001011|412|0.6142806555579505|0|26|145|-80.826724|22|35.195689|MILK-CANNED|1.82|1|CARNATION EVAPORATED MILK|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00050000010110|PACKAGED MILKS & MODIFIERS|G1 GROCERY|-80.826724|1.4106924574007214|412|4
35.195689|1c1c92c5133054062a5eb7d2e2604d98ee851e2a|0.75|2015-02-27 12:37:00|1.4094857484078087|1||412|0.6142806555579505|0|26|1635|-80.826724|375|35.195689|BULK (BAGELS)|0.25|14|BULK  BAGELS|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00072036955500|BAGELS|BAKERY|-80.826724|1.4106924574007214|412|1
35.195689|507b8137d334253bbeb8d2290b033827b3e097f3|3.0|2014-09-30 18:28:00|1.4094857484078087|1||412|0.6142806555579505|0|26|1635|-80.826724|375|35.195689|BULK (BAGELS)|0.0|14|BULK  BAGELS|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00072036955500|BAGELS|BAKERY|-80.826724|1.4106924574007214|412|4
35.195689|5c2d630f4916396ccddbfb4897a4a38263f1e8d8|3.0|2014-11-02 08:40:00|1.4094857484078087|1||412|0.6142806555579505|0|26|1635|-80.826724|375|35.195689|BULK (BAGELS)|0.0|14|BULK  BAGELS|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00072036955500|BAGELS|BAKERY|-80.826724|1.4106924574007214|412|4
35.195689|071651a58b4253d7cdec6eee7a48c504f68542d3|7.98|2014-09-11 19:30:00|80.828402574597021|1|71575620002|412|35.205805382112153|0|8|504|-80.80146|64|35.17739|FRESH BERRIES|0.98|4|STRAWBERRIES 1LB CLAM|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|35.209978091326001|00665290001184|FRESH PRODUCE|PRODUCE|-80.826724|80.826724940034225|208|2
35.195689|2e30d7dfd5b77b02254a63dc7ae380e58ae506a9|8.45|2014-11-15 15:37:00|1.4094857484078087|1|7800014645|412|0.6142806555579505|0|26|55|-80.826724|8|35.195689|REGULAR|2.2|23|CANADA DRY CLUB SODA 1 LTR|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00078000146455|CARBONATED BEVERAGES|BEVERAGE|-80.826724|1.4106924574007214|412|5
35.195689|ea1ec4b6748b86ca96cfc7aad6bfe7c2f058f7f9|4.45|2014-10-17 14:29:00|1.4094857484078087|1|7218063473|412|0.6142806555579505|0|26|254|-80.826724|892|35.195689|PREMIUM PIZZA|0.0|5|RED BARON PEPPERONI|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00072180634733|FROZEN PIZZA|FROZEN|-80.826724|1.4106924574007214|412|1
35.195689|95741cbc5f0524c9ee18ed37f25682daf883166c|3.69|2014-11-07 13:14:00|1.4094857484078087|1|7240071124|412|0.6142806555579505|0|26|25|-80.826724|3|35.195689|BAKING SYRUPS|0.7|1|GRANDMA'S ORIGINAL MOLASSES|11ed418aa421367a74da40d43a08fa23e3b83e91|0.6990175757768262|0.61471665291522548|00072400711244|BAKING SUPPLIES|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.03469|a7fb1158769d2a03b8d8bee995fbc1c8786af146|1.5|2014-09-16 19:49:00|80.970590786568081|1|7203663107|82|35.077344170799897|0|55|1262|-80.994596|57|35.061685|HALF N HALF WHIPPING CREAM|0.0|3|HT HALF & HALF|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00072036632036|MILK|DAIRY|-80.97058|80.970588998988319|475|1
35.03469|1279012ab1b16ce4343ab9fa50669474e22876ff|3.34|2014-11-18 19:22:00|80.970590786568081|1|7203670851|82|35.077344170799897|0|55|1262|-80.994596|57|35.061685|HALF N HALF WHIPPING CREAM|0.0|3|HIGHLAND CREST HALF&HALF|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00072036708519|MILK|DAIRY|-80.97058|80.970588998988319|475|2
35.03469|2a8ddbbebd454599f7d7ad9e1b2de305d1bd704c|1.67|2014-11-02 16:21:00|80.970590786568081|1|7203670851|82|35.077344170799897|0|55|1262|-80.994596|57|35.061685|HALF N HALF WHIPPING CREAM|0.0|3|HIGHLAND CREST HALF&HALF|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00072036708519|MILK|DAIRY|-80.97058|80.970588998988319|475|1
35.03469|944823d27e137ba8b2f1ec4bc58a77beecec746f|3.74|2014-12-22 19:39:00|80.970590786568081|1|7203670851|82|35.077344170799897|0|55|1262|-80.994596|57|35.061685|HALF N HALF WHIPPING CREAM|0.0|3|HIGHLAND CREST HALF&HALF|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00072036708519|MILK|DAIRY|-80.97058|80.970588998988319|475|2
35.03469|ea14451800b9ddef81a810c0bfaca57c2238eca1|1.87|2014-12-17 19:51:00|80.970590786568081|1|7203670851|82|35.077344170799897|0|55|1262|-80.994596|57|35.061685|HALF N HALF WHIPPING CREAM|0.0|3|HIGHLAND CREST HALF&HALF|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00072036708519|MILK|DAIRY|-80.97058|80.970588998988319|475|1
35.03469|8a5afdbf1e35984dc3ce6b1bc95ee1cef002ce65|6.68|2014-11-23 17:03:00|80.970590786568081|1|7203670851|82|35.077344170799897|0|55|1262|-80.994596|57|35.061685|HALF N HALF WHIPPING CREAM|0.0|3|HIGHLAND CREST HALF&HALF|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00072036708519|MILK|DAIRY|-80.97058|80.970588998988319|475|4
35.03469|59db5497b226a83a7da794d810904ffaf74763cb|1.67|2014-10-10 19:20:00|80.970590786568081|1|7203670851|82|35.077344170799897|0|55|1262|-80.994596|57|35.061685|HALF N HALF WHIPPING CREAM|0.0|3|HIGHLAND CREST HALF&HALF|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00072036708519|MILK|DAIRY|-80.97058|80.970588998988319|475|1
35.03469|28f9233338c946d27a4675d5e39adf180d016510|1.67|2014-10-26 19:06:00|80.970590786568081|1|7203670851|82|35.077344170799897|0|55|1262|-80.994596|57|35.061685|HALF N HALF WHIPPING CREAM|0.0|3|HIGHLAND CREST HALF&HALF|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00072036708519|MILK|DAIRY|-80.97058|80.970588998988319|475|1
35.03469|d90f031321d67e16744e910c1b2189e940c6600d|1.67|2014-09-12 19:17:00|80.970590786568081|1|7203670851|82|35.077344170799897|0|55|1262|-80.994596|57|35.061685|HALF N HALF WHIPPING CREAM|0.0|3|HIGHLAND CREST HALF&HALF|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00072036708519|MILK|DAIRY|-80.97058|80.970588998988319|475|1
35.03469|d2eafb43937e01d6a6bfa21627fc8366b6894fcb|3.74|2015-02-17 17:12:00|80.970590786568081|1|7203670851|82|35.077344170799897|0|55|1262|-80.994596|57|35.061685|HALF N HALF WHIPPING CREAM|0.0|3|HIGHLAND CREST HALF&HALF|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00072036708519|MILK|DAIRY|-80.97058|80.970588998988319|475|2
35.03469|20ff532194d87966f6326e8c709b51e22d3e7221|4.23|2015-01-27 18:47:00|1.4132775322775095|1||82|0.6114706929155321|0|58|529|-80.97058|64|35.03469|FRESH ASPARAGUS|0.21|4|GREEN  ASPARAGUS|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|0.61177642288969325|00204080000008|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|2d34c6978bbd76220c5565fb8618da1ab71405f3|4.89|2015-01-13 19:07:00|80.970590786568081|1||82|35.077344170799897|0|55|529|-80.994596|64|35.061685|FRESH ASPARAGUS|0.0|4|GREEN  ASPARAGUS|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00204080000008|FRESH PRODUCE|PRODUCE|-80.97058|80.970588998988319|475|1
35.03469|66ed3d592924d302e04f165ca64f0547ea54afed|8.53|2014-09-13 19:03:00|80.970590786568081|1||82|35.077344155951799|0|55|529|-81.027334|64|34.977331|FRESH ASPARAGUS|0.38|4|GREEN  ASPARAGUS|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00204080000008|FRESH PRODUCE|PRODUCE|-80.97058|80.970624398999078|149|1
35.03469|fdbe84cd34e17886cbaba641bb6ddf8ebc1c793c|3.67|2015-02-08 19:30:00|80.970590786568081|1||82|35.077344170799897|0|55|529|-80.994596|64|35.061685|FRESH ASPARAGUS|0.92|4|GREEN  ASPARAGUS|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00204080000008|FRESH PRODUCE|PRODUCE|-80.97058|80.970588998988319|475|1
35.03469|961566ecdcfdc501bb74aaad3bc939aa109e5b2e|8.78|2014-10-29 19:49:00|80.970590786568081|1||82|35.077344170799897|0|55|529|-80.994596|64|35.061685|FRESH ASPARAGUS|0.44|4|GREEN  ASPARAGUS|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00204080000008|FRESH PRODUCE|PRODUCE|-80.97058|80.970588998988319|475|1
35.03469|a21af8d94685a78545ebb300b62b63938fbd0507|10.58|2014-12-29 18:52:00|80.970590786568081|1||82|35.077344170799897|0|55|529|-80.994596|64|35.061685|FRESH ASPARAGUS|0.0|4|GREEN  ASPARAGUS|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00204080000008|FRESH PRODUCE|PRODUCE|-80.97058|80.970588998988319|475|1
35.03469|c0588705f1cf06db98693ff4c1b3ffbaf2f21ade|2.19|2015-02-14 18:43:00|80.970590786568081|1|4900005010|82|35.077344170799897|0|55|55|-80.994596|8|35.061685|REGULAR|0.2|23|SPRITE  2 LITER|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00049000050158|CARBONATED BEVERAGES|BEVERAGE|-80.97058|80.970588998988319|475|1
35.03469|4104774a28b1586ed529cc3e05376101b4845cbc|2.38|2014-10-30 21:58:00|80.970590786568081|1|3940001747|82|35.077344170799897|0|55|242|-80.994596|39|35.061685|CANNED BEANS|0.38|1|BUSH BEAN SND BLACK|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00039400018841|VEGETABLES-CAN/JAR|G1 GROCERY|-80.97058|80.970588998988319|475|2
35.03469|c9ab7165a2fd809867e4bec162bb5f40899c4a21|1.19|2014-12-23 21:20:00|80.970590786568081|1|3940001747|82|35.077344170799897|0|55|242|-80.994596|39|35.061685|CANNED BEANS|0.19|1|BUSH BEAN BLACK MILD CHILI SC|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00039400015024|VEGETABLES-CAN/JAR|G1 GROCERY|-80.97058|80.970588998988319|475|1
35.03469|47fd902a12b7f0c761dfddcdcc111e1292d747e2|3.99|2015-01-07 07:17:00|1.4132775322775095|1|4650075764|82|0.6114706929155321|0|58|393|-80.97058|68|35.03469|NFS-AIR FRESHENERS|1.49|1|GLADE WAX MELTS-LAV PCH BLOSSM|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|0.61177642288969325|00046500750946|FRESHENERS/DEODORIZERS|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|7f2b20e3c1161078138a0181940cde3bda79e291|3.29|2015-01-25 16:41:00|80.970590786568081|1|7203644036|82|35.077344170799897|0|55|273|-80.994596|43|35.061685|PREMIUM NOVELTIES|0.0|5|HT ICE CREAM SANDWICH-12PK|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00072036440365|FROZEN NOVELTIES|FROZEN|-80.97058|80.970588998988319|475|1
35.03469|b761bb928214af50e38d41d90d5961845c17da11|2.79|2014-11-02 16:31:00|80.970590786568081|1|7203698374|82|35.077344170799897|0|55|423|-80.994596|72|35.061685|NFS-DISPOSE PLATES/BOWLS|0.79|1|YH ULTRA DESIGNER BOWLS 20 OZ|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00072036983749|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.97058|80.970588998988319|475|1
35.03469|3ca0c9dfa3039dac738b4db8dcf92c4a6efd7746|9.29|2015-01-20 20:29:00|80.970590786568081|1|3160401285|82|35.077344158902214|0|55|4594|-80.8062|1215|35.037115|VITAMIN B|4.65|17|NM VITAMIN B6 100MG|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00031604012854|VITAMINS & SUPPLEMENTS|HBC|-80.97058|80.970619945703035|27|1
35.03469|73f2e974229d9781b8acc54fe48ae2eefb129345|3.99|2014-11-21 21:26:00|80.970590786568081|1|4400002854|82|35.077344163304957|0|55|1248|-80.992182|12|35.103409|SANDWICH COOKIES|0.49|1|OREO GOLDEN|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00044000032586|COOKIES|G1 GROCERY|-80.97058|80.97061217377869|88|1
35.03469|dea56113a59e9de231191b486a737008b474eeb6|1.99|2014-11-15 08:26:00|80.970590786568081|1|5100000524|82|35.077344170799897|0|55|1201|-80.994596|33|35.061685|RTS CANNED|0.49|1|CHUNKY POTATO CHEDDAR BACON|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00051000128041|SOUP|G1 GROCERY|-80.97058|80.970588998988319|475|1
35.03469|11b39a2bf15b9db0b741c6ef496aefd5582d909b|3.19|2014-12-01 17:33:00|80.970590786568081|1|5150005722|82|35.077344170799897|0|55|123|-80.994596|19|35.061685|JELLY/JAMS|1.19|1|SMUCKER'S STRAWBERRY SQUEEZE|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00051500057223|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.97058|80.970588998988319|475|1
35.03469|6e069924a94e4390c9ad5afc1b673ac28ca5de99|0.77|2014-09-28 16:01:00|80.970590786568081|1|7203610114|82|35.077344170799897|0|55|55|-80.994596|8|35.061685|REGULAR|0.0|23|HT CRANBERRY GINGER AL 2 LITER|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00072036983916|CARBONATED BEVERAGES|BEVERAGE|-80.97058|80.970588998988319|475|1
35.03469|c3f6f979db00b8eb7a4228a7c8fdfab7a7f14848|2.69|2014-10-04 17:20:00|80.970590786568081|1|7203698161|82|35.077344170799897|0|55|124|-80.994596|16|35.061685|APPLESAUCE MULTISERVE|0.0|1|HT APPLESAUCE (UNSWTND)|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00072036981622|FRUIT-CAN/JAR|G1 GROCERY|-80.97058|80.970588998988319|475|1
35.03469|3d426d423f731b5704cb01492c811db574847b30|2.39|2014-11-15 16:56:00|80.970590786568081|1|7203697771|82|35.077344170799897|0|55|239|-80.994596|38|35.061685|RICE-PACKAGED & BULK|0.0|1|HT RICE WHITE 80|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00072036977717|RICE GRAINS AND BEANS|G1 GROCERY|-80.97058|80.970588998988319|475|1
35.03469|25fd81e3ed4ba1cb7bcc46701dd840c0560e9a31|1.99|2014-11-13 19:17:00|80.970590786568081|1|7127915101|82|35.077344170799897|0|55|555|-80.994596|64|35.061685|PACKAGED SALADS|0.0|4|F.E. SHREDS|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00071279151014|FRESH PRODUCE|PRODUCE|-80.97058|80.970588998988319|475|1
35.03469|3e03f6132a5ac29058ac1d38d53d68b91b2ddad5|1.89|2014-11-04 22:27:00|80.970590786568081|1|31254662380|82|35.077344170799897|0|55|4207|-80.994596|1200|35.061685|COUGH DROP-ADULT|0.0|17|HALLS ICE BLUE 30'S  -62928|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00312546629288|COUGH/COLD/SINUS|HBC|-80.97058|80.970588998988319|475|1
35.03469|155a8775ea2dbf202db3ae4ffb40e9bf4e2f2ab9|1.89|2014-11-07 21:16:00|80.970590786568081|1|31254662380|82|35.077344155951799|0|55|4207|-81.027334|1200|34.977331|COUGH DROP-ADULT|0.7|17|HALLS ICE BLUE 30'S  -62928|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00312546629288|COUGH/COLD/SINUS|HBC|-80.97058|80.970624398999078|149|1
35.03469|30131cbb58b5bedda51e4a6f25f6dafcb8f57890|4.69|2014-12-14 12:46:00|80.970590786568081|1|4900002468|82|35.077344170799897|0|55|54|-80.994596|8|35.061685|DIET|4.69|23|DIET COKE .5 LITER/6 PK.|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.97058|80.970588998988319|475|1
35.03469|2efd5175081531d71eb93524c149dca41890f490|2.79|2014-10-25 10:46:00|80.970590786568081|1|5210000245|82|35.077344170799897|0|55|1246|-80.994596|34|35.061685|SPICE BLENDS|0.0|1|MC GRILL MATES MONTREAL CHICKN|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00052100002460|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.97058|80.970588998988319|475|1
35.03469|839021f9f1b106cf0d9eb5dc9a940a3966db3a63|5.99|2015-02-15 13:44:00|80.970590786568081|1|7756725423|82|35.077344170799897|0|55|252|-80.994596|45|35.061685|PREMIUM ICE CREAM|3.0|5|BREYERS EX CREAMY VANILLA|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00077567250049|ICE CREAM|FROZEN|-80.97058|80.970588998988319|475|1
35.03469|f8b8385d2b50050e029fc126fe79b064bb962ce6|2.78|2015-01-12 18:28:00|1.4132775322775095|1|3710003578|82|0.6114706929155321|0|58|245|-80.97058|39|35.03469|VEGETABLES-CORE|1.39|1|LIBBY CORN CREAM STYLE|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|0.61177642288969325|00037100036134|VEGETABLES-CAN/JAR|G1 GROCERY|-80.97058|1.4132032182494703|82|2
35.03469|13c07d551f19d9af4b2c4eb601ce3241e0a01ae9|9.89|2014-10-18 20:20:00|1.4132775322775095|1|7023011720|82|0.6114706929155321|0|58|730|-80.97058|24|35.03469|NFS-CAT LITTER|1.1|1|TIDY CAT IOC CAT LITTER 20 #JU|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|0.61177642288969325|00070230117205|PET FOOD/SUPPLIES|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|2dc7bd44effbf56e6e719c93c56d0859f04c335e|4.99|2015-01-13 22:29:00|80.970590786568081|1|4900002468|82|35.077344170799897|0|55|54|-80.994596|8|35.061685|DIET|4.99|23|COKE ZERO .5L 6PK PET|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00049000045840|CARBONATED BEVERAGES|BEVERAGE|-80.97058|80.970588998988319|475|1
35.03469|2a7ffd62cf425f3249beb2fe19273e144dacd18f|1.79|2015-01-22 08:41:00|80.970590786568081|1|5200033875|82|35.077344170799897|0|55|171|-80.994596|20|35.061685|ISOTONIC DRINKS|0.41|1|GATORADE AM TROPICAL MANGO|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00052000322132|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.97058|80.970588998988319|475|1
35.03469|d7637fe12357ab87aaccf0018c3b399880598480|7.98|2015-02-23 19:08:00|80.970590786568081|1|4470003050|82|35.077344170799897|0|55|840|-80.994596|102|35.061685|TUBS|0.98|19|OM DELI FRESH MESQUITE TURKEY|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00044700030707|LUNCHMEATS|CASE READY MEATS|-80.97058|80.970588998988319|475|2
35.03469|6afb1e4bf64ec8da2496f04e6a2507410e9b9898|1.25|2014-11-23 17:05:00|80.970590786568081|1|76866330908|82|35.077344170799897|0|55|8598|-80.994596|1792|35.061685|NEWSPAPERS|0.0|18|THE HERALD SUNDAY|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00768663309082|NEWSPAPERS|GM|-80.97058|80.970588998988319|475|1
35.03469|ba0a686638dd765f3292744883a1ccdd56bf944d|5.99|2014-11-27 11:58:00|80.970590786568081|1|1650053764|82|35.077344155951799|0|55|4236|-81.027334|1200|34.977331|DEX ADULT/CHILDREN|0.0|17|ALKA SELTZER PLUS COLD 50586|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00016500537649|COUGH/COLD/SINUS|HBC|-80.97058|80.970624398999078|149|1
35.03469|e5b3fa7955127067b365da1174f27c379d2513f3|7.78|2014-09-15 09:09:00|1.4132775322775095|1|2100060464|82|0.6114706929155321|0|58|315|-80.97058|52|35.03469|CHEESE-PROCESSED-SLICED|1.78|3|KRAFT SHARP CHEDDAR SINGLES|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|0.61177642288969325|00021000616480|CHEESE|DAIRY|-80.97058|1.4132032182494703|82|2
35.03469|f40793ed55bf6b92f074fcd4fbdde486a1c11694|3.85|2015-01-14 18:04:00|80.970590786568081|1|4812127620|82|35.077344170799897|0|55|1037|-80.994596|164|35.061685|ENGLISH MUFFINS|1.93|7|THOMAS SEASONAL EM PP|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00048121221003|BREAKFAST|COMMERCIAL BAKERY|-80.97058|80.970588998988319|475|1
35.03469|dca50ecba6efcc9e3379ef3b97b89ba2cdfb3f3f|2.85|2015-01-27 12:25:00|1.4132775322775095|1|4400000055|82|0.6114706929155321|0|58|88|-80.97058|13|35.03469|FLAKED SODA CRACKERS|0.35|1|NABISCO PREMIUMS|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|0.61177642288969325|00044000000578|CRACKERS|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|3f17534b8505f3109312babb513549a7fde313cb|1.39|2015-02-28 13:14:00|80.970590786568081|1|7203602056|82|35.077344170799897|0|55|78|-80.994596|11|35.061685|MUSTARD|0.7|1|HT MUSTARD YELLOW 14 OZ|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00072036020567|CONDIMENTS|G1 GROCERY|-80.97058|80.970588998988319|475|1
35.03469|3010f0fe3641f8e1ad645ab0b8f5a6068ce4db4c|7.92|2015-02-28 13:06:00|80.970590786568081|1|20496000000|82|35.077344170799897|0|55|755|-80.994596|87|35.061685|NFS-BALLOONS|0.0|9|*BALLOONS|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00204960000005|FLORAL|FLORAL|-80.97058|80.970588998988319|475|1
35.03469|c4484d0f1f945d431171ad5799ea40b42e304f1a|1.49|2015-01-23 21:59:00|80.970590786568081|1|4900005537|82|35.077344170799897|0|55|55|-80.994596|8|35.061685|REGULAR|0.49|23|DR PEPPER 1.25 LITER BOTTLE|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00078000082395|CARBONATED BEVERAGES|BEVERAGE|-80.97058|80.970588998988319|475|1
35.03469|0ff90bb091fafb4a0efe4734a1f37b3edc3dc5cd|6.79|2014-10-23 20:14:00|1.4132775322775095|1|1200080994|82|0.6114706929155321|0|58|55|-80.97058|8|35.03469|REGULAR|6.79|23|MTN DEW CODE RED FRIDGEMATE|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|0.61177642288969325|00012000809989|CARBONATED BEVERAGES|BEVERAGE|-80.97058|1.4132032182494703|82|1
35.03469|257e6e26182728ebff3fd01b05d51f4723a85422|5.69|2014-10-17 09:42:00|1.4132775322775095|1|5190001602|82|0.6114706929155321|0|58|839|-80.97058|102|35.03469|STACK PACKS|0.0|19|LOF PREMIUM BLACK FOREST HAM|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|0.61177642288969325|00051900016134|LUNCHMEATS|CASE READY MEATS|-80.97058|1.4132032182494703|82|1
35.03469|2c6492369b0ab3c6141fa6ac44643c74c2b7b948|2.19|2014-10-04 15:51:00|80.970590786568081|1|1200000496|82|35.077344170799897|0|55|54|-80.994596|8|35.061685|DIET|0.69|23|DIET PEPSI MAX 2LTR|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00012000018817|CARBONATED BEVERAGES|BEVERAGE|-80.97058|80.970588998988319|475|1
35.03469|114bc3d3233fb3b80f1122ddf87b95086faea0d1|5.37|2014-09-15 18:34:00|80.970590786568081|1|20165900000|82|35.077344170799897|0|55|297|-80.994596|49|35.061685|GROUND BEEF|1.54|2|GROUND BEEF 93% LEAN|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00201659000001|BEEF|MEAT|-80.97058|80.970588998988319|475|1
35.03469|c3d562232da783f43e470de7f5c161c98f80ff4e|1.69|2014-10-22 18:25:00|80.970590786568081|1|1200000129|82|35.077344170799897|0|55|54|-80.994596|8|35.061685|DIET|0.0|23|CB DIET PEPSI 20 OZ NR|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00012000001307|CARBONATED BEVERAGES|BEVERAGE|-80.97058|80.970588998988319|475|1
35.03469|93f08390ff3d3ee222a1d38fd5bb36a5d0c173f8|4.99|2014-09-11 19:44:00|80.970590786568081|1|2410044068|82|35.077344170799897|0|55|87|-80.994596|13|35.061685|CHEESE CRACKERS|1.49|1|CHEEZ-IT WHITE CHEDDAR|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00024100789382|CRACKERS|G1 GROCERY|-80.97058|80.970588998988319|475|1
35.03469|9edbd9d632800e7c817073f78b4926236a1e938d|29.99|2014-12-24 17:54:00|80.970590786568081|1|20310600000|82|35.077344170799897|0|55|1153|-80.994596|87|35.061685|NFS-FRESH CUT ARRANGE|0.0|9|*FOAM ARRANGEMENTS|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00203106000008|FLORAL|FLORAL|-80.97058|80.970588998988319|475|1
35.03469|8f8ccf813443558cbe069a3bdeb352a17fc90e39|5.13|2014-11-21 19:47:00|80.970590786568081|1||82|35.077344170799897|0|55|529|-80.994596|64|35.061685|FRESH ASPARAGUS|0.0|4|GREEN  ASPARAGUS|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00204080000008|FRESH PRODUCE|PRODUCE|-80.97058|80.970588998988319|475|1
35.03469|8dc95ed8b8557b707c98a360c884c2b4feaf9012|4.0|2014-10-19 16:43:00|80.970590786568081|1||82|35.077344170799897|0|55|511|-80.994596|64|35.061685|FRESH AVOCADOS|0.21|4|AVOCADOS, HASS XL 36CT|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00204770000004|FRESH PRODUCE|PRODUCE|-80.97058|80.970588998988319|475|2
35.03469|22c85488b12b303fc059d0b47a8cebf79dc40275|3.49|2014-11-07 08:53:00|80.970590786568081|1|20496400000|82|35.077344170799897|0|55|756|-80.994596|87|35.061685|NFS-FLORAL ACCESSORIES|0.0|9|*ACCESSORIES|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00204964000001|FLORAL|FLORAL|-80.97058|80.970588998988319|475|1
35.03469|2d1b8ee4aee6cb5613402b0a2c0328e868ce69ac|2.0|2014-09-21 08:12:00|80.970590786568081|1|7203663118|82|35.077344170799897|0|55|1262|-80.994596|57|35.061685|HALF N HALF WHIPPING CREAM|0.0|3|HT HALF & HALF|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00072036632043|MILK|DAIRY|-80.97058|80.970588998988319|475|1
35.03469|b33427f8aa7d709eb21003de382b94b877587b74|2.19|2014-10-14 20:07:00|80.970590786568081|1|1200000496|82|35.077344170799897|0|55|54|-80.994596|8|35.061685|DIET|0.2|23|DIET PEPSI 2 LTR NR|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00012000002311|CARBONATED BEVERAGES|BEVERAGE|-80.97058|80.970588998988319|475|1
35.03469|3d563f56fb2fe5ce379922be0ed040b393474435|4.38|2014-12-13 18:59:00|80.970590786568081|1|1200000496|82|35.077344170799897|0|55|54|-80.994596|8|35.061685|DIET|0.4|23|DIET PEPSI 2 LTR NR|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00012000002311|CARBONATED BEVERAGES|BEVERAGE|-80.97058|80.970588998988319|475|2
35.03469|94f4e5c1657cb459c7e6b8d4f9a83f0b34e42546|2.19|2015-02-22 13:15:00|80.970590786568081|1|1200000496|82|35.077344170799897|0|55|54|-80.994596|8|35.061685|DIET|0.2|23|DIET PEPSI 2 LTR NR|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00012000002311|CARBONATED BEVERAGES|BEVERAGE|-80.97058|80.970588998988319|475|1
35.03469|bcff5bcd2d34e0690486d49d28436ee5e0a29037|13.9|2015-02-28 13:14:00|80.970590786568081|1|76211104952|82|35.077344170799897|0|55|1600|-80.994596|370|35.061685|PACKAGED FOOD|3.92|22|CHOC HEARTS|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00762111049520|STARBUCKS|COFFEE SHOP|-80.97058|80.970588998988319|475|2
35.03469|b06d3e0b76e98064ec829d2d451fd5a9f1fea22c|1.37|2015-01-31 18:29:00|80.970590786568081|1|7203690020|82|35.077344170799897|0|55|1034|-80.994596|163|35.061685|HOT DOG|0.0|7|H T HOT DOG BUNS|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00072036900203|BUNS/ROLLS|COMMERCIAL BAKERY|-80.97058|80.970588998988319|475|1
35.03469|3f86284276db8e328c2fcc29c344989583884b68|8.0|2014-10-12 20:53:00|80.970590786568081|1|89307700194|82|35.077344170799897|0|55|1165|-80.994596|87|35.061685|NFS-FRESH CONSUMER BUNCH|0.0|9|BUNCHES - ASST. LILY BUNCHES|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00893077001946|FLORAL|FLORAL|-80.97058|80.970588998988319|475|2
35.03469|953de28858c60fe329d40a151718fc5b6118f31c|13.58|2014-11-04 13:51:00|80.970590786568081|1|1200080994|82|35.077344167697291|0|55|55|-80.837892|8|34.937113|REGULAR|3.4|23|DR. PEPPER FRIDGEMATE|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00078000082166|CARBONATED BEVERAGES|BEVERAGE|-80.97058|80.97060181673956|372|2
35.03469|f4ae99675db8c8d6d2dfc0b5a9db4d3839635039|1.99|2014-09-28 16:03:00|80.970590786568081|1|7203648011|82|35.077344170799897|0|55|274|-80.994596|44|35.061685|ICE|0.0|5|HT BAGGED ICE 10LB (456)|128891d5c73515994509aa846993ae2cf8cc4b64|2.947300240091429|35.077427448337218|00000000004560|ICE|FROZEN|-80.97058|80.970588998988319|475|1
35.4437|3e5e1b793df01c96b1e5e66b1cc2fdaf048ceb70|4.9|2014-12-10 20:09:00|1.4102725052409182|3|1450000253|272|0.6186092640891142|0|1|1272|-80.8955|50|35.4437|BAG VEG STEAM|0.9|5|BE STEAMFRESH PREM GRN BEANS|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00014500011572|VEGETABLES-FROZEN|FROZEN|-80.8955|1.4118928250470728|272|2
35.4437|10114800955ba0931be59c2e07d713f177506acc|4.9|2014-11-30 18:02:00|1.4102725052409182|3|1450000253|272|0.6186092640891142|0|1|1272|-80.8955|50|35.4437|BAG VEG STEAM|1.22|5|BE STEAMFRESH PREM GRN BEANS|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00014500011572|VEGETABLES-FROZEN|FROZEN|-80.8955|1.4118928250470728|272|2
35.4437|98344e7577a1fb141b0c5a00b66760de426c0f29|2.69|2015-02-10 14:48:00|80.89430079996653|3|1450000253|272|35.456943265423064|0|32|1272|-80.861571|50|35.444615|BAG VEG STEAM|1.35|5|BE STEAMFRESH PREM GRN BEANS|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00014500011572|VEGETABLES-FROZEN|FROZEN|-80.8955|80.895502661736458|340|1
35.4437|e8e6efacafc539a0c4f203b856ec70d3bc170545|4.9|2014-10-03 16:37:00|80.89430079996653|3|1450000253|272|35.456943251192634|0|32|1272|-80.945176|50|35.323246|BAG VEG STEAM|0.9|5|BE STEAMFRESH PREM GRN BEANS|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00014500011572|VEGETABLES-FROZEN|FROZEN|-80.8955|80.895523980537376|166|2
35.4437|ff1977c27aa44cb90117518abef4a79d1afaa6a9|4.9|2014-09-16 22:39:00|1.4102725052409182|3|1450000253|272|0.6186092640891142|0|1|1272|-80.8955|50|35.4437|BAG VEG STEAM|1.23|5|BE STEAMFRESH PREM GRN BEANS|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00014500011572|VEGETABLES-FROZEN|FROZEN|-80.8955|1.4118928250470728|272|2
35.4437|c343f8325000f03ad3434adff2c5ec7a3e5e8367|4.9|2014-12-19 06:16:00|80.89430079996653|3|1450000253|272|35.456943265332697|0|32|1272|-80.86175|50|35.40953|BAG VEG STEAM|1.23|5|BE STEAMFRESH PREM GRN BEANS|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00014500011572|VEGETABLES-FROZEN|FROZEN|-80.8955|80.895503269802148|209|2
35.4437|13a0264ffa939dce5200544e39489e4dae5efd27|4.9|2014-09-13 16:19:00|1.4102725052409182|3|1450000253|272|0.6186092640891142|0|1|1272|-80.8955|50|35.4437|BAG VEG STEAM|1.22|5|BE STEAMFRESH PREM GRN BEANS|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00014500011572|VEGETABLES-FROZEN|FROZEN|-80.8955|1.4118928250470728|272|2
35.4437|7d697ce11ee9a8b1904a56d63ebf409370da7d43|4.9|2014-12-02 20:33:00|1.4102725052409182|3|1450000253|272|0.6186092640891142|0|1|1272|-80.8955|50|35.4437|BAG VEG STEAM|1.22|5|BE STEAMFRESH PREM GRN BEANS|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00014500011572|VEGETABLES-FROZEN|FROZEN|-80.8955|1.4118928250470728|272|2
35.4437|3b7ab63d6995782829da5190bb365771c27ccb8e|4.9|2014-09-27 11:43:00|80.89430079996653|3|1450000253|272|35.456943265423064|0|32|1272|-80.861571|50|35.444615|BAG VEG STEAM|0.9|5|BE STEAMFRESH PREM GRN BEANS|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00014500011572|VEGETABLES-FROZEN|FROZEN|-80.8955|80.895502661736458|340|2
35.4437|3cba22a73ea79e864648cd8c737f340231359117|4.9|2015-01-30 16:00:00|80.89430079996653|3|1450000253|272|35.456943264724117|0|32|1272|-80.893784|50|35.478031|BAG VEG STEAM|0.9|5|BE STEAMFRESH PREM GRN BEANS|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00014500011572|VEGETABLES-FROZEN|FROZEN|-80.8955|80.895505914557205|179|2
35.4437|33081523a5fa90b3021312707f2eead034c08898|4.9|2014-10-24 21:28:00|1.4102725052409182|3|1450000253|272|0.6186092640891142|0|1|1272|-80.8955|50|35.4437|BAG VEG STEAM|0.9|5|BE STEAMFRESH PREM GRN BEANS|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00014500011572|VEGETABLES-FROZEN|FROZEN|-80.8955|1.4118928250470728|272|2
35.4437|36968638338b60db5c727641e33f05b5b4c070d7|3.69|2015-02-03 17:13:00|80.89430079996653|3|2500005542|272|35.456943264724117|0|32|335|-80.893784|56|35.478031|ORANGE JUICE-REGRIGERATED|0.69|3|SIMPLY ORANGE ORIGINAL|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00025000055423|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.8955|80.895505914557205|179|1
35.4437|932b78388abfac7257f1d4f32d29608e62d3f030|7.91|2015-02-05 22:01:00|1.4102725052409182|3|20869700000|272|0.6186092640891142|0|1|648|-80.8955|154|35.4437|FISH FLTS/STK FARM RAISD|0.99|12|TEQUILA LIME CATFISH FILLETS|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00208697000000|FISH FILLETS/STEAKS|SEAFOOD|-80.8955|1.4118928250470728|272|1
35.4437|2f60a4ff35740c365897f749a589951a27193599|1.0|2015-01-02 15:33:00|80.89430079996653|3|5360000178|272|35.456943264724117|0|32|687|-80.893784|61|35.478031|BLENDED|0.2|3|LA CHOCOLAT MINT YOGURT|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00053600001793|YOGURT|DAIRY|-80.8955|80.895505914557205|179|1
35.4437|e44f0e49b47df2856352c876722e9848eac68335|4.39|2014-10-17 17:12:00|80.89430079996653|3|5480001008|272|35.456943265332697|0|32|239|-80.86175|38|35.40953|RICE-PACKAGED & BULK|1.2|1|UNCLE BENS RICE CONVERTED 32|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00054800010080|RICE GRAINS AND BEANS|G1 GROCERY|-80.8955|80.895503269802148|209|1
35.4437|e5c41a2bf03b377cf41b29108c54589af8c5f653|1.55|2015-01-18 17:10:00|80.89430079996653|3|68954408205|272|35.456943264724117|0|32|685|-80.893784|61|35.478031|GREEK|0.55|3|FAGE 0% FRUYO PEACH GREEK YOG|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00689544082040|YOGURT|DAIRY|-80.8955|80.895505914557205|179|1
35.4437|24309dc36b714fa74f6e72213b0e803cde6aafdb|3.39|2015-01-25 18:11:00|80.89430079996653|3|2529300098|272|35.456943240683792|0|32|1263|-80.810056|57|35.219587|GOOD FOR YOU MILK|0.39|3|SILK PURE CASHEW MILK|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00025293002746|MILK|DAIRY|-80.8955|80.895531535804167|401|1
35.4437|b30f1f4749d483d3ec7082fb340f36979c1b7b4a|71.96|2015-01-03 16:29:00|80.89430079996653|3|7203678085|272|35.45694326165696|0|32|665|-80.814133|145|35.333742|PACKAGED RAW|17.99|12|FISHERMANS SHRIMP 21/30 EZP WH|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00072036780850|SHRIMP|SEAFOOD|-80.8955|80.895512545992858|472|2
35.4437|2819f63bc72c61f401d9ba7b331ae87fda2116c6|23.96|2015-01-06 18:38:00|80.89430079996653|3|20931700000|272|35.456943264724117|0|32|676|-80.893784|148|35.478031|TAILS|0.0|12|WC LOBSTER TAILS 4.2 OZ  (CA)|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00209317000004|LOBSTERS|SEAFOOD|-80.8955|80.895505914557205|179|1
35.4437|f0929e1e9ca09e9bca52efc2b455da5a870c716e|3.29|2014-11-18 20:19:00|80.89430079996653|3|7225091171|272|35.456943265423064|0|32|1033|-80.861571|163|35.444615|HAMBURGER|0.0|7|NATOWN WHITEWHEAT HAMS|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00072250911719|BUNS/ROLLS|COMMERCIAL BAKERY|-80.8955|80.895502661736458|340|1
35.4437|f2398d6199d0b5bf01fda1fb0c0513436012414e|3.29|2015-01-15 20:42:00|1.4102725052409182|3|7225091171|272|0.6186092640891142|0|1|1033|-80.8955|163|35.4437|HAMBURGER|0.0|7|NATOWN WHITEWHEAT HAMS|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00072250911719|BUNS/ROLLS|COMMERCIAL BAKERY|-80.8955|1.4118928250470728|272|1
35.4437|ab66ae32c4bd0520dd92bb183afb8ac6d161e972|3.29|2014-11-11 22:36:00|80.89430079996653|3|7225091171|272|35.456943264724117|0|32|1033|-80.893784|163|35.478031|HAMBURGER|0.0|7|NATOWN WHITEWHEAT HAMS|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00072250911719|BUNS/ROLLS|COMMERCIAL BAKERY|-80.8955|80.895505914557205|179|1
35.4437|8b1cd5d5614c63848d0b00b9fc2327fe279e6d63|1.2|2014-11-02 18:53:00|80.89430079996653|3|7047000100|272|35.456943264724117|0|32|687|-80.893784|61|35.478031|BLENDED|0.0|3|YOPLAIT ORIG  STRAWBERRY/BANA|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00070470003139|YOGURT|DAIRY|-80.8955|80.895505914557205|179|2
35.4437|317bea9460665cb1c03c9ca6ef4f453db428b571|2.4|2014-11-18 19:37:00|80.89430079996653|3|7047000100|272|35.456943265423064|0|32|687|-80.861571|61|35.444615|BLENDED|0.4|3|YOPLAIT ORG. FRENCH VANILLA|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00070470003238|YOGURT|DAIRY|-80.8955|80.895502661736458|340|4
35.4437|9bce73e59d0b043bdf26c89dab87f6df3a2fa487|1.2|2014-12-23 10:12:00|80.89430079996653|3|7047000100|272|35.456943265423064|0|32|687|-80.861571|61|35.444615|BLENDED|0.0|3|YOPLAIT ORIG  STRAWBERRY/BANA|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00070470003139|YOGURT|DAIRY|-80.8955|80.895502661736458|340|2
35.4437|1523d0b9ad5ea4f361e9ff2bdb40dcce1c311751|0.8|2014-10-11 11:31:00|80.89430079996653|3|7047000100|272|35.456943265423064|0|32|687|-80.861571|61|35.444615|BLENDED|0.3|3|YOPLAIT ORIG  STRAWBERRY/BANA|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00070470003139|YOGURT|DAIRY|-80.8955|80.895502661736458|340|1
35.4437|7d93b1bd53ab5f5f24167cc570bc2347dd41e44e|1.6|2014-10-14 22:57:00|80.89430079996653|3|7047000100|272|35.456943265423064|0|32|687|-80.861571|61|35.444615|BLENDED|0.6|3|YOPLAIT ORIG  STRAWBERRY/BANA|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00070470003139|YOGURT|DAIRY|-80.8955|80.895502661736458|340|2
35.4437|bff2feab38e19298d3f4083bdea5cdbd9a89b405|1.2|2015-02-23 23:05:00|80.89430079996653|3|7047000100|272|35.456943265423064|0|32|687|-80.861571|61|35.444615|BLENDED|0.2|3|YOPLAIT ORIG  STRAWBERRY/BANA|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00070470003139|YOGURT|DAIRY|-80.8955|80.895502661736458|340|2
35.4437|48cb949302fb4ad73b3136692bacf220d98eee0b|2.4|2014-12-28 16:10:00|1.4102725052409182|3|7047000100|272|0.6186092640891142|0|1|687|-80.8955|61|35.4437|BLENDED|0.0|3|YOPLAIT ORG. FRENCH VANILLA|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00070470003238|YOGURT|DAIRY|-80.8955|1.4118928250470728|272|4
35.4437|2333c13a3e780d34ab4be1f74d3fe846090804ae|1.8|2015-03-09 19:47:00|1.4102725052409182|3|7047000100|272|0.6186092640891142|0|1|687|-80.8955|61|35.4437|BLENDED|0.0|3|YOPLAIT ORG. FRENCH VANILLA|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00070470003238|YOGURT|DAIRY|-80.8955|1.4118928250470728|272|3
35.4437|05b52bee2d48a656962c0a85d8d6b172e5ae88df|1.7999999999999998|2015-01-20 20:38:00|80.89430079996653|3|7047000100|272|35.456943264724117|0|32|687|-80.893784|61|35.478031|BLENDED|0.30000000000000004|3|YOPLAIT ORG. FRENCH VANILLA|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00070470003238|YOGURT|DAIRY|-80.8955|80.895505914557205|179|3
35.4437|82027c7ac5889904bec674b326cdcc091e5cd514|2.45|2015-01-20 19:44:00|80.89430079996653|3|1450000253|272|35.456943265423064|0|32|1272|-80.861571|50|35.444615|BAG VEG STEAM|0.45|5|BE STEAMFRESH PEAS&MUSHROOMS|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00014500011619|VEGETABLES-FROZEN|FROZEN|-80.8955|80.895502661736458|340|1
35.4437|a29cf42707a2fe5ae4b49818f53e55fc418250e6|2.45|2014-09-23 20:50:00|1.4102725052409182|3|1450000253|272|0.6186092640891142|0|1|1272|-80.8955|50|35.4437|BAG VEG STEAM|0.45|5|BE STEAMFRESH PEAS&MUSHROOMS|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00014500011619|VEGETABLES-FROZEN|FROZEN|-80.8955|1.4118928250470728|272|1
35.4437|d523a7c795a3e425c834eb27678ba567bcc5aeaa|3.99|2014-12-02 20:20:00|80.89430079996653|3|7203663995|272|35.456943264724117|0|32|342|-80.893784|57|35.478031|FRESH MILK|1.52|3|HARRIS TEETER 1% MILK|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00072036631275|MILK|DAIRY|-80.8955|80.895505914557205|179|1
35.4437|335d9dca5420a210f2f8b0cf430c47f5c8348ced|3.49|2015-02-08 16:03:00|1.4102725052409182|3|7203663995|272|0.6186092640891142|0|1|342|-80.8955|57|35.4437|FRESH MILK|0.72|3|HARRIS TEETER 1% MILK|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00072036631275|MILK|DAIRY|-80.8955|1.4118928250470728|272|1
35.4437|6584bf39829b76b7efb8755b0a2f8f0591bc03cc|3.65|2015-01-24 20:23:00|1.4102725052409182|3|4400002827|272|0.6186092640891142|0|1|1251|-80.8955|12|35.4437|WHOLESOME COOKIES|0.65|1|BELVITA BREAKFAST BITES CHOCOL|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00044000033323|COOKIES|G1 GROCERY|-80.8955|1.4118928250470728|272|1
35.4437|68a0c0912acd20641c75425c222d0d0965c0c257|2.85|2015-03-07 19:01:00|80.89430079996653|3|4400000055|272|35.456943264724117|0|32|88|-80.893784|13|35.478031|FLAKED SODA CRACKERS|0.35|1|NABISCO PREMIUM UNSALTED|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00044000000554|CRACKERS|G1 GROCERY|-80.8955|80.895505914557205|179|1
35.4437|ac2d0e63aed7f4471371de8c1adaba705d99a926|2.52|2014-09-26 19:06:00|80.89430079996653|3|20540400000|272|35.456943265423064|0|32|1832|-80.861571|415|35.444615|BH SLICING CHEESE|0.0|6|BOARS HEAD HORSERADISH CHEDDAR|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00205404000001|SLICING CHEESE|DELI|-80.8955|80.895502661736458|340|1
35.4437|9900d3c247525a27f0416f477782b0af4dc1c68d|7.139999999999999|2015-01-24 17:58:00|1.4102725052409182|3|3940001747|272|0.6186092640891142|0|1|242|-80.8955|39|35.4437|CANNED BEANS|1.14|1|BUSH BEAN SND BLACK|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00039400018841|VEGETABLES-CAN/JAR|G1 GROCERY|-80.8955|1.4118928250470728|272|6
35.4437|e8a97ef2585dcdf6d428064cd72bbcc92740c2e2|2.69|2015-02-15 18:34:00|1.4102725052409182|3|1450000253|272|0.6186092640891142|0|1|1272|-80.8955|50|35.4437|BAG VEG STEAM|0.69|5|BE STEAMFRESH ITALIAN BLEND|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00014500012913|VEGETABLES-FROZEN|FROZEN|-80.8955|1.4118928250470728|272|1
35.4437|d3ef4ff23334ed16c0b7b6f307b17daf9e45908a|2.45|2015-01-04 18:14:00|1.4102725052409182|3|1450000253|272|0.6186092640891142|0|1|1272|-80.8955|50|35.4437|BAG VEG STEAM|0.78|5|BE STEAMFRESH ITALIAN BLEND|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00014500012913|VEGETABLES-FROZEN|FROZEN|-80.8955|1.4118928250470728|272|1
35.4437|87ae2cc989b6f52004f35906d67a232a0b4d15ac|2.45|2014-10-06 19:46:00|1.4102725052409182|3|1450000253|272|0.6186092640891142|0|1|1272|-80.8955|50|35.4437|BAG VEG STEAM|0.45|5|BE STEAMFRESH ITALIAN BLEND|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00014500012913|VEGETABLES-FROZEN|FROZEN|-80.8955|1.4118928250470728|272|1
35.4437|cd648a9a229b8ddadcab960cf242a0f86828010e|2.29|2014-12-15 12:16:00|1.4102725052409182|3|7800023046|272|0.6186092640891142|0|1|55|-80.8955|8|35.4437|REGULAR|1.29|23|CANADA DRY GINGER ALE NR 2LTR|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00078000152463|CARBONATED BEVERAGES|BEVERAGE|-80.8955|1.4118928250470728|272|1
35.4437|011973ca4d9788d8c9c4bc0bebfe78616cd54fd0|2.02|2015-01-26 20:21:00|1.4102725052409182|3||272|0.6186092640891142|0|1|502|-80.8955|64|35.4437|FRESH BANANAS|0.0|4|BANANAS, YELLOW|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.8955|1.4118928250470728|272|1
35.4437|15c0ae9389ab3847552c4b1a28401f9e3d4ac415|6.98|2014-10-20 09:49:00|1.4102725052409182|3|3000001190|272|0.6186092640891142|0|1|60|-80.8955|9|35.4437|HOT CEREAL|1.98|1|QUAKER OATML RAISIN SPICE|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00030000013205|CEREAL|G1 GROCERY|-80.8955|1.4118928250470728|272|2
35.4437|d36d6e9d9de7e82db6886acb12d30c0aa6266f5c|2.59|2014-09-30 20:04:00|80.89430079996653|3|7047041381|272|35.456943264724117|0|32|687|-80.893784|61|35.478031|BLENDED|0.92|3|YOPLAIT FRENCH VANILLA 4PK|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00070470434810|YOGURT|DAIRY|-80.8955|80.895505914557205|179|1
35.4437|b9346572f88331162f35c88da2aa91c26acfc6bb|7.77|2014-09-30 20:17:00|1.4102725052409182|3|7047041381|272|0.6186092640891142|0|1|687|-80.8955|61|35.4437|BLENDED|2.77|3|YOPLAIT FRENCH VANILLA 4PK|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00070470434810|YOGURT|DAIRY|-80.8955|1.4118928250470728|272|3
35.4437|488630426fca5a2693c86bc149b3fde21174143f|5.85|2015-01-20 20:21:00|1.4102725052409182|3|1450001098|272|0.6186092640891142|0|1|1272|-80.8955|50|35.4437|BAG VEG STEAM|1.85|5|BE STEAMFRESH SWEET PEAS|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00014500011008|VEGETABLES-FROZEN|FROZEN|-80.8955|1.4118928250470728|272|3
35.4437|432ecf6d9eea3a00fd375663da92f2ff67624428|2.29|2015-01-06 19:32:00|80.89430079996653|3|7203663996|272|35.456943265423064|0|32|342|-80.861571|57|35.444615|FRESH MILK|0.82|3|HARRIS TEETER 1%  MILK|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00072036631305|MILK|DAIRY|-80.8955|80.895502661736458|340|1
35.4437|d73d9b11443ea9957b10e2bea561fca1911ff740|2.0|2015-03-02 12:17:00|1.4102725052409182|3|5100000524|272|0.6186092640891142|0|1|1201|-80.8955|33|35.4437|RTS CANNED|0.5|1|CHUNKY HR OLD FASH VEG BEEF|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00051000167767|SOUP|G1 GROCERY|-80.8955|1.4118928250470728|272|1
35.4437|8a104d43b7eadc576d6ea7288fbd0023c6c61e2f|3.79|2015-01-27 19:01:00|80.89430079996653|3|4850002013|272|35.456943263286576|0|32|335|-80.762919|56|35.442529|ORANGE JUICE-REGRIGERATED|1.29|3|TROPICANA PP ORIGINAL|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00048500301029|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.8955|80.895509610344121|471|1
35.4437|366e3fb695e754e9443ed866e640851d5224f3b0|11.879999999999999|2015-01-30 16:16:00|1.4102725052409182|3|20822400000|272|0.6186092640891142|0|1|669|-80.8955|146|35.4437|CRAB VALUE ADDED|1.19|12|CRAB STUFFED FLOUNDER|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00208224000008|CRAB|SEAFOOD|-80.8955|1.4118928250470728|272|2
35.4437|575ed3d10a50a22f3069dca5f3a3e7ae01292030|1.99|2014-10-30 17:43:00|80.89430079996653|3|7127900105|272|35.456943251192634|0|32|555|-80.945176|64|35.323246|PACKAGED SALADS|0.0|4|F.E. COLE SLAW 16OZ|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00071279123004|FRESH PRODUCE|PRODUCE|-80.8955|80.895523980537376|166|1
35.4437|7dfc35cab86dedeb251b05b016be086b8e00beea|1.99|2014-11-20 19:36:00|80.89430079996653|3|7127900105|272|35.456943263286576|0|32|555|-80.762919|64|35.442529|PACKAGED SALADS|0.0|4|F.E. COLE SLAW 16OZ|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00071279123004|FRESH PRODUCE|PRODUCE|-80.8955|80.895509610344121|471|1
35.4437|78a0b08e465c47cb532de3d957985cd4e52132ce|1.99|2015-02-13 18:54:00|80.89430079996653|3|7127900105|272|35.456943265332697|0|32|555|-80.86175|64|35.40953|PACKAGED SALADS|0.0|4|F.E. COLE SLAW 16OZ|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00071279123004|FRESH PRODUCE|PRODUCE|-80.8955|80.895503269802148|209|1
35.4437|1d58d67c51fcbd7b026edcb6be661106484af867|1.99|2014-09-26 18:59:00|1.4102725052409182|3|7127900105|272|0.6186092640891142|0|1|555|-80.8955|64|35.4437|PACKAGED SALADS|0.0|4|F.E. COLE SLAW 16OZ|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00071279123004|FRESH PRODUCE|PRODUCE|-80.8955|1.4118928250470728|272|1
35.4437|41d00937caf3971b14a5a21863f981727cee5f1c|6.5|2014-09-16 22:54:00|80.89430079996653|3|1380016610|272|35.456943265423064|0|32|1278|-80.861571|48|35.444615|SINGLE SERVE NUTRITIONAL|2.5|5|LC STEAK TIPS PORTABELLO|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00013800156501|FROZEN MEALS|FROZEN|-80.8955|80.895502661736458|340|2
35.4437|5a1e9a4d4988c99d8b5b1f083dc7710daafce06d|1.76|2015-01-05 13:05:00|80.89430079996653|3||272|35.456943264724117|0|32|502|-80.893784|64|35.478031|FRESH BANANAS|0.0|4|BANANAS, YELLOW|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00204011000008|FRESH PRODUCE|PRODUCE|-80.8955|80.895505914557205|179|1
35.4437|3c27f61c98e1cdc629005e8819582644138215c6|1.33|2014-11-28 22:06:00|80.89430079996653|3||272|35.456943265423064|0|32|502|-80.861571|64|35.444615|FRESH BANANAS|0.0|4|BANANAS, YELLOW|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00204011000008|FRESH PRODUCE|PRODUCE|-80.8955|80.895502661736458|340|1
35.4437|332acc7ccb25f3f5226bc8c5af92d452c6f1ea4d|1.05|2014-12-07 20:56:00|1.4102725052409182|3||272|0.6186092640891142|0|1|502|-80.8955|64|35.4437|FRESH BANANAS|0.0|4|BANANAS, YELLOW|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.8955|1.4118928250470728|272|1
35.4437|9ad4d701dff7cfdbf3060697b52d7edcf246c839|19.45|2014-10-15 19:34:00|1.4102725052409182|3|4400002827|272|0.6186092640891142|0|1|1251|-80.8955|12|35.4437|WHOLESOME COOKIES|4.45|1|BELVITA BREAKFAST CHOCOLATE|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00044000031947|COOKIES|G1 GROCERY|-80.8955|1.4118928250470728|272|5
35.4437|33bb15d2a39ab1a5cd7bb0704c3724b1ca4ab577|1.27|2014-11-12 19:03:00|1.4102725052409182|3|7203628032|272|0.6186092640891142|0|1|163|-80.8955|25|35.4437|RELISHES|0.0|1|HT RELISH SWEET 16|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|0.61833652052202714|00072036280329|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.8955|1.4118928250470728|272|1
35.4437|e82366ab21e5cc83791474c4439e7b6b55049a2b|1.32|2015-03-02 19:25:00|80.89430079996653|3||272|35.456943265423064|0|32|524|-80.861571|64|35.444615|FRESH PROD FRESH ONIONS|0.22|4|COO RED ONIONS|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00204082000006|FRESH PRODUCE|PRODUCE|-80.8955|80.895502661736458|340|1
35.4437|dc5e2db9fe385463514a222f5c6b1f46348c3c4c|2.4|2014-12-24 13:37:00|80.89430079996653|3|7047000100|272|35.456943264724117|0|32|687|-80.893784|61|35.478031|BLENDED|0.0|3|YOPLAIT ORG MIXED BERRY|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00070470003108|YOGURT|DAIRY|-80.8955|80.895505914557205|179|4
35.4437|bbd7624d4887314c2f269b7dda06f75b0f55134a|1.5|2014-11-20 19:39:00|80.89430079996653|3|81204900640|272|35.456943263286576|0|32|504|-80.762919|64|35.442529|FRESH BERRIES|0.0|4|BLUEBERRIES 6 OZ|134d5adaaf94c7021091dcb5e1489541e193618f|0.9150776716574354|35.45572462568753|00033383222288|FRESH PRODUCE|PRODUCE|-80.8955|80.895509610344121|471|1
35.478031|75204f2f638fe573183897101624f167c7b11689|1.55|2014-12-19 11:22:00|80.8939826282094|1|2920000307|179|35.485912169994826|0|2|149|-80.861571|23|35.444615|WHSE PASTA CORE|0.0|1|MUELLER PENNE RIGATE BOX|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00029200003079|PASTA|G1 GROCERY|-80.893784|80.893785936476448|340|1
35.478031|f88d4bb1a1d6b0d454a1332387d0123ad83a6ef9|3.79|2015-02-01 12:54:00|1.4102725052409182|1|2100062503|179|0.6192084530746164|0|1|318|-80.893784|52|35.478031|SHREDDED/GRATED CHEESE|1.89|3|KRAFT FINELY SHREDDED SHARP C|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00021000638741|CHEESE|DAIRY|-80.893784|1.4118628751971085|179|1
35.478031|9ceefabffbdb5d337abba20de2047c1a6018f781|7.79|2014-11-06 18:21:00|80.8939826282094|1|2279691005|179|35.485912169631028|0|2|3533|-80.8955|1045|35.4437|SHAMPOO-NATURAL|1.8|17|ORGANIX TEATREE MINT SHAMPOO|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00022796910141|HAIR & SCALP CARE|HBC|-80.893784|80.89378752106721|272|1
35.478031|1b8cf5b1463ace40060c56766d21dc98cccda648|8.33|2014-10-03 08:22:00|80.8939826282094|1|20249700000|179|35.485912168894963|0|2|297|-80.86175|49|35.40953|GROUND BEEF|0.42|2|NY STRIP STEAKBURGER 80% LEAN|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00202497000000|BEEF|MEAT|-80.893784|80.893789467652809|209|1
35.478031|af23418addf605299a9e5bbcb991f9674f2a7554|6.15|2014-11-13 13:37:00|1.4102725052409182|1|20337400000|179|0.6192084530746164|0|1|641|-80.893784|137|35.478031|PREMIUM PORK|0.0|2|PORK LOIN BNLS BUTTERFLY CHOPS|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00203382000006|PORK|MEAT|-80.893784|1.4118628751971085|179|1
35.478031|719aa5e634f29702e811de70ad723923d6ba771f|4.0|2015-02-25 12:38:00|80.8939826282094|1||179|35.485912169631028|0|2|531|-80.8955|64|35.4437|FRESH CORN|0.0|4|COO YELLOW CORN|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00204078000003|FRESH PRODUCE|PRODUCE|-80.893784|80.89378752106721|272|5
35.478031|97e1d5aee5ecfbf266a2a2d935b7b65affc8a8fe|6.99|2015-01-21 16:44:00|1.4102725052409182|1|8346724624|179|0.6192084530746164|0|1|4913|-80.893784|1240|35.478031|WART REMOVERS|0.0|17|WARTSTICK WART REMOVER|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00083467246242|FOOT CARE|HBC|-80.893784|1.4118628751971085|179|1
35.478031|1f8333725e3184fec4558bf902b24f2e567313a3|4.01|2015-02-05 10:21:00|80.8939826282094|1|20337400000|179|35.485912169631028|0|2|641|-80.8955|137|35.4437|PREMIUM PORK|0.0|2|PORK LOIN BNLS BUTTERFLY CHOPS|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00203382000006|PORK|MEAT|-80.893784|80.89378752106721|272|1
35.478031|661f1455381d2605a565cfdfb5ec91b6379cef07|5.99|2015-02-21 22:01:00|80.8939826282094|1|7756725423|179|35.485912169631028|0|2|252|-80.8955|45|35.4437|PREMIUM ICE CREAM|1.41|5|BREYERS S&D NSA BUTTER PECAN|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00077567281968|ICE CREAM|FROZEN|-80.893784|80.89378752106721|272|1
35.478031|b5c25614eca7f65e8e10ecccd235d175009a1e95|2.29|2015-01-31 13:46:00|1.4102725052409182|1|7800023046|179|0.6192084530746164|0|1|54|-80.893784|8|35.478031|DIET|0.79|23|CANADA DRY DT G/ALE 2 LITER|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00078000148466|CARBONATED BEVERAGES|BEVERAGE|-80.893784|1.4118628751971085|179|1
35.478031|069873a75d915a3bd8be9e446d96ca02d8c091db|2.99|2014-12-31 15:37:00|1.4102725052409182|1|7482064552|179|0.6192084530746164|0|1|6785|-80.893784|1568|35.478031|MAGAZINES WEEKLY|0.0|18|IN TOUCH WEEKLY|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00074820645529|MAGAZINES|GM|-80.893784|1.4118628751971085|179|1
35.478031|7274ed0a5eacf1e79124f4a47086f8ea3913f560|2.29|2014-12-17 10:48:00|1.4102725052409182|1|7800023046|179|0.6192084530746164|0|1|54|-80.893784|8|35.478031|DIET|1.29|23|CANADA DRY DT G/ALE 2 LITER|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00078000148466|CARBONATED BEVERAGES|BEVERAGE|-80.893784|1.4118628751971085|179|1
35.478031|0062a1360b4c21a755e4dcb19fa4c8f67e2ab93a|2.29|2014-12-06 21:16:00|1.4102725052409182|1|7800023046|179|0.6192084530746164|0|1|54|-80.893784|8|35.478031|DIET|1.29|23|CANADA DRY DT G/ALE 2 LITER|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00078000148466|CARBONATED BEVERAGES|BEVERAGE|-80.893784|1.4118628751971085|179|1
35.478031|7b51b225ec4c54da99e95cc2d60c6db6fdc75d3f|7.15|2015-02-26 15:26:00|80.8939826282094|1|4470003128|179|35.485912169631028|0|2|840|-80.8955|102|35.4437|TUBS|1.16|19|OM 1LB HONEY SMOKED TURKEY|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00044700058640|LUNCHMEATS|CASE READY MEATS|-80.893784|80.89378752106721|272|1
35.478031|66a127cc111fb7714253d53dcce97a56e256f204|2.99|2015-01-22 13:35:00|1.4102725052409182|1|4411544801|179|0.6192084530746164|0|1|1878|-80.893784|435|35.478031|HUMMUS|0.0|6|ORIGINAL ORGANIC HOMMUS|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00044115448012|SALADS|DELI|-80.893784|1.4118628751971085|179|1
35.478031|70b0a400106b144d041cd7f478e4439cad23dc6e|7.15|2014-10-31 12:05:00|1.4102725052409182|1|4470003128|179|0.6192084530746164|0|1|840|-80.893784|102|35.478031|TUBS|0.66|19|OM 1LB HONEY SMOKED TURKEY|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00044700058640|LUNCHMEATS|CASE READY MEATS|-80.893784|1.4118628751971085|179|1
35.478031|47f088675e615269e95391bd02070f806702410d|7.15|2015-02-09 11:28:00|80.8939826282094|1|4470003128|179|35.485912169631028|0|2|840|-80.8955|102|35.4437|TUBS|0.0|19|OM 1LB HONEY SMOKED TURKEY|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00044700058640|LUNCHMEATS|CASE READY MEATS|-80.893784|80.89378752106721|272|1
35.478031|514e8f2de9d50ea468176f9b24d900a081437d9b|2.99|2014-10-07 13:47:00|1.4102725052409182|1|4411544801|179|0.6192084530746164|0|1|1878|-80.893784|435|35.478031|HUMMUS|0.0|6|ORIGINAL ORGANIC HOMMUS|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00044115448012|SALADS|DELI|-80.893784|1.4118628751971085|179|1
35.478031|7d8b2eb7c11b43a943de8bad88c77bb067f3ae00|2.98|2014-10-13 13:25:00|80.8939826282094|1|5000000457|179|35.485912169631028|0|2|168|-80.8955|24|35.4437|NFS-CAT TREATS|0.0|1|FF APPETIZER WHT MEAT CHICKEN|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00050000004591|PET FOOD/SUPPLIES|G1 GROCERY|-80.893784|80.89378752106721|272|2
35.478031|8c94bc3f94b8c5c07724ab5cda678c43ba45954e|2.98|2014-12-05 13:09:00|80.8939826282094|1|5000000457|179|35.485912169631028|0|2|168|-80.8955|24|35.4437|NFS-CAT TREATS|0.48|1|FF APPETIZER WHT MEAT CHICKEN|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00050000004591|PET FOOD/SUPPLIES|G1 GROCERY|-80.893784|80.89378752106721|272|2
35.478031|7d6f29ac479aeb7c7e2181dd202b42c8546dd04b|5.96|2014-10-23 14:23:00|80.8939826282094|1|5000000457|179|35.485912169631028|0|2|168|-80.8955|24|35.4437|NFS-CAT TREATS|0.0|1|FF APPETIZER WHT MEAT CHICKEN|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00050000004591|PET FOOD/SUPPLIES|G1 GROCERY|-80.893784|80.89378752106721|272|4
35.478031|460730abd993e55f7e41b1d8e0ebbbda2897786e|4.47|2014-12-26 19:31:00|1.4102725052409182|1|5000000457|179|0.6192084530746164|0|1|168|-80.893784|24|35.478031|NFS-CAT TREATS|0.24|1|FF APPETIZER WHT MEAT CHICKEN|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00050000004591|PET FOOD/SUPPLIES|G1 GROCERY|-80.893784|1.4118628751971085|179|3
35.478031|0a6cdd2e32ecdd4b7fcabbf479e80516f0e4c56e|11.92|2014-10-08 11:12:00|80.8939826282094|1|5000000457|179|35.485912169631028|0|2|168|-80.8955|24|35.4437|NFS-CAT TREATS|0.0|1|FF APPETIZER WHT MEAT CHICKEN|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00050000004591|PET FOOD/SUPPLIES|G1 GROCERY|-80.893784|80.89378752106721|272|8
35.478031|ab5d2029a3fa08713b4f8a19746734b11c45e7ab|5.96|2015-01-10 16:01:00|80.8939826282094|1|5000000457|179|35.485912169631028|0|2|168|-80.8955|24|35.4437|NFS-CAT TREATS|0.0|1|FF APPETIZER WHT MEAT CHICKEN|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00050000004591|PET FOOD/SUPPLIES|G1 GROCERY|-80.893784|80.89378752106721|272|4
35.478031|446512848b3e86a159347b46a2684ac02b825267|4.47|2015-02-14 16:31:00|80.8939826282094|1|5000000457|179|35.485912169631028|0|2|168|-80.8955|24|35.4437|NFS-CAT TREATS|0.72|1|FF APPETIZER WHT MEAT CHICKEN|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00050000004591|PET FOOD/SUPPLIES|G1 GROCERY|-80.893784|80.89378752106721|272|3
35.478031|3d5d0b8754168830e0aece5753de53e7cce5552e|6.58|2015-01-25 16:38:00|80.8939826282094|1|5410000400|179|35.485912169631028|0|2|162|-80.8955|25|35.4437|PICKLES|1.65|1|VLASIC WHL KOSHER BABY DILL|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00054100004000|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.893784|80.89378752106721|272|2
35.478031|5b51c670755d6a3ff5d923b45cdedb94e174bf73|6.99|2014-11-26 11:04:00|80.8939826282094|1|7050106095|179|35.485912169631028|0|2|3249|-80.8955|1020|35.4437|FACIAL CLEANSER|0.0|17|(E)NEUTRO DP CLN GENTLE SCRB|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00070501050354|FACIAL CLEANSER & MOISTURIZER|HBC|-80.893784|80.89378752106721|272|1
35.478031|99eca4e1d4bcfd75f6849d7acc1033862be5b4ef|1.89|2014-12-31 10:15:00|1.4102725052409182|1|7069002210|179|0.6192084530746164|0|1|757|-80.893784|3|35.478031|BAKING NUTS|0.0|1|FISHER ALMONDS SLIVERED|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00070690022101|BAKING SUPPLIES|G1 GROCERY|-80.893784|1.4118628751971085|179|1
35.478031|c883aa9d7a6c88fcffcb8fd16d9bb8e617b4e2ac|3.99|2014-11-04 12:15:00|80.8939826282094|1|7056097799|179|35.485912169994826|0|2|1272|-80.861571|50|35.444615|BAG VEG STEAM|0.0|5|PCTSWT STM DLX ASPARAGUS SPEAR|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00070560977999|VEGETABLES-FROZEN|FROZEN|-80.893784|80.893785936476448|340|1
35.478031|4e181d54c79f99a25928cdc97dc48d1c9b4490d1|3.99|2015-01-29 10:38:00|1.4102725052409182|1|7203602701|179|0.6192084530746164|0|1|1878|-80.893784|435|35.478031|HUMMUS|0.5|6|FFM ARTISAN SMK PAPRIKA HUMMUS|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00072036027061|SALADS|DELI|-80.893784|1.4118628751971085|179|1
35.478031|7c574957b9a17b14e16ca5fb26cb1c24d7760bc9|3.99|2015-01-03 18:30:00|1.4102725052409182|1|7203602701|179|0.6192084530746164|0|1|1878|-80.893784|435|35.478031|HUMMUS|0.5|6|FFM ARTISAN SMK PAPRIKA HUMMUS|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00072036027061|SALADS|DELI|-80.893784|1.4118628751971085|179|1
35.478031|2ad5a4a4a2747ed7e20a682a76850999bf65357a|7.98|2014-10-27 12:42:00|80.8939826282094|1|7056097799|179|35.485912169631028|0|2|1272|-80.8955|50|35.4437|BAG VEG STEAM|1.98|5|PCTSWT STM DLX ASPARAGUS SPEAR|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00070560977999|VEGETABLES-FROZEN|FROZEN|-80.893784|80.89378752106721|272|2
35.478031|76aaee5636b46e018505f8e4d8e1b33ef258773c|3.99|2014-12-17 21:48:00|1.4102725052409182|1|7203602701|179|0.6192084530746164|0|1|1878|-80.893784|435|35.478031|HUMMUS|0.5|6|FFM ARTISAN SMK PAPRIKA HUMMUS|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00072036027061|SALADS|DELI|-80.893784|1.4118628751971085|179|1
35.478031|9ca70fe6e533396de786465ee37e2101cf53b6d3|3.99|2015-03-08 11:33:00|1.4102725052409182|1|7203602701|179|0.6192084530746164|0|1|1878|-80.893784|435|35.478031|HUMMUS|0.3|6|FFM ARTISAN SMK PAPRIKA HUMMUS|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00072036027061|SALADS|DELI|-80.893784|1.4118628751971085|179|1
35.478031|46f5e6e8c71b6533d5d15e4cd0e7027362d61af2|3.79|2014-11-02 16:48:00|80.8939826282094|1|5210000698|179|35.485912169631028|0|2|1245|-80.8955|34|35.4437|SINGLE SPICES|0.0|1|MC BAY LEAVES|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00052100006987|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.893784|80.89378752106721|272|1
35.478031|26ccb3f0182f68257d198ec9c4b70c3c8315bb6f|2.52|2015-02-22 12:49:00|80.8939826282094|1||179|35.485912169631028|0|2|522|-80.8955|64|35.4437|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00204664000004|FRESH PRODUCE|PRODUCE|-80.893784|80.89378752106721|272|1
35.478031|a863963f8eb593eda9c14463543370b0e31d16fc|2.29|2014-11-22 12:05:00|1.4102725052409182|1||179|0.6192084530746164|0|1|522|-80.893784|64|35.478031|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00204664000004|FRESH PRODUCE|PRODUCE|-80.893784|1.4118628751971085|179|1
35.478031|b534c02b55615bd172228002452bfa6e195b89fb|2.28|2015-01-04 16:13:00|1.4102725052409182|1||179|0.6192084530746164|0|1|522|-80.893784|64|35.478031|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00204664000004|FRESH PRODUCE|PRODUCE|-80.893784|1.4118628751971085|179|1
35.478031|65dab11dcb1871a5374eaaaf516f3eb32c8336ba|2.07|2015-01-29 11:53:00|80.8939826282094|1||179|35.485912169994826|0|2|522|-80.861571|64|35.444615|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00204664000004|FRESH PRODUCE|PRODUCE|-80.893784|80.893785936476448|340|1
35.478031|0c028db2f88e725f6d82a9ae84a6cc3941d806eb|7.0|2015-01-27 16:26:00|80.8939826282094|1|20943300000|179|35.485912169631028|0|2|664|-80.8955|145|35.4437|SHRIMP WILD CAUGHT|2.01|12|WC P & D ARGENTINA PINK SHRMP|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00209433000001|SHRIMP|SEAFOOD|-80.893784|80.89378752106721|272|1
35.478031|175c3c0e042f6d63e257cb3bc4243ffbf690453a|1.69|2014-10-28 13:40:00|1.4102725052409182|1|7203688003|179|0.6192084530746164|0|1|527|-80.893784|64|35.478031|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00072036880031|FRESH PRODUCE|PRODUCE|-80.893784|1.4118628751971085|179|1
35.478031|9b48c4f4291e775b39cc29b5433c939be7a175ca|3.38|2014-12-24 08:49:00|1.4102725052409182|1|7203688003|179|0.6192084530746164|0|1|527|-80.893784|64|35.478031|FRESH CARROTS|0.38|4|HT BABY CARROTS 1LB BAG|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00072036880031|FRESH PRODUCE|PRODUCE|-80.893784|1.4118628751971085|179|2
35.478031|ba1e2f1dc44a1b87d96dbff548eb9dfbfd8edacc|12.99|2015-02-14 10:48:00|1.4102725052409182|1|7203695587|179|0.6192084530746164|0|1|1707|-80.893784|387|35.478031|MESSAGE|3.0|14|12 INCH MESSAGE COOKIE|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00072036955876|COOKIES|BAKERY|-80.893784|1.4118628751971085|179|1
35.478031|4d97b4ce09d4851df2caaa6c2dadcbed4abf74c4|5.25|2014-10-30 14:29:00|80.8939826282094|1|7203633086|179|35.485912169631028|0|2|1148|-80.8955|21|35.4437|ALMONDS|0.4|1|HT ROASTED ALMONDS LIGHT SALT|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00072036979537|NUTS|G1 GROCERY|-80.893784|80.89378752106721|272|1
35.478031|3688c6644490719a8b20ab9f40bcb648acd303be|4.19|2014-10-05 09:12:00|80.8939826282094|1|4812127620|179|35.485912169631028|0|2|1037|-80.8955|164|35.4437|ENGLISH MUFFINS|0.0|7|THOMAS LITE MULTIGRAIN EM PP|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00048121276201|BREAKFAST|COMMERCIAL BAKERY|-80.893784|80.89378752106721|272|1
35.478031|95a09ee6a04f0b2d4a7cd78f8d873ac3c83a5bbe|3.99|2014-12-10 20:11:00|1.4102725052409182|1|4450097650|179|0.6192084530746164|0|1|840|-80.893784|102|35.478031|TUBS|0.0|19|HF THIN LS O/R TURKEY BREAST|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00044500976441|LUNCHMEATS|CASE READY MEATS|-80.893784|1.4118628751971085|179|1
35.478031|b6eb639164157416845f3f2c800c6a3d7898938d|3.95|2014-12-02 15:01:00|1.4102725052409182|1|4450097650|179|0.6192084530746164|0|1|840|-80.893784|102|35.478031|TUBS|0.0|19|HF THIN LS O/R TURKEY BREAST|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00044500976441|LUNCHMEATS|CASE READY MEATS|-80.893784|1.4118628751971085|179|1
35.478031|7bb427f6ea630e62b2cb68c0a03e85e6285b8a67|3.75|2014-11-11 14:35:00|80.8939826282094|1|4139000107|179|35.485912169994826|0|2|79|-80.861571|273|35.444615|ASIAN SAUCES/SEASONINGS|0.0|1|KIKKOMAN SOY SAUCE LT 15|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00041390001079|ASIAN PREP. FOODS|G1 GROCERY|-80.893784|80.893785936476448|340|1
35.478031|7a0882dd7e3d8b00eca94cb7d14ec210a95c18e3|3.99|2015-01-15 18:59:00|1.4102725052409182|1|4450097650|179|0.6192084530746164|0|1|840|-80.893784|102|35.478031|TUBS|0.65|19|HF THIN LS O/R TURKEY BREAST|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00044500976441|LUNCHMEATS|CASE READY MEATS|-80.893784|1.4118628751971085|179|1
35.478031|a96aa8f2e36103123b55fcb28bf2eb5176bcaa41|3.25|2015-03-03 13:49:00|80.8939826282094|1|1980020133|179|35.485912169631028|0|2|405|-80.8955|69|35.4437|NFS-WINDOW CLEANERS|0.0|1|WINDEX TRIGGER BLUE|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00019800201333|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.893784|80.89378752106721|272|1
35.478031|0d3dfba4dbfad26600d8ad10bc0d523e7e4e5617|2.79|2015-03-05 10:49:00|80.8939826282094|1|4133500053|179|35.485912169631028|0|2|184|-80.8955|28|35.4437|SALAD DRESSINGS-LIQUID|0.0|1|KENS DRS LT HONEY MUSTARD|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00041335335177|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.893784|80.89378752106721|272|1
35.478031|d028e9219da8b33d20676c6518b84e7d26f17077|3.49|2014-12-10 11:24:00|1.4102725052409182|1|5150004042|179|0.6192084530746164|0|1|126|-80.893784|19|35.478031|PRESERVES/MARMALADE|0.0|1|SMUCKERS S/F RED RASPBERRY|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00051500040010|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.893784|1.4118628751971085|179|1
35.478031|fd07bb609cefb9c6cfd43a0ab466ea86566c1961|2.29|2015-01-07 16:12:00|1.4102725052409182|1|7203663996|179|0.6192084530746164|1|1|342|-80.893784|57|35.478031|FRESH MILK|0.23|3|HARRIS TEETER FF SKIM MILK|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00072036631299|MILK|DAIRY|-80.893784|1.4118628751971085|179|1
35.478031|6e92f730b530d55ba7c5c67c1baaa18704790d4d|2.29|2015-01-19 19:03:00|1.4102725052409182|1|7203663996|179|0.6192084530746164|0|1|342|-80.893784|57|35.478031|FRESH MILK|0.23|3|HARRIS TEETER FF SKIM MILK|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00072036631299|MILK|DAIRY|-80.893784|1.4118628751971085|179|1
35.478031|b2bf65a0e19c62dedc89140f28d9042b38df30e3|3.99|2015-02-23 17:09:00|80.8939826282094|1|7203678108|179|35.485912169631028|0|2|670|-80.8955|146|35.4437|CRAB PACKAGED|1.02|12|FISHERMANS MKT CRAB-FLAKE|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00072036781086|CRAB|SEAFOOD|-80.893784|80.89378752106721|272|1
35.478031|ee540ca6e9f3bfa9ae02b57fccf1f9406045a7a3|1.29|2014-11-09 12:47:00|1.4102725052409182|1|4920005675|179|0.6192084530746164|0|1|224|-80.893784|35|35.478031|SUGAR-BROWN|0.3|1|DOMINO LT BRWN SUGAR-BOX|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00049200056752|SUGAR/SUBSTITUTES|G1 GROCERY|-80.893784|1.4118628751971085|179|1
35.478031|cea7594a9b2ef6dd5793826a69ab7a3803c97415|3.35|2015-02-18 16:10:00|80.8939826282094|1|5000012734|179|35.485912169631028|0|2|341|-80.8955|57|35.4437|CREAMERS|0.0|3|COFFEEMATE SF FRENCH VANILLA|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00050000848119|MILK|DAIRY|-80.893784|80.89378752106721|272|1
35.478031|f47c0fbe4c8614aa835abbe76ebdfe0008e19f44|3.35|2015-02-16 13:51:00|1.4102725052409182|1|5000012734|179|0.6192084530746164|0|1|341|-80.893784|57|35.478031|CREAMERS|0.0|3|COFFEEMATE SF FRENCH VANILLA|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00050000848119|MILK|DAIRY|-80.893784|1.4118628751971085|179|1
35.478031|1eeff85178b729c9b1fd0a8d6865c361ee37ab2a|4.99|2014-10-04 16:22:00|80.8939826282094|1|4082201114|179|35.485912169631028|0|2|1878|-80.8955|435|35.4437|HUMMUS|2.5|6|ROASTED RED PEPPER HUMMUS|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00040822011549|SALADS|DELI|-80.893784|80.89378752106721|272|1
35.478031|78c7e75523b83efc33d4e0423f8ceaaa35907fc0|5.99|2014-09-17 16:50:00|1.4102725052409182|1|4525513785|179|0.6192084530746164|0|1|561|-80.893784|64|35.478031|FR PROD ORGANIC PRODUCE|0.0|4|ORG EDAMAME SOYBEAN SHELL|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00045255137859|FRESH PRODUCE|PRODUCE|-80.893784|1.4118628751971085|179|1
35.478031|c7192b91e543bb7f8d1249069778be1d65f3a339|3.99|2014-10-30 15:52:00|1.4102725052409182|1|7203602701|179|0.6192084530746164|0|1|1878|-80.893784|435|35.478031|HUMMUS|0.5|6|FFM ARTISAN RED PEPPER HUMMUS|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00072036027030|SALADS|DELI|-80.893784|1.4118628751971085|179|1
35.478031|88ee0346c81877d328b7f9edd2e878e3f7889bcf|1.2|2014-11-20 19:00:00|1.4102725052409182|1|68954408205|179|0.6192084530746164|0|1|685|-80.893784|61|35.478031|GREEK|0.0|3|FAGE 0% FRUYO CHERRY GREEK YOG|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00689544082033|YOGURT|DAIRY|-80.893784|1.4118628751971085|179|1
35.478031|58731bb8c1e7d47a7b3e477ad3c530e712c109ed|1.99|2014-11-12 13:02:00|1.4102725052409182|1|82415040108|179|0.6192084530746164|0|1|577|-80.893784|136|35.478031|OTHER MERCH FR MSC JUICE|0.2|4|POM POMEGRANATE JUICE 8 OZ|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00824150401087|OTHER MERCHANDISE|PRODUCE|-80.893784|1.4118628751971085|179|1
35.478031|a65c04656e588823c8f764ee5e7027c8919da48b|10.99|2015-02-20 18:28:00|80.8939826282094|1|82415040148|179|35.485912169994826|0|2|577|-80.861571|136|35.444615|OTHER MERCH FR MSC JUICE|0.0|4|POM POMEGRANATE JUICE 48 OZ|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00824150401483|OTHER MERCHANDISE|PRODUCE|-80.893784|80.893785936476448|340|1
35.478031|331729fe889a997726057f22209be44436f43c43|8.79|2014-11-29 15:18:00|1.4102725052409182|1|9955508520|179|0.6192084530746164|0|1|37|-80.893784|10|35.478031|PODS/CUPS/SINGLES|0.0|1|CARIBOU BLEND K-CUPS|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00099555089929|COFFEE|G1 GROCERY|-80.893784|1.4118628751971085|179|1
35.478031|724fd4ced595be0d4369a79ba71c29c7c7044a87|2.49|2014-10-10 18:01:00|80.8939826282094|1|60504939530|179|35.485912169631028|0|2|509|-80.8955|64|35.4437|FRESH CITRUS-REMAINING|0.0|4|LEMONS, SMALL 1LB BAG|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00605049395300|FRESH PRODUCE|PRODUCE|-80.893784|80.89378752106721|272|1
35.478031|27c7be4ff1030aa1076f016d3b32ebe6c6dd803b|2.69|2014-10-11 13:37:00|1.4102725052409182|1|30041080200|179|0.6192084530746164|0|1|4056|-80.893784|1080|35.478031|TOOTH BRUSH-PREMIUM|0.7|17|ORAL-B INDICATR SFT#10 CMPT|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00300410841003|ORAL HYGIENE|HBC|-80.893784|1.4118628751971085|179|1
35.478031|870f403b0c4dcc62544c628bc66735fd7249b5e1|3.49|2014-10-02 17:34:00|1.4102725052409182|1|3000001499|179|0.6192084530746164|0|1|60|-80.893784|9|35.478031|HOT CEREAL|0.5|1|QUAKER OATML LS MAPLE BRWN|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00030000268728|CEREAL|G1 GROCERY|-80.893784|1.4118628751971085|179|1
35.478031|903ac6c4312f11d3750a7e9584370d840d9898cf|4.79|2014-11-28 18:24:00|80.8939826282094|1|4100005152|179|35.485912168894963|0|2|273|-80.86175|43|35.40953|PREMIUM NOVELTIES|0.0|5|GH STRWBERRY SHORTCAKE BAR 6CT|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00041000053153|FROZEN NOVELTIES|FROZEN|-80.893784|80.893789467652809|209|1
35.478031|64e445c61a59321ea7e2f04974a0cad9cc7227b1|1.79|2015-01-02 14:25:00|1.4102725052409182|1|5200033875|179|0.6192084530746164|0|1|171|-80.893784|20|35.478031|ISOTONIC DRINKS|0.41|1|GATORADE LEMON LIME|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00052000338775|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.893784|1.4118628751971085|179|1
35.478031|1e1e6b5f11a7a2fffcc021ea8a2bfc205d81e724|1.79|2015-01-03 18:03:00|1.4102725052409182|1|5200033875|179|0.6192084530746164|0|1|171|-80.893784|20|35.478031|ISOTONIC DRINKS|0.41|1|GATORADE LEMON LIME|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00052000338775|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.893784|1.4118628751971085|179|1
35.478031|bca94dc25c9513d425f5c66ae0b5c333ba4512c2|1.79|2014-12-29 17:22:00|1.4102725052409182|1|5200033875|179|0.6192084530746164|0|1|171|-80.893784|20|35.478031|ISOTONIC DRINKS|0.41|1|GATORADE LEMON LIME|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00052000338775|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.893784|1.4118628751971085|179|1
35.478031|8a1bb98829e7c42e257d4199847320046c4ff727|2.29|2014-11-10 11:54:00|80.8939826282094|1|3400000007|179|35.485912169994826|0|2|48|-80.861571|7|35.444615|REGISTER GUM|0.0|1|ICE BREAKER WINTERGREEN MINTS|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00034000000098|CANDY|G1 GROCERY|-80.893784|80.893785936476448|340|1
35.478031|96fe16471320f4f1c62c7a123768ab3bfd1b00f8|5.39|2014-11-10 13:17:00|80.8939826282094|1|7027200217|179|35.485912169994826|0|2|1132|-80.861571|55|35.444615|EGGS SUBSTITUTES|0.0|3|EGGBEATER CARTON 32|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00070272002170|EGGS FRESH|DAIRY|-80.893784|80.893785936476448|340|1
35.478031|2b9ea45a9a2ed1c8a496034459dd0142476f0129|11.49|2015-03-09 10:00:00|80.8939826282094|1|20219900000|179|35.485912169631028|0|2|299|-80.8955|49|35.4437|ANGUS BEEF|1.17|2|ANGUS BEEF TOP SIRLOIN FILET|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|35.490689277687849|00202199000001|BEEF|MEAT|-80.893784|80.89378752106721|272|1
35.478031|7e99211f4d158b7a756b8496cb0663a0ebe011c3|21.99|2014-09-10 15:19:00|1.4102725052409182|1|85516500507|179|0.6192084530746164|0|1|9981|-80.893784|888|35.478031|NFS-U/PREM-OTHER RED|0.0|13|MEIOMI SONOMA PINOT NOIR|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00855165005076|ULTRA PREMIUM ($15-$19.99)|WINE|-80.893784|1.4118628751971085|179|1
35.478031|1e836a4130b33d374bf745330f1e053818597123|9.78|2014-12-17 12:16:00|1.4102725052409182|1|8660000001|179|0.6192084530746164|0|1|190|-80.893784|29|35.478031|TUNA-CANNED|1.8|1|B BEE TUNA 12 SOLID WHT ALB|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00086600000015|SEAFOOD-CANNED|G1 GROCERY|-80.893784|1.4118628751971085|179|2
35.478031|18194ce3c93897f5e5253df9085c42aa6884d06e|1.99|2014-12-29 20:21:00|1.4102725052409182|1|78616200387|179|0.6192084530746164|0|1|31|-80.893784|4|35.478031|NON CARBONATED WATER|1.0|1|FRUITWATER STRAWBERRY KIWI|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00786162003843|BOTTLED WATER|G1 GROCERY|-80.893784|1.4118628751971085|179|1
35.478031|f52fd78ebc51dd993176e78314c4b0714bfb4d5d|1.79|2014-12-30 19:01:00|1.4102725052409182|1|5200033875|179|0.6192084530746164|0|1|171|-80.893784|20|35.478031|ISOTONIC DRINKS|0.41|1|GATORADE FRUIT PUNCH|206946d510c65b5731f41e9f14c3433a83fa6341|0.544569825198699|0.61833652052202714|00052000338751|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.893784|1.4118628751971085|179|1
35.17335|03b97b8e960d708669ff0d732df4e50438fd676c|2.29|2014-12-11 21:19:00|80.709059419360486|4|2073509279|174|35.211125887094234|0|31|365|-80.780702|56|35.318911|REFRIGERATED TEAS|0.8|3|TURKEY HILL DT BLKBRY SWT TEA|225cb8f6d08d41a5afbd5f7482dbd56f6a4f5cf2|2.6102244175914993|35.187384292804154|00020735094051|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.70901|80.709064958464353|167|1
35.603432|bd8e2581fe6a1d694fd8e7fab9391ae6cd13c149|2.19|2014-10-31 15:05:00|80.895431304315082|2|7203698771|274|35.809602818987813|0|10|176|-80.875654|72|35.585842|NFS-DISPOSE CUPS|0.0|1|YH FOAM CUPS 10 OZ|2347556843de98291f71dda4542d7168a7dc9663|14.245905770413879|35.810118468028598|00072036987716|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.895009|80.895032889436251|99|1
35.603432|2b77794f99374ae2418137412f4e118937cce2dc|11.99|2014-11-18 16:25:00|80.895431304315082|2|2301286481|274|35.809602818987813|0|10|1477|-80.875654|485|35.585842|SUSHI HYBRID|0.0|6|"CHEF SAMPLER ""A"""|2347556843de98291f71dda4542d7168a7dc9663|14.245905770413879|35.810118468028598|00023012864811|SUSHI|DELI|-80.895009|80.895032889436251|99|1
35.603432|bf8a3e304f0e182aa44373a10b06ba3810f9017b|1.39|2014-10-11 16:34:00|80.895431304315082|2|2100000667|274|35.809602818987813|0|10|320|-80.875654|53|35.585842|COTTAGE CHEESE|0.39|3|BREAKSTONE 100 CAL CD PINEAPPL|2347556843de98291f71dda4542d7168a7dc9663|14.245905770413879|35.810118468028598|00021000006670|CULTURES|DAIRY|-80.895009|80.895032889436251|99|1
35.603432|2a092340ee814bfb430955d23d50f8839abd0656|2.99|2015-01-14 11:49:00|80.895431304315082|2|7090020822|274|35.809602818987813|0|10|257|-80.875654|39|35.585842|TOMATOES|0.0|1|DEI FRTLI TOMATO SC|2347556843de98291f71dda4542d7168a7dc9663|14.245905770413879|35.810118468028598|00070900501501|VEGETABLES-CAN/JAR|G1 GROCERY|-80.895009|80.895032889436251|99|1
35.603432|be39f1df02d19bbf3ba5da7908a211092e0a2e9d|3.69|2015-01-04 19:05:00|80.895431304315082|2|7127921100|274|35.809602818987813|0|10|555|-80.875654|64|35.585842|PACKAGED SALADS|0.0|4|F.E. ITALIAN SALAD MIX|2347556843de98291f71dda4542d7168a7dc9663|14.245905770413879|35.810118468028598|00071279211008|FRESH PRODUCE|PRODUCE|-80.895009|80.895032889436251|99|1
35.603432|fbdb9d721eff9f851f7afabba1cd985af10c43d2|5.39|2014-12-17 18:05:00|80.895431304315082|2|5000001547|274|35.809602818987813|0|10|152|-80.875654|24|35.585842|NFS-CAT FOOD DRY|0.6|1|FRISKIES GOURMET|2347556843de98291f71dda4542d7168a7dc9663|14.245905770413879|35.810118468028598|00050000051472|PET FOOD/SUPPLIES|G1 GROCERY|-80.895009|80.895032889436251|99|1
35.603432|62b5f4a0a5399298b59839cf8d83ab794de9df22|12.99|2014-10-16 17:23:00|80.895431304315082|2|4179021426|274|35.809602818987813|0|10|194|-80.875654|30|35.585842|OLIVE OIL|0.0|1|BERTOLLI EX VIRGIN OLIVE OIL|2347556843de98291f71dda4542d7168a7dc9663|14.245905770413879|35.810118468028598|00041790214260|SHORTENING/OIL|G1 GROCERY|-80.895009|80.895032889436251|99|1
35.603432|07af560e22a87a4dfb788d1c4ab07bc6203e25da|5.59|2015-02-01 17:06:00|80.895431304315082|2|4850002141|274|35.809602818987813|0|10|1407|-80.875654|57|35.585842|ICED COFFEE|1.1|3|STARBCKS ESPRESSO SKINNY VAN|2347556843de98291f71dda4542d7168a7dc9663|14.245905770413879|35.810118468028598|00048500021422|MILK|DAIRY|-80.895009|80.895032889436251|99|1
35.603432|ee2ddfcf0785ff7dd6847eae3bd731b11f27502c|3.49|2014-12-26 21:37:00|80.895431304315082|2|4834100016|274|35.809602818987813|0|10|3172|-80.875654|1010|35.585842|COTTON-COSMETICS-MISC|0.0|17|SWISSPERS PREM COTTON OVAL|2347556843de98291f71dda4542d7168a7dc9663|14.245905770413879|35.810118468028598|00048341000167|NAIL CARE|HBC|-80.895009|80.895032889436251|99|1
35.603432|a8028df848ead8177f89ca66bd48214d2deaf422|25.139999999999997|2015-02-10 12:17:00|80.895431304315082|2|27086500000|274|35.809602818987813|0|10|973|-80.875654|201|35.585842|FRESH PERDUE CHICKEN|1.91|2|PERDUE BONELESS CHICKEN THIGHS|2347556843de98291f71dda4542d7168a7dc9663|14.245905770413879|35.810118468028598|00270865000006|POULTRY|MEAT|-80.895009|80.895032889436251|99|4
35.603432|d522863bf96b9d556088a1b63e4ca842b4fd0769|1.82|2014-09-30 15:41:00|80.895431304315082|2||274|35.809602589256912|0|10|522|-80.861571|64|35.444615|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|2347556843de98291f71dda4542d7168a7dc9663|14.245905770413879|35.810118468028598|00204664000004|FRESH PRODUCE|PRODUCE|-80.895009|80.895388782095523|340|1
35.603432|099c21bb2ee8da539b7babed1688e3958f570f53|5.15|2014-11-07 16:59:00|80.895431304315082|2|7778200870|274|35.809602818987813|0|10|355|-80.875654|104|35.585842|FRESH GRILLING SAUSAGE|0.0|19|JVILLE GROUND SAUSAGE HOT|2347556843de98291f71dda4542d7168a7dc9663|14.245905770413879|35.810118468028598|00077782008685|DINNER SAUSAGE|CASE READY MEATS|-80.895009|80.895032889436251|99|1
35.603432|b58cfb6383da9caa20d6cf54851e23f43bbdb41b|17.98|2014-09-12 12:13:00|80.895431304315082|2|8130859207|274|35.809602818987813|0|10|9947|-80.875654|886|35.585842|NFS-PREM-CHARDONNAY|0.0|13|CB-CUPCAKE CHARDONNAY|2347556843de98291f71dda4542d7168a7dc9663|14.245905770413879|35.810118468028598|00081308592077|PREMIUM ($8-$10.99)|WINE|-80.895009|80.895032889436251|99|2
35.603432|457466fc121697c6cf167d8e90920e82bcda17ea|8.99|2015-02-10 12:14:00|80.895431304315082|2|8130859207|274|35.809602818987813|0|10|9947|-80.875654|886|35.585842|NFS-PREM-CHARDONNAY|0.0|13|CB-CUPCAKE CHARDONNAY|2347556843de98291f71dda4542d7168a7dc9663|14.245905770413879|35.810118468028598|00081308592077|PREMIUM ($8-$10.99)|WINE|-80.895009|80.895032889436251|99|1
35.603432|3437f55ee3ed8ecbe9e7d2220994c5328fd2c253|4.59|2014-09-12 19:29:00|80.895431304315082|2|5000088600|274|35.809602818987813|0|10|341|-80.875654|57|35.585842|CREAMERS|0.6|3|I/O COFFEEMATE PUMPKIN SPICE|2347556843de98291f71dda4542d7168a7dc9663|14.245905770413879|35.810118468028598|00050000886005|MILK|DAIRY|-80.895009|80.895032889436251|99|1
35.603432|6197f9577566b7d54b36f2df8d58344d3194581f|1.5|2014-11-06 18:28:00|1.4102725052409182|2|7800014945|274|0.6213971134099097|0|1|54|-80.895009|8|35.603432|DIET|0.0|23|DIET CANADA DRY TONIC WTR 1LTR|2347556843de98291f71dda4542d7168a7dc9663|14.245905770413879|0.61833652052202714|00078000149456|CARBONATED BEVERAGES|BEVERAGE|-80.895009|1.4118842554804456|274|1
35.603432|9d9da3f7ffa745293fc9a2bd88e0bc9d4a67eede|17.99|2014-11-01 15:55:00|80.895431304315082|2|3774125400|274|35.809602818987813|0|10|6965|-80.875654|1586|35.585842|GM READING GLASSES|0.0|18|GREEN READERS-BAMBOO TEMPLE|2347556843de98291f71dda4542d7168a7dc9663|14.245905770413879|35.810118468028598|00037741254027|READING GLASSES|GM|-80.895009|80.895032889436251|99|1
35.219587|18d00f53a397819d4e97a64e991927ce66b837c0|1.69|2014-12-05 07:48:00|80.810069425230125|4|4900000044|401|35.25592770327497|0|23|55|-80.86175|8|35.40953|REGULAR|0.0|23|CB COKE SINGLE 20 OZ.|2652315c0c7f49a1b4a347b32fdb2627dd1c0a2b|2.511058633269311|35.240679762029046|00049000000443|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.810133371722287|209|1
35.219587|a5e6a3670f76d34909534b52a0ac871c84e37d17|3.65|2014-12-04 07:57:00|80.810069425230125|4|3010067264|401|35.25592770327497|0|23|91|-80.86175|13|35.40953|SPRAYED BUTTER CRACKERS|1.15|1|TOWN HOUSE FLATBRD ITALIAN HRB|2652315c0c7f49a1b4a347b32fdb2627dd1c0a2b|2.511058633269311|35.240679762029046|00030100506591|CRACKERS|G1 GROCERY|-80.810056|80.810133371722287|209|1
35.152722|6bd8906d9f84dafbea874dddb4edfba9efe2d8cb|4.99|2014-11-04 17:48:00|1.4094857484078087|1|7597140209|160|0.613530739938246|0|26|1845|-80.825175|425|35.152722|FFM PRESLICED CHEESE|0.0|6|F.F.COLBY JACK CHEDDAR  CHEESE|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00072036010315|PRESLICED CHEESE|DELI|-80.825175|1.4106654222506079|160|1
35.152722|0e5d6e8d6bc210eed84e154d27e769d995472580|4.99|2014-11-15 13:41:00|1.4094857484078087|1|7597140209|160|0.613530739938246|0|26|1845|-80.825175|425|35.152722|FFM PRESLICED CHEESE|0.0|6|F.F.COLBY JACK CHEDDAR  CHEESE|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00072036010315|PRESLICED CHEESE|DELI|-80.825175|1.4106654222506079|160|1
35.152722|9e101adfc029439927b25063eb75edeb38e9d8ce|4.99|2014-09-16 16:24:00|1.4094857484078087|1|7597140209|160|0.613530739938246|0|26|1845|-80.825175|425|35.152722|FFM PRESLICED CHEESE|0.0|6|F.F.COLBY JACK CHEDDAR  CHEESE|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00072036010315|PRESLICED CHEESE|DELI|-80.825175|1.4106654222506079|160|1
35.152722|137d9273385eea7b353a7ad32e6a99b92874474e|3.99|2014-11-16 10:37:00|1.4094857484078087|1|7127927100|160|0.613530739938246|0|26|555|-80.825175|64|35.152722|PACKAGED SALADS|0.0|4|F.E. BABY SPINACH|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00071279271002|FRESH PRODUCE|PRODUCE|-80.825175|1.4106654222506079|160|1
35.152722|d608932d9d0c9a9c6e6e4958d0b08b445c20b315|4.99|2014-10-15 18:32:00|1.4094857484078087|1|7597140209|160|0.613530739938246|0|26|1845|-80.825175|425|35.152722|FFM PRESLICED CHEESE|0.0|6|F.F.COLBY JACK CHEDDAR  CHEESE|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00072036010315|PRESLICED CHEESE|DELI|-80.825175|1.4106654222506079|160|1
35.152722|028053d3f8ded0b24996b30570a956e1f1a71693|4.59|2014-09-13 11:28:00|1.4094857484078087|1|7203636053|160|0.613530739938246|0|26|31|-80.825175|4|35.152722|NON CARBONATED WATER|1.59|1|(U)HT SPRING WATER .5 LTR 24PK|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00072036360533|BOTTLED WATER|G1 GROCERY|-80.825175|1.4106654222506079|160|1
35.152722|50c4e2e9f8bcb70ba4dc9c1227e7f6dcec66dd86|4.49|2014-11-25 16:48:00|1.4094857484078087|1|7203636053|160|0.613530739938246|0|26|31|-80.825175|4|35.152722|NON CARBONATED WATER|1.15|1|(U)HT SPRING WATER .5 LTR 24PK|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00072036360533|BOTTLED WATER|G1 GROCERY|-80.825175|1.4106654222506079|160|1
35.152722|5c81f7e4b3b6a509b2a4a746bdd89a10b3337fc1|4.49|2014-10-07 16:28:00|1.4094857484078087|1|7203636053|160|0.613530739938246|0|26|31|-80.825175|4|35.152722|NON CARBONATED WATER|1.49|1|(U)HT SPRING WATER .5 LTR 24PK|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00072036360533|BOTTLED WATER|G1 GROCERY|-80.825175|1.4106654222506079|160|1
35.152722|464be150e57e8b87170d2610283956f290c38eca|13.47|2015-01-28 17:42:00|1.4094857484078087|1|7203636053|160|0.613530739938246|0|26|31|-80.825175|4|35.152722|NON CARBONATED WATER|3.4699999999999998|1|(U)HT SPRING WATER .5 LTR 24PK|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00072036360533|BOTTLED WATER|G1 GROCERY|-80.825175|1.4106654222506079|160|3
35.152722|921fad8016bd106ebca189d876b6f2325f083fd3|2.99|2014-12-22 19:08:00|1.4094857484078087|1|4760001111|160|0.613530739938246|0|26|1246|-80.825175|34|35.152722|SPICE BLENDS|0.0|1|WEBER KICK'N CHICKEN|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00047600011036|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.825175|1.4106654222506079|160|1
35.152722|b7175b657beffbfc5b22a0f58ba29d5c2053d407|7.99|2015-02-08 10:12:00|1.4094857484078087|1|4175705920|160|0.613530739938246|0|26|2018|-80.825175|505|35.152722|PRESSED CHEESE|0.0|6|MINI BABYBEL GOUDA 10CT|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00041757680473|SPECIALTY CHEESE|DELI|-80.825175|1.4106654222506079|160|1
35.152722|49103f2a2e05785c5133c780b1180a2e351b82f1|7.99|2014-12-29 22:57:00|1.4094857484078087|1|3680025145|160|0.613530739938246|0|26|4885|-80.825175|1240|35.152722|ANTI-FUNGAL TREATMENTS/DEOD|2.4|17|TC ATHLETES FT CRM|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00036800251458|FOOT CARE|HBC|-80.825175|1.4106654222506079|160|1
35.152722|66e2b0c0f03fcf51c8a221bafce87033b7de006a|1.99|2014-11-21 18:44:00|1.4094857484078087|1|3900004504|160|0.613530739938246|0|26|114|-80.825175|14|35.152722|PUMPKIN|0.2|1|LIBBY SOLID PACK PUMPKIN|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00039000045049|DESSERTS/GELS/SYRUPS|G1 GROCERY|-80.825175|1.4106654222506079|160|1
35.152722|e646a33927de408d595ce998bc67d3b050b1bed6|3.75|2014-12-14 12:38:00|1.4094857484078087|1|4139000107|160|0.613530739938246|0|26|79|-80.825175|273|35.152722|ASIAN SAUCES/SEASONINGS|0.96|1|KIKKOMAN SOY SAUCE LT 15|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00041390001079|ASIAN PREP. FOODS|G1 GROCERY|-80.825175|1.4106654222506079|160|1
35.152722|d6a70cd76f25df3262c1c06c7792a3a231712bd0|3.34|2014-11-27 08:52:00|1.4094857484078087|1||160|0.613530739938246|0|26|562|-80.825175|64|35.152722|FRESH CUT FRUIT|0.0|4|SLICED STRAWBERRIES BY/LB|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00204217000000|FRESH PRODUCE|PRODUCE|-80.825175|1.4106654222506079|160|1
35.152722|3472dae267331fefef4c102c9002a5b3155a28d0|1.29|2015-02-21 18:40:00|1.4094857484078087|1||160|0.613530739938246|0|26|508|-80.825175|64|35.152722|FRESH GRAPEFRUIT|0.29|4|RED GRAPEFRUIT, FL  LRG|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00204281000005|FRESH PRODUCE|PRODUCE|-80.825175|1.4106654222506079|160|1
35.152722|44e44de43de10483258a7f11b23e980bd0aef85f|29.99|2014-09-23 19:34:00|1.4094857484078087|1|20545100000|160|0.613530739938246|0|26|1290|-80.825175|381|35.152722|LOCAL CAKES|0.0|14|"TIZ'S 8""  DECO CHOC TRUFF CAKE"|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00205451000009|CAKES|BAKERY|-80.825175|1.4106654222506079|160|1
35.152722|81ccd97a9e7db66b6d9cb652b9b84a68c60be7ab|8.44|2014-12-13 18:27:00|80.825044058860698|1||160|35.1702275358397|0|29|529|-80.85013|64|35.175855|FRESH ASPARAGUS|0.0|4|GREEN  ASPARAGUS|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00204080000008|FRESH PRODUCE|PRODUCE|-80.825175|80.825177734975583|218|2
35.152722|b324193311c637b8b7ffe336c7ce837ba846453d|2.58|2014-11-11 16:29:00|1.4094857484078087|1||160|0.613530739938246|0|26|508|-80.825175|64|35.152722|FRESH GRAPEFRUIT|0.29|4|RED GRAPEFRUIT, FL  LRG|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00204281000005|FRESH PRODUCE|PRODUCE|-80.825175|1.4106654222506079|160|2
35.152722|35afa41e31f5cb76932b30a8313f9fa9492806b5|12.9|2015-02-23 19:31:00|1.4094857484078087|1||160|0.613530739938246|0|26|508|-80.825175|64|35.152722|FRESH GRAPEFRUIT|0.29|4|RED GRAPEFRUIT, FL  LRG|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00204281000005|FRESH PRODUCE|PRODUCE|-80.825175|1.4106654222506079|160|10
35.152722|da94e680311be093c89507b4d65b8d663366fe4c|4.49|2014-12-23 15:19:00|1.4094857484078087|1|74759930652|160|0.613530739938246|0|26|62|-80.825175|7|35.152722|SPECIALTY BAR/BOX CHOCOLATE|0.0|1|GHIRADELLI DK CHOC MINT SQUARE|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00747599306525|CANDY|G1 GROCERY|-80.825175|1.4106654222506079|160|1
35.152722|6a11eee129307888128592720a72ad299b5f3237|7.99|2014-12-26 16:39:00|1.4094857484078087|1|30067208611|160|0.613530739938246|0|26|4243|-80.825175|1200|35.152722|NASAL PRODUCT-ADULT|0.0|17|4-WAY FAST ACTING NASAL SPRAY|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00300672086112|COUGH/COLD/SINUS|HBC|-80.825175|1.4106654222506079|160|1
35.152722|dda167890409e353dd09307359ae025bba827ee2|2.17|2014-10-12 18:07:00|80.825044058860698|1||160|35.17022753420661|0|29|524|-80.844274|64|35.204336|FRESH PROD FRESH ONIONS|0.0|4|COO PEELED RED ONIONS|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00204667000001|FRESH PRODUCE|PRODUCE|-80.825175|80.825184645071957|61|1
35.152722|11fa8c88f22006072f26d401e55a7a991048b846|1.55|2014-11-13 15:33:00|1.4094857484078087|1|8000051306|160|0.613530739938246|0|26|189|-80.825175|29|35.152722|TUNA-POUCH|0.05|1|STARKIST TUNA PCH LS CHNK LGHT|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00080000505279|SEAFOOD-CANNED|G1 GROCERY|-80.825175|1.4106654222506079|160|1
35.152722|5766c9cfc0f92c5ca6f196f0cdd375edaf53bac8|4.29|2015-03-05 15:57:00|1.4094857484078087|1|9418456083|160|0.613530739938246|0|26|583|-80.825175|136|35.152722|NUTS|0.0|4|TROPICAL CRYSTALLIZED GINGER|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00094184560832|OTHER MERCHANDISE|PRODUCE|-80.825175|1.4106654222506079|160|1
35.152722|b9f9b63bb9ade272a6acf5d518356e2cc3f31126|4.79|2014-11-19 21:16:00|80.825044058860698|1|18685200031|160|35.170227533599295|0|29|275|-80.85753|45|35.116638|SUPER PREMIUM ICE CREAM|2.4|5|TALENTI SIMPLY STRWBRRY GELATO|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00186852000488|ICE CREAM|FROZEN|-80.825175|80.825186173210739|204|1
35.152722|e3fd6c064e503444b36a98a47911e4eb066a5f0c|3.49|2014-12-20 13:42:00|1.4094857484078087|1|4178000211|160|0.613530739938246|0|26|202|-80.825175|31|35.152722|PRETZELS|0.99|1|UTZ POLY BAG WHEEL PRETZELS|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00041780002587|SNACKS|G1 GROCERY|-80.825175|1.4106654222506079|160|1
35.152722|945dfdaf525a1107e99495ef1ae43f808ed70ba9|3.59|2014-09-12 16:44:00|1.4094857484078087|1|4850002013|160|0.613530739938246|0|26|335|-80.825175|56|35.152722|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA PP HOMESTYLE|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00048500301395|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.825175|1.4106654222506079|160|1
35.152722|78a8e20af4b2f353c37928558d068d0327cab3ce|4.49|2014-12-10 20:38:00|80.825044058860698|1|70897191697|160|35.1702275358397|0|29|1703|-80.85013|387|35.175855|SEASONAL COOKIES|1.0|14|RED VELVET FRSTD SUGAR COOKIES|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00708971916978|COOKIES|BAKERY|-80.825175|80.825177734975583|218|1
35.152722|1341d91f786d68594a0f5ea82e44bd1a2d5d33cc|15.98|2015-01-21 22:48:00|1.4094857484078087|1|76722602504|160|0.613530739938246|0|26|1279|-80.825175|48|35.152722|SINGLE SERVE FLAVOR|0.0|5|SUKHIS CHICKEN CURRY|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00767226025049|FROZEN MEALS|FROZEN|-80.825175|1.4106654222506079|160|2
35.152722|2cccdfa9cbe26d8f50a690d4b5d4f6c6b152ba08|7.49|2015-02-12 18:52:00|80.825044058860698|1|76108880053|160|35.170227534767925|0|29|1941|-80.824767|465|35.116751|COLD PREP FOODS MEALS|0.0|6|CHICKEN TIKKA W/JASMINE RICE|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00761088800530|COLD PREPARED FOODS|DELI|-80.825175|80.825182976425793|294|1
35.152722|e23915f017756a1f0b63e65c2b170f44bee39c16|3.99|2015-01-07 17:21:00|1.4094857484078087|1|75535500511|160|0.613530739938246|0|26|205|-80.825175|31|35.152722|REMAINING SNACKS|2.0|1|GOOD HEALTH NAT VEGGIE CHIPS|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00755355005155|SNACKS|G1 GROCERY|-80.825175|1.4106654222506079|160|1
35.152722|6ae25cff10c616276f74dfd33208d6437deb8366|2.85|2015-02-15 16:37:00|1.4094857484078087|1|1380010321|160|0.613530739938246|0|26|1279|-80.825175|48|35.152722|SINGLE SERVE FLAVOR|0.0|5|STOUFFER CREAMED CHIP BEEF|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00013800100184|FROZEN MEALS|FROZEN|-80.825175|1.4106654222506079|160|1
35.152722|dc58734573214bab28f3d43ddd4a499c1f424afc|5.78|2014-11-08 10:54:00|1.4094857484078087|1|1380010321|160|0.613530739938246|0|26|1279|-80.825175|48|35.152722|SINGLE SERVE FLAVOR|0.78|5|STOUFFER CREAMED CHIP BEEF|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00013800100184|FROZEN MEALS|FROZEN|-80.825175|1.4106654222506079|160|2
35.152722|64d02d73bf3b66a640d1e79ea226e440705d5854|4.49|2014-09-28 21:35:00|80.825044058860698|1|88491201426|160|35.170227503380175|0|29|74|-80.780702|9|35.318911|RTE CEREAL ALL FAMILY|0.0|1|POST HNY BUNCHES FAM HNY RSTD|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00884912014269|CEREAL|G1 GROCERY|-80.825175|80.825216325854655|167|1
35.152722|803bb9c7c7186e687ccaf92ebff672a6c9353794|2.99|2015-01-21 16:43:00|1.4094857484078087|1|1380004717|160|0.613530739938246|0|26|1278|-80.825175|48|35.152722|SINGLE SERVE NUTRITIONAL|0.0|5|LC CAFE CLSSC PEPPERONI PIZZA|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00013800047175|FROZEN MEALS|FROZEN|-80.825175|1.4106654222506079|160|1
35.152722|6f8092de7b4d2d1dcef30e3f5c49726624fc452e|9.99|2014-11-22 13:53:00|1.4094857484078087|1|3700080900|160|0.613530739938246|0|26|403|-80.825175|69|35.152722|NFS-RUG CLEANERS|0.0|1|SWIFFER DUSTER EXT HANDLE|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00037000809005|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.825175|1.4106654222506079|160|1
35.152722|4258d2ee520733d84fc4ddb0b1ca311b2e43ecb3|2.99|2014-11-10 11:29:00|80.825044058860698|1|5250006714|160|35.170227491957206|0|29|182|-80.764523|28|35.341927|MAYO|0.0|1|DUKES MAYO 11.5 SQZ|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00052500067144|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.825175|80.825223022923083|220|1
35.152722|2cf51a50d8423a6d8f7b1a6086bf6a6b98c4866d|13.58|2014-09-20 14:50:00|1.4094857484078087|1|4900002890|160|0.613530739938246|0|26|54|-80.825175|8|35.152722|DIET|3.4|23|DIET COKE W/SPLENDA 12 OZ FRID|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00049000042696|CARBONATED BEVERAGES|BEVERAGE|-80.825175|1.4106654222506079|160|2
35.152722|0167de3e31203e338ee5208edec4157769319d9a|5.89|2014-10-26 16:26:00|1.4094857484078087|1|5210082791|160|0.613530739938246|0|26|1245|-80.825175|34|35.152722|SINGLE SPICES|0.0|1|MC GOURMET ORG OREGANO LEAVES|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00052100827919|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.825175|1.4106654222506079|160|1
35.152722|4709e26daef00b6278d133be096cb5fc89333dee|2.19|2015-03-05 21:04:00|80.825044058860698|1|4900005010|160|35.1702275358397|0|29|54|-80.85013|8|35.175855|DIET|0.2|23|DT CLASSIC 2 LITER|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00049000050110|CARBONATED BEVERAGES|BEVERAGE|-80.825175|80.825177734975583|218|1
35.152722|22f146ebf3ab1d7abfb5f7df785dc32e2e0aa1cc|2.49|2015-02-12 13:00:00|1.4094857484078087|1|7156766109|160|0.613530739938246|0|26|52|-80.825175|7|35.152722|PKG NON CHOC|0.0|1|JBELLY 20 FLAVORS|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00071567661096|CANDY|G1 GROCERY|-80.825175|1.4106654222506079|160|1
35.152722|ac5200c97ac796f590d99e4b87ae1373225db167|5.69|2014-11-11 16:02:00|80.825044058860698|1|1450000711|160|35.170227491957206|0|29|1274|-80.764523|50|35.341927|BAG VEG PROTEIN|0.0|5|BE VOILA 3 CHS CHICKEN|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00014500007131|VEGETABLES-FROZEN|FROZEN|-80.825175|80.825223022923083|220|1
35.152722|26e1356acc72db17b28789b22d56bdfdeb0e280b|6.78|2014-12-18 15:47:00|1.4094857484078087|1|2113150605|160|0.613530739938246|0|26|1279|-80.825175|48|35.152722|SINGLE SERVE FLAVOR|1.78|5|M CALLENDER CHICKEN TERIYAKI|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00021131800406|FROZEN MEALS|FROZEN|-80.825175|1.4106654222506079|160|2
35.152722|3df935dbf61ecd117d775bd32847e220a8f90bed|3.39|2014-11-25 08:11:00|80.825044058860698|1|2113150605|160|35.170227491957206|0|29|1279|-80.764523|48|35.341927|SINGLE SERVE FLAVOR|0.0|5|M CALLENDER CHICKEN TERIYAKI|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00021131800406|FROZEN MEALS|FROZEN|-80.825175|80.825223022923083|220|1
35.152722|be4590365adff9a9d8bb4d9ca9f3f72f2837c47d|3.39|2014-12-30 15:57:00|1.4094857484078087|1|2113150605|160|0.613530739938246|0|26|1279|-80.825175|48|35.152722|SINGLE SERVE FLAVOR|0.0|5|M CALLENDER CHICKEN TERIYAKI|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00021131800406|FROZEN MEALS|FROZEN|-80.825175|1.4106654222506079|160|1
35.152722|48c019275022bc2e60cacccb9b89339168bbf961|3.35|2014-11-11 08:29:00|80.825044058860698|1|1600045723|160|35.170227491957206|0|29|42|-80.764523|6|35.341927|GRANOLA/YOGURT BARS|0.0|1|NV BAR PROT COCONUT ALMOND|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00016000485426|BREAKFAST FOODS|G1 GROCERY|-80.825175|80.825223022923083|220|1
35.152722|c38da040300c6e9346ab9bf30d37a8d6d4728447|3.39|2015-01-02 09:31:00|80.825044058860698|1|2113150605|160|35.170227491957206|0|29|1279|-80.764523|48|35.341927|SINGLE SERVE FLAVOR|0.0|5|M CALLENDER CHICKEN TERIYAKI|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00021131800406|FROZEN MEALS|FROZEN|-80.825175|80.825223022923083|220|1
35.152722|d544e5c06b2c3e8fc36634586bca07e7463f1795|3.39|2014-12-04 10:59:00|80.825044058860698|1|2113150605|160|35.170227503380175|0|29|1279|-80.780702|48|35.318911|SINGLE SERVE FLAVOR|0.0|5|M CALLENDER COUNTRY PRK RIBLET|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00021131800307|FROZEN MEALS|FROZEN|-80.825175|80.825216325854655|167|1
35.152722|140d6dca089a415e3d43801a13ad907613a079ae|3.99|2014-10-19 09:03:00|1.4094857484078087|1|1600027534|160|0.613530739938246|0|26|81|-80.825175|9|35.152722|RTE CEREAL KIDS|0.0|1|GM LUCKY CHARMS  11.5OZ|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00016000275348|CEREAL|G1 GROCERY|-80.825175|1.4106654222506079|160|1
35.152722|e35208331537709932553ea408f5c5b0a03fc6ac|3.39|2014-12-04 14:37:00|1.4094857484078087|1|2113150605|160|0.613530739938246|0|26|1279|-80.825175|48|35.152722|SINGLE SERVE FLAVOR|0.0|5|M CALLENDER CHICKEN TERIYAKI|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00021131800406|FROZEN MEALS|FROZEN|-80.825175|1.4106654222506079|160|1
35.152722|232dba165c5a8b18681f6eeacad458d73252dd9d|6.29|2015-01-15 17:21:00|1.4094857484078087|1|5150072001|160|0.613530739938246|0|26|125|-80.825175|19|35.152722|PEANUT BUTTER|0.0|1|JIF CREAMY PEANUT BUTTER|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00051500720011|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.825175|1.4106654222506079|160|1
35.152722|8e7ed3a3647351d87ff7ce262150866685da1d1b|89.99|2014-11-01 15:06:00|1.4094857484078087|1|7217923171|160|0.613530739938246|0|26|6034|-80.825175|1544|35.152722|COFFEE APPLIANCE|0.0|18|MR. COFFEE SINGLE SERVE SYSTEM|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00072179231714|APPLIANCES|GM|-80.825175|1.4106654222506079|160|1
35.152722|cb1092fa6c5f7b29abd9e9acf7d8048baec34d90|3.79|2014-12-22 21:09:00|80.825044058860698|1|7203688184|160|35.170227491957206|0|29|555|-80.764523|64|35.341927|PACKAGED SALADS|0.0|4|HTT ASIAN CHOP SALAD KIT|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00072036881847|FRESH PRODUCE|PRODUCE|-80.825175|80.825223022923083|220|1
35.152722|e552fa545ccd1703b79419fba7b496c65928d351|2.29|2014-11-26 18:16:00|1.4094857484078087|1|7675311860|160|0.613530739938246|0|26|5852|-80.825175|1538|35.152722|KITCHEN GAD CAN OPENERS|1.15|18|GOODCOOK CAN TAPPER SET 11860|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00076753118606|KITCHEN GADGETS|GM|-80.825175|1.4106654222506079|160|1
35.152722|e9fb089742d5396724006c1297c65023dc186e7f|2.87|2014-11-28 22:21:00|80.825044058860698|1|8130831863|160|35.170227534617439|0|29|9935|-80.806073|885|35.106477|NFS POP CAB SAUV|0.0|13|OAK CREEK CABERNET|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00081308318639|POPULAR (4-$7.99)|WINE|-80.825175|80.82518345614416|4|1
35.152722|75fcf81bffd8864109fe1eee4755a32339ce95af|16.58|2015-01-12 11:31:00|1.4094857484078087|1|9955508510|160|0.613530739938246|0|26|1247|-80.825175|37|35.152722|SINGLES PODS CUPS TEA|0.0|1|BIGELOW K CUP TEA GREEN|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00099555085136|TEA|G1 GROCERY|-80.825175|1.4106654222506079|160|2
35.152722|69eb8422d0477c4af164897791230a7aebb78edd|9.99|2014-12-05 16:15:00|1.4094857484078087|1|8858660384|160|0.613530739938246|0|26|9947|-80.825175|886|35.152722|NFS-PREM-CHARDONNAY|0.0|13|CB-CH ST MICH CHARDONNAY|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00088586603846|PREMIUM ($8-$10.99)|WINE|-80.825175|1.4106654222506079|160|1
35.152722|d30ef953b67a32f0415b854bd1d33c9aa7b6f726|5.99|2015-03-02 19:36:00|80.825044058860698|1|1834175105|160|35.170227534767925|0|29|9934|-80.824767|885|35.116751|NFS POP CHARDONNAY|0.0|13|CB-BAREFOOT CHARDONNAY|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00018341751055|POPULAR (4-$7.99)|WINE|-80.825175|80.825182976425793|294|1
35.152722|90dea0728acaae8d36fb1026413575d36c7a28fb|3.39|2015-01-09 10:03:00|80.825044058860698|1|2113150605|160|35.170227491957206|0|29|1279|-80.764523|48|35.341927|SINGLE SERVE FLAVOR|0.89|5|M CALLENDER MTBALL SAUS MARINA|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00021131800369|FROZEN MEALS|FROZEN|-80.825175|80.825223022923083|220|1
35.152722|d027645b1bde40523df44ebe0a656c083ca3b6df|6.78|2014-12-02 18:57:00|1.4094857484078087|1|2113150605|160|0.613530739938246|0|26|1279|-80.825175|48|35.152722|SINGLE SERVE FLAVOR|0.0|5|M CALLENDER MTBALL SAUS MARINA|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00021131800369|FROZEN MEALS|FROZEN|-80.825175|1.4106654222506079|160|2
35.152722|a2753eadc49f8014b7dcf537ae531894be1423a5|3.39|2014-10-14 12:28:00|80.825044058860698|1|2113150605|160|35.170227491957206|0|29|1279|-80.764523|48|35.341927|SINGLE SERVE FLAVOR|0.89|5|M CALLENDER MTBALL SAUS MARINA|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00021131800369|FROZEN MEALS|FROZEN|-80.825175|80.825223022923083|220|1
35.152722|af03a33053bacebc1e3abd638f7e4a6b4b518890|20.97|2015-01-04 10:40:00|1.4094857484078087|1|4900002890|160|0.613530739938246|0|26|54|-80.825175|8|35.152722|DIET|4.99|23|DIET COKE 12OZ 12PK FRIDGE CAN|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00049000028911|CARBONATED BEVERAGES|BEVERAGE|-80.825175|1.4106654222506079|160|3
35.152722|9cddbb6e75c78ab2c8c634602c1637e41d72a085|6.79|2014-12-09 14:28:00|1.4094857484078087|1|4900002890|160|0.613530739938246|0|26|54|-80.825175|8|35.152722|DIET|1.8|23|DIET COKE 12OZ 12PK FRIDGE CAN|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00049000028911|CARBONATED BEVERAGES|BEVERAGE|-80.825175|1.4106654222506079|160|1
35.152722|5f09407d4621c204bda0e507f6fb1348b24565a3|4.99|2015-02-09 18:00:00|80.825044058860698|1|5210000247|160|35.170227534767925|0|29|1245|-80.824767|34|35.116751|SINGLE SPICES|0.0|1|MC CURRY POWDER|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00052100002477|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.825175|80.825182976425793|294|1
35.152722|a4f95f64ba657b2797e27928b9d2a2740e2306cc|6.79|2014-11-09 18:31:00|80.825044058860698|1|4900002890|160|35.1702275358397|0|29|54|-80.85013|8|35.175855|DIET|1.8|23|DIET COKE 12OZ 12PK FRIDGE CAN|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00049000028911|CARBONATED BEVERAGES|BEVERAGE|-80.825175|80.825177734975583|218|1
35.152722|9b5ae8139a0c0169751bb833d3267c6ca8c4308c|13.58|2014-12-16 15:43:00|80.825044058860698|1|4900002890|160|35.170227491957206|0|29|54|-80.764523|8|35.341927|DIET|3.6|23|DIET COKE 12OZ 12PK FRIDGE CAN|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00049000028911|CARBONATED BEVERAGES|BEVERAGE|-80.825175|80.825223022923083|220|2
35.152722|952a7c30fb788cdabbc3ece24d091d2048c916dc|1.2|2014-11-20 17:28:00|1.4094857484078087|1|7047000641|160|0.613530739938246|0|26|688|-80.825175|61|35.152722|LIGHT|0.0|3|YOPLAIT LIGHT CHERRY|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00070470006536|YOGURT|DAIRY|-80.825175|1.4106654222506079|160|2
35.152722|47c135aff5e940a5f824ccb30f90bcdc359f8f04|8.99|2014-12-31 16:03:00|1.4094857484078087|1|8500001437|160|0.613530739938246|0|26|9939|-80.825175|885|35.152722|NFS POP PINOT NOIR|0.0|13|BELLA SERA PINOT NOIR|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00085000014370|POPULAR (4-$7.99)|WINE|-80.825175|1.4106654222506079|160|1
35.152722|87ad96e17100c12da857d27e4c407fb96b45a1bc|8.19|2015-01-12 19:03:00|80.825044058860698|1|9955509849|160|35.170227534822438|0|29|1247|-80.80146|37|35.17739|SINGLES PODS CUPS TEA|0.0|1|CELESTIAL K CUP SLEEPYTIME|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00099555098495|TEA|G1 GROCERY|-80.825175|80.825182795370594|208|1
35.152722|1e8b968ca1ce4e6474ff538b38ca15477ae33ab7|6.49|2014-09-27 12:31:00|1.4094857484078087|1|76108880034|160|0.613530739938246|0|26|1941|-80.825175|465|35.152722|COLD PREP FOODS MEALS|0.0|6|HAND ROLLED CHICKEN BURRITTOS|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00761088800349|COLD PREPARED FOODS|DELI|-80.825175|1.4106654222506079|160|1
35.152722|b4f207ab8289569506556164116158901aff91ab|5.49|2014-09-28 09:56:00|1.4094857484078087|1|72822912347|160|0.613530739938246|0|26|201|-80.825175|31|35.152722|POTATO CHIPS|0.0|1|TERRA CHIPS MEDITERRANEAN|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00728229123477|SNACKS|G1 GROCERY|-80.825175|1.4106654222506079|160|1
35.152722|f6ee70a867e2e6d3434216b5b8dc9998f588e53d|0.95|2014-10-09 09:55:00|80.825044058860698|1|61300871771|160|35.170227533599295|0|29|99|-80.85753|32|35.116638|LIQUID TEA|0.0|1|ARIZONA DIET GREEN TEA|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00613008720711|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.825175|80.825186173210739|204|1
35.152722|62b2667293609912ecf5829b9fc7ea58dd0dbe97|0.95|2014-10-14 09:52:00|80.825044058860698|1|61300871771|160|35.170227533599295|0|29|99|-80.85753|32|35.116638|LIQUID TEA|0.48|1|ARIZONA DIET GREEN TEA|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00613008720711|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.825175|80.825186173210739|204|1
35.152722|98d99a7e331f01c65e3c01b1b78c1909cf98aaa3|0.95|2014-12-09 09:53:00|80.825044058860698|1|61300871771|160|35.170227533599295|0|29|99|-80.85753|32|35.116638|LIQUID TEA|0.2|1|ARIZONA DIET GREEN TEA|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00613008720711|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.825175|80.825186173210739|204|1
35.152722|8a865e262d7232106499675822f0e4abc36d29ce|3.69|2014-11-05 17:53:00|1.4094857484078087|1|71514172928|160|0.613530739938246|0|26|330|-80.825175|55|35.152722|EGGS|0.0|3|EGGLAND BEST GRADE A EX-LG EGG|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00715141729283|EGGS FRESH|DAIRY|-80.825175|1.4106654222506079|160|1
35.152722|2b4c52d3d1964d77c3293865c9647c388f016e19|0.95|2015-02-05 09:46:00|80.825044058860698|1|61300871771|160|35.170227533599295|0|29|99|-80.85753|32|35.116638|LIQUID TEA|0.15|1|ARIZONA DIET GREEN TEA|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00613008720711|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.825175|80.825186173210739|204|1
35.152722|066b9ebb875eb7625417c27955c1c04591ba465d|0.95|2015-01-03 13:36:00|80.825044058860698|1|61300871771|160|35.170227533599295|0|29|99|-80.85753|32|35.116638|LIQUID TEA|0.15|1|ARIZONA DIET GREEN TEA|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00613008720711|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.825175|80.825186173210739|204|1
35.152722|f3c1290bfe45155cb713396c9ce5bacc25b70b22|0.95|2015-02-10 09:45:00|80.825044058860698|1|61300871771|160|35.170227533599295|0|29|99|-80.85753|32|35.116638|LIQUID TEA|0.15|1|ARIZONA DIET GREEN TEA|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00613008720711|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.825175|80.825186173210739|204|1
35.152722|a7ca2a0d9eea12761080f46df5b5789fc2a01d0d|5.74|2015-03-08 16:42:00|1.4094857484078087|1|7203698594|160|0.613530739938246|0|26|403|-80.825175|69|35.152722|NFS-RUG CLEANERS|0.0|1|YH FLOOR MOPPING CLOTHS|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00072036985965|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.825175|1.4106654222506079|160|2
35.152722|ff80e71649273fa2fede69cb01192e7494a493b2|7.02|2014-12-06 14:06:00|1.4094857484078087|1||160|0.613530739938246|0|26|500|-80.825175|64|35.152722|FRESH APPLES|0.0|4|HONEY CRISP APPLE|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00233283000003|FRESH PRODUCE|PRODUCE|-80.825175|1.4106654222506079|160|1
35.152722|e33344e89e5224de2ba74ed342465d99e95ce220|9.58|2014-10-28 13:25:00|1.4094857484078087|1||160|0.613530739938246|0|26|500|-80.825175|64|35.152722|FRESH APPLES|2.88|4|HONEY CRISP APPLE|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00233283000003|FRESH PRODUCE|PRODUCE|-80.825175|1.4106654222506079|160|1
35.152722|b1a32e6d6e8bc8567c37797654c906a901f3a4ff|6.94|2014-12-12 18:04:00|1.4094857484078087|1||160|0.613530739938246|0|26|500|-80.825175|64|35.152722|FRESH APPLES|0.0|4|HONEY CRISP APPLE|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00233283000003|FRESH PRODUCE|PRODUCE|-80.825175|1.4106654222506079|160|1
35.152722|5811c1eb534ae4c4904afae1c2554e75783e7faf|3.49|2014-11-28 15:32:00|1.4094857484078087|1|85225100001|160|0.613530739938246|0|26|339|-80.825175|57|35.152722|EGGNOGS/DRINKS|0.5|3|I/O SUTHRN COMF EGG NOG|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00852251000014|MILK|DAIRY|-80.825175|1.4106654222506079|160|1
35.152722|44c096c098a48bf86a64ae7154f3a117619fc96e|16.99|2015-01-31 17:38:00|80.825044058860698|1|71280845554|160|35.170227504438287|0|29|458|-80.737839|82|35.297134|CRAFT BEER|0.0|16|HIGHLAND MTN MEDLEY SMPLR 12PK|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00712808455547|DOMESTIC BEER|BEER|-80.825175|80.825215649707076|258|1
35.152722|ead5cdb20dd815a6bfb9b0319c3b84f1d31a39e9|5.48|2014-10-14 18:27:00|80.825044058860698|1|20165700000|160|35.170227534767925|0|29|297|-80.824767|49|35.116751|GROUND BEEF|0.61|2|HT GROUND BEEF CHUCK 80% LEAN|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00201657000003|BEEF|MEAT|-80.825175|80.825182976425793|294|1
35.152722|868bc8d87b66c1b384254f30fdd5a4bc51aa0e9d|3.65|2015-01-19 20:20:00|1.4094857484078087|1|7585600110|160|0.613530739938246|0|26|273|-80.825175|43|35.152722|PREMIUM NOVELTIES|0.0|5|KLONDIKE HEATH BAR|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00075856011135|FROZEN NOVELTIES|FROZEN|-80.825175|1.4106654222506079|160|1
35.152722|1b8f506873e4c8d88d532186f7470b89c5a40614|3.65|2015-02-11 14:45:00|1.4094857484078087|1|7585600110|160|0.613530739938246|0|26|273|-80.825175|43|35.152722|PREMIUM NOVELTIES|0.0|5|KLONDIKE HEATH BAR|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00075856011135|FROZEN NOVELTIES|FROZEN|-80.825175|1.4106654222506079|160|1
35.152722|25844b372be444cc90d1d3ea82726aa8b3ff607a|7.99|2015-02-14 20:33:00|80.825044058860698|1|8190863007|160|35.170227534288045|0|29|9964|-80.826724|887|35.195689|NFS-S/PREM-PINOT NOIR|0.0|13|CONCANNON PINOT NOIR|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00081908630070|SUPER PREMIUM ($11-$14.99)|WINE|-80.825175|80.825184421307398|412|1
35.152722|e236cb5e20020bdf323b5cd8603342b31544a3a0|3.65|2015-01-29 19:29:00|1.4094857484078087|1|7585600110|160|0.613530739938246|0|26|273|-80.825175|43|35.152722|PREMIUM NOVELTIES|0.0|5|KLONDIKE HEATH BAR|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00075856011135|FROZEN NOVELTIES|FROZEN|-80.825175|1.4106654222506079|160|1
35.152722|9544da6fab1d66987ef159bc001703849ffdb5a9|2.39|2014-10-31 17:32:00|1.4094857484078087|1|7084781116|160|0.613530739938246|0|26|97|-80.825175|8|35.152722|ENERGY DRINKS|0.89|23|MONSTER ABSOLUTELY ZERO CAN|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00070847000037|CARBONATED BEVERAGES|BEVERAGE|-80.825175|1.4106654222506079|160|1
35.152722|e4490917c952b2660073c18262cc728828e1cadc|4.78|2014-09-13 21:44:00|1.4094857484078087|1|7084781116|160|0.613530739938246|0|26|97|-80.825175|8|35.152722|ENERGY DRINKS|0.0|23|MONSTER ABSOLUTELY ZERO CAN|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00070847000037|CARBONATED BEVERAGES|BEVERAGE|-80.825175|1.4106654222506079|160|2
35.152722|eb60c58f8fdb5f74c012312c0612bee799a8a7b4|10.99|2014-11-06 15:20:00|80.825044058860698|1|4740000126|160|35.170227534822438|0|29|3917|-80.80146|1075|35.17739|DISPOSABLE RAZOE-MEN|2.0|17|(FE) GIL FUSION DISPOSBL RZR|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00047400001268|SHAVING NEEDS/MEN HAIR|HBC|-80.825175|80.825182795370594|208|1
35.152722|3c60df4a4d3cd275323574729db9ab047632226e|4.39|2015-01-11 16:34:00|80.825044058860698|1|4400002796|160|35.170227534822438|0|29|90|-80.80146|13|35.17739|SNACK CRACKERS|1.39|1|TRISCUIT SWT POTATO RST ONION|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00044000031596|CRACKERS|G1 GROCERY|-80.825175|80.825182795370594|208|1
35.152722|2f81c85384ac926ea8740e1f4d8cac9bd94f404c|3.49|2014-10-24 16:30:00|80.825044058860698|1|4178001502|160|35.170227534617439|0|29|199|-80.806073|31|35.106477|DIPS & SALSAS|0.8|1|UTZ MILD SALSA|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00041780015020|SNACKS|G1 GROCERY|-80.825175|80.82518345614416|4|1
35.152722|acd8011010dda631a9af8bdebb186e984fa09e8e|3.99|2014-10-08 08:31:00|80.825044058860698|1|7127923100|160|35.170227491957206|0|29|555|-80.764523|64|35.341927|PACKAGED SALADS|0.0|4|F.E. BABY SPRING SALAD MIX|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00071279231006|FRESH PRODUCE|PRODUCE|-80.825175|80.825223022923083|220|1
35.152722|8e03e0c97217734aedb398387c5bccbcff6ae400|5.5|2014-12-21 08:41:00|1.4094857484078087|1|2800021010|160|0.613530739938246|0|26|16|-80.825175|3|35.152722|BAKING CHOCOLATE/CHIPS/MORSELS|0.0|1|NESTLE PREM.WHITE CHOC CHIP|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00028000210106|BAKING SUPPLIES|G1 GROCERY|-80.825175|1.4106654222506079|160|2
35.152722|94c089e455f79c73fe61f2819a5c43f31faa3010|5.55|2015-03-03 10:25:00|1.4094857484078087|1|3700006194|160|0.613530739938246|0|26|3527|-80.825175|1045|35.152722|HAIR CARE SHPOO-MED|0.56|17|H&S ITCHY SCALP SHAMPOO|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00037000473657|HAIR & SCALP CARE|HBC|-80.825175|1.4106654222506079|160|1
35.152722|2f57fa23928f8361f3f816e7fd7bd8d60cd08e15|11.99|2014-12-27 16:43:00|1.4094857484078087|1|2301286481|160|0.613530739938246|0|26|1477|-80.825175|485|35.152722|SUSHI HYBRID|0.0|6|"CHEF SAMPLER ""A"""|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00023012864811|SUSHI|DELI|-80.825175|1.4106654222506079|160|1
35.152722|4e8a92d6c68eef5c1d332af922937b1d9d980fbc|11.99|2014-11-12 21:08:00|80.825044058860698|1|8600300340|160|35.170227533599295|0|29|9939|-80.85753|885|35.116638|NFS POP PINOT NOIR|0.0|13|WOODBRIDGE PINOT NOIR 1.5L|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00086003003408|POPULAR (4-$7.99)|WINE|-80.825175|80.825186173210739|204|1
35.152722|23461353f4c87bfbca85cfc759da26ac2529e362|3.39|2014-12-12 09:32:00|80.825044058860698|1|2113150605|160|35.170227491957206|0|29|1279|-80.764523|48|35.341927|SINGLE SERVE FLAVOR|0.89|5|M CALLENDER PENNE GARLIC CHKN|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00021131800376|FROZEN MEALS|FROZEN|-80.825175|80.825223022923083|220|1
35.152722|b38f92e6497f12a9a79abd8692b143daa182a581|6.3|2014-11-30 12:21:00|1.4094857484078087|1|7203603083|160|0.613530739938246|0|26|30|-80.825175|4|35.152722|CARBONATED WATER|0.96|1|HT LEMON LIME SELTZER 12 PK|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00072036030849|BOTTLED WATER|G1 GROCERY|-80.825175|1.4106654222506079|160|2
35.152722|cef4a7760661748811d047d6288e9be1a3ba644d|3.69|2014-09-10 17:39:00|1.4094857484078087|1|7518500700|160|0.613530739938246|0|26|1030|-80.825175|162|35.152722|SLICED BREAD POTATO|0.0|7|MARTINS POTATO BREAD|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00075185007007|SLICED BREAD|COMMERCIAL BAKERY|-80.825175|1.4106654222506079|160|1
35.152722|c8ba9d230f6e3bfb32f4370bf7009ee2e8634cef|3.69|2015-03-03 12:30:00|1.4094857484078087|1|7518500700|160|0.613530739938246|0|26|1030|-80.825175|162|35.152722|SLICED BREAD POTATO|0.0|7|MARTINS POTATO BREAD|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00075185007007|SLICED BREAD|COMMERCIAL BAKERY|-80.825175|1.4106654222506079|160|1
35.152722|c13363c60f6bfb47e9ab29aad79fc2b86659a015|6.3|2015-02-14 18:11:00|1.4094857484078087|1|7203603083|160|0.613530739938246|0|26|30|-80.825175|4|35.152722|CARBONATED WATER|0.3|1|HT LEMON LIME SELTZER 12 PK|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00072036030849|BOTTLED WATER|G1 GROCERY|-80.825175|1.4106654222506079|160|2
35.152722|072bb471f3cc9eef2d773e1a7d77834a0bd1509d|19.99|2014-11-16 19:59:00|80.825044058860698|1|1820096715|160|35.17022753420661|0|29|455|-80.844274|82|35.204336|DOMESTIC PREMIUM 12PK&>|0.0|16|MICHELOB ULTRA 24PK CANS|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00018200967153|DOMESTIC BEER|BEER|-80.825175|80.825184645071957|61|1
35.152722|814bf0cbfde451fc33e73e0619b1f143657b3f37|7.98|2014-12-01 08:26:00|80.825044058860698|1|3400021303|160|35.170227491957206|0|29|46|-80.764523|7|35.341927|PKG CHOC|1.0|1|KIT KAT MINIATURES BAG 11 OZ|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00034000225392|CANDY|G1 GROCERY|-80.825175|80.825223022923083|220|2
35.152722|ce7792841cfc58e507fee11f94f8a751712b4dbe|3.99|2014-10-02 21:41:00|80.825044058860698|1|2500005542|160|35.170227534617439|0|29|335|-80.806073|56|35.106477|ORANGE JUICE-REGRIGERATED|0.99|3|SIMPLY ORANGE CALCIUM|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00025000055430|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.825175|80.82518345614416|4|1
35.152722|6edc037e09a0647f409de72d76e3458ebb445508|7.98|2014-09-15 13:50:00|1.4094857484078087|1|3338300005|160|0.613530739938246|0|26|500|-80.825175|64|35.152722|FRESH APPLES|0.0|4|RED DEL APPLE 3LB BAG|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00072036880116|FRESH PRODUCE|PRODUCE|-80.825175|1.4106654222506079|160|2
35.152722|b12a7e27dfcae6b44aa6037219b0831871202486|3.99|2014-09-10 16:56:00|80.825044058860698|1|3338300005|160|35.170227491957206|0|29|500|-80.764523|64|35.341927|FRESH APPLES|0.0|4|RED DEL APPLE 3LB BAG|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00072036880116|FRESH PRODUCE|PRODUCE|-80.825175|80.825223022923083|220|1
35.152722|e360b800681496e4139dfb0b1a91e0a82c6443e5|0.95|2014-10-03 12:52:00|80.825044058860698|1|61300871771|160|35.170227533599295|0|29|99|-80.85753|32|35.116638|LIQUID TEA|0.0|1|ARIZONA GINSENG TEA|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00613008715267|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.825175|80.825186173210739|204|1
35.152722|9f126295693ec504fb839e72c1077b238e41a26f|0.95|2014-10-01 09:54:00|80.825044058860698|1|61300871771|160|35.170227533599295|0|29|99|-80.85753|32|35.116638|LIQUID TEA|0.0|1|ARIZONA GINSENG TEA|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00613008715267|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.825175|80.825186173210739|204|1
35.152722|4b90a7376005070a721b2d62dccdaf48db471ee2|0.95|2014-11-10 09:49:00|80.825044058860698|1|61300871771|160|35.170227533599295|0|29|99|-80.85753|32|35.116638|LIQUID TEA|0.0|1|ARIZONA GINSENG TEA|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00613008715267|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.825175|80.825186173210739|204|1
35.152722|255de5b14991aec6c7370d4c71ab37ad750bee83|15.99|2015-02-14 23:30:00|1.4094857484078087|1|1820053349|160|0.613530739938246|0|26|455|-80.825175|82|35.152722|DOMESTIC PREMIUM 12PK&>|0.0|16|BUD LIGHT 24PK 12OZ BOTTLES|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00018200533495|DOMESTIC BEER|BEER|-80.825175|1.4106654222506079|160|1
35.152722|1fb9d7ce32d9b10f17d0896f9a48560a5dc9e99c|12.0|2014-10-01 10:27:00|80.825044058860698|1||160|35.170227533599295|0|29|511|-80.85753|64|35.116638|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00204770000004|FRESH PRODUCE|PRODUCE|-80.825175|80.825186173210739|204|6
35.152722|700ee59d8a59f6d8e30e651157bd4906d5ace09d|0.99|2014-10-12 06:49:00|80.825044058860698|1|7203698116|160|35.170227525044652|0|29|31|-80.8062|4|35.037115|NON CARBONATED WATER|0.24|1|HT SMPLY ACAI/BLU/POM VIT WATR|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00072036981189|BOTTLED WATER|G1 GROCERY|-80.825175|80.825198936651461|27|1
35.152722|9ba380a8d7e57d0f0680426bec1d97c61a680fac|1.99|2014-09-14 18:25:00|1.4094857484078087|1|7203688083|160|0.613530739938246|0|26|526|-80.825175|64|35.152722|FRESH MUSHROOMS|0.2|4|HT WHITE MUSHROOMS, 8 OZ WHOLE|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00072036880833|FRESH PRODUCE|PRODUCE|-80.825175|1.4106654222506079|160|1
35.152722|4c0e7859dc6e10479a66c273232ff4589f84e890|3.39|2014-12-19 09:47:00|80.825044058860698|1|2113150605|160|35.170227491957206|0|29|1279|-80.764523|48|35.341927|SINGLE SERVE FLAVOR|0.89|5|M CALLENDER STUFF RIGATONI CKN|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00021131507305|FROZEN MEALS|FROZEN|-80.825175|80.825223022923083|220|1
35.152722|144bff2b6f65c9a1686bc31321ec0644c83e376f|0.99|2014-12-03 09:55:00|80.825044058860698|1|7203695306|160|35.170227533599295|0|29|1895|-80.85753|450|35.116638|TEA|0.0|6|FFM DIET TEA W/SPLENDA|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00072036018892|BEVERAGES|DELI|-80.825175|80.825186173210739|204|1
35.152722|c5b87b0d2c2c238e7b9f56523ac0e6a6318dad6e|5.39|2014-11-16 22:24:00|1.4094857484078087|1|3450015193|160|0.613530739938246|0|26|312|-80.825175|51|35.152722|BUTTER|0.0|3|LOL W/OLV OIL SEA SALT HF STKS|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00034500151931|BUTTER & MARGARINE|DAIRY|-80.825175|1.4106654222506079|160|1
35.152722|067c0d69bad824d07851987a3226f2965005a5d4|14.91|2014-09-19 23:08:00|1.4094857484078087|1|7203688105|160|0.613530739938246|0|26|500|-80.825175|64|35.152722|FRESH APPLES|0.0|4|HT RED DEL 5LB BAG|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00072036881052|FRESH PRODUCE|PRODUCE|-80.825175|1.4106654222506079|160|3
35.152722|4239779957e00e2598cfea9931f60a8a2c7f7851|23.96|2015-01-31 18:41:00|1.4094857484078087|1|7203688105|160|0.613530739938246|0|26|500|-80.825175|64|35.152722|FRESH APPLES|0.0|4|HT RED DEL 5LB BAG|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00072036881052|FRESH PRODUCE|PRODUCE|-80.825175|1.4106654222506079|160|4
35.152722|b30ee90f0e7dbc2a81602c09c69c9d5cfda6d09c|24.85|2014-09-27 00:37:00|1.4094857484078087|1|7203688105|160|0.613530739938246|0|26|500|-80.825175|64|35.152722|FRESH APPLES|0.0|4|HT RED DEL 5LB BAG|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00072036881052|FRESH PRODUCE|PRODUCE|-80.825175|1.4106654222506079|160|5
35.152722|429c6b9d5114b7bb03f1e082ce6a6d81016e7f41|2.39|2014-09-09 23:52:00|1.4094857484078087|1|7084781116|160|0.613530739938246|0|26|97|-80.825175|8|35.152722|ENERGY DRINKS|0.0|23|MONSTER LOW CARB ENRGY CAN|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00070847811268|CARBONATED BEVERAGES|BEVERAGE|-80.825175|1.4106654222506079|160|1
35.152722|930c4d027bc86e821026cf8a06433f1e8f4afd92|12.99|2015-02-13 23:25:00|80.825044058860698|1|7199009554|160|35.170227530872587|0|29|458|-80.810056|82|35.219587|CRAFT BEER|0.0|16|BLUE MOON VARIETY 12PK|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00071990095543|DOMESTIC BEER|BEER|-80.825175|80.825191360781005|401|1
35.152722|f414a914f5eeec3e11c238db2ca613727c63df5b|6.49|2014-11-01 21:33:00|80.825044058860698|1|2301200005|160|35.170227534617439|0|29|1479|-80.806073|485|35.106477|SUSHI HYBRID SPECIALTY|0.0|6|TROPICAL SALAD|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00023012000059|SUSHI|DELI|-80.825175|80.82518345614416|4|1
35.152722|d15586b78b09b3eb7a4020f9c2325611450bc3ea|16.98|2015-02-04 13:05:00|1.4094857484078087|1|84105802507|160|0.613530739938246|0|26|3917|-80.825175|1075|35.152722|DISPOSABLE RAZOE-MEN|0.0|17|SCHICK SLM TWN SENSITVE GRIP|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00841058025078|SHAVING NEEDS/MEN HAIR|HBC|-80.825175|1.4106654222506079|160|2
35.152722|3cdb632c81c313f30ea3be79820e5da132e1b236|7.99|2015-02-28 21:46:00|80.825044058860698|1|2210000170|160|35.1702275358397|0|29|454|-80.85013|82|35.175855|DOMESTIC ECONOMY 12PK&>|0.0|16|PABST 12PK 12OZ CAN|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00022100001701|DOMESTIC BEER|BEER|-80.825175|80.825177734975583|218|1
35.152722|545496b72a71b55d56730875e305bc1e204269cb|23.97|2015-01-16 12:17:00|80.825044058860698|1|3600025830|160|35.170227491957206|0|29|424|-80.764523|72|35.341927|NFS-FACIAL TISSUE|0.0|1|KLEENEX LOTION UPRIGHT 4PK|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00036000258325|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.825175|80.825223022923083|220|3
35.152722|03aa459b720046df0973dd7d04ba4b2000bc0d2c|14.99|2015-02-01 19:10:00|1.4094857484078087|1|946808164|160|0.613530739938246|0|26|458|-80.825175|82|35.152722|CRAFT BEER|0.0|16|SARANAC TRAIL MIX 12PK BTL|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00009468081644|DOMESTIC BEER|BEER|-80.825175|1.4106654222506079|160|1
35.152722|13166e378f8a0d77ba90d826cd47c630b69c1c2f|3.49|2014-10-10 16:36:00|1.4094857484078087|1|4850002115|160|0.613530739938246|0|26|338|-80.825175|56|35.152722|OTHER FRUIT JUICES|0.99|3|DOLE BLENDS-ORANGE STWBRY BANA|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00048500021118|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.825175|1.4106654222506079|160|1
35.152722|662b18ea4309ae1c5721ba83a125d6c6458ec9bb|0.99|2014-09-11 09:50:00|80.825044058860698|1|7203695306|160|35.170227533599295|0|29|1895|-80.85753|450|35.116638|TEA|0.0|6|FFM SWEET TEA|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00072036953063|BEVERAGES|DELI|-80.825175|80.825186173210739|204|1
35.152722|ec23dfa25104204fe55d1b5fd03f752f1f10c5a8|0.99|2014-10-07 09:47:00|80.825044058860698|1|7203695306|160|35.170227533599295|0|29|1895|-80.85753|450|35.116638|TEA|0.0|6|FFM SWEET TEA|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00072036953063|BEVERAGES|DELI|-80.825175|80.825186173210739|204|1
35.152722|cfed5f660b4fd5364a42b9153707964a9fdacecd|7.99|2015-01-18 19:36:00|1.4094857484078087|1|8600309193|160|0.613530739938246|0|26|9952|-80.825175|886|35.152722|NFS-PREM-PINOT NOIR|0.0|13|R. MONDAVI P.S. PINOT NOIR|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00086003091931|PREMIUM ($8-$10.99)|WINE|-80.825175|1.4106654222506079|160|1
35.152722|6bf6a13843a61258f625869430dce22857fc1fb3|6.76|2014-12-20 14:19:00|80.825044058860698|1|4430012171|160|35.170227534822438|0|29|1216|-80.80146|273|35.17739|ASIAN RICE/NOODLES|1.76|1|LACHOY NOODLES CHOW MEIN|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00044300121713|ASIAN PREP. FOODS|G1 GROCERY|-80.825175|80.825182795370594|208|4
35.152722|bb738a4d0e70768712323f54d71d6c43cbc83cc4|18.99|2014-10-26 21:36:00|1.4094857484078087|1|3700088207|160|0.613530739938246|0|26|426|-80.825175|72|35.152722|NFS-PAPER TOWELS|0.0|1|BOUNTY TOWEL 12 WHITE|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|0.61471665291522548|00037000882077|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.825175|1.4106654222506079|160|1
35.152722|409c8fad53688edd715e0784d64cc87627c23302|14.99|2014-11-23 16:52:00|80.825044058860698|1|946831513|160|35.1702275358397|0|29|459|-80.85013|83|35.175855|IMPORT BEER|0.0|16|SARANAC TRAIL MIX 13PK|2e429b227264060e0e932e4456acadfe0289e843|1.2095902620343821|35.157881615307893|00009468315138|IMPORT BEER|BEER|-80.825175|80.825177734975583|218|1
35.082768|3e3b4d4cba72925c868d069d2837b46540292190|3.85|2015-02-22 15:46:00|1.4091206135396188|2|4812127620|147|0.6123098123133061|0|47|1037|-80.732725|164|35.082768|ENGLISH MUFFINS|0.0|7|THOMAS LITE MULTIGRAIN EM PP|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|0.61242566243833529|00048121276201|BREAKFAST|COMMERCIAL BAKERY|-80.732725|1.409051865357139|147|1
35.082768|88f908270abfdef97541e8d7ca23451fc512cf07|6.98|2014-12-01 18:34:00|80.732732175546019|2|4812127620|147|35.104380197732347|0|35|1037|-80.771677|164|35.066546|ENGLISH MUFFINS|1.74|7|THOMAS LITE MULTIGRAIN EM PP|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00048121276201|BREAKFAST|COMMERCIAL BAKERY|-80.732725|80.732734120956124|45|2
35.082768|515adc05b397e368c57ef9a4b2acb34b94ef708f|6.98|2014-11-10 18:34:00|80.732732175546019|2|4812127620|147|35.104380197732347|0|35|1037|-80.771677|164|35.066546|ENGLISH MUFFINS|1.74|7|THOMAS LITE MULTIGRAIN EM PP|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00048121276201|BREAKFAST|COMMERCIAL BAKERY|-80.732725|80.732734120956124|45|2
35.082768|a6f4d89ef033de40a5355c7d8c2ce6176b953061|3.85|2015-02-09 18:55:00|80.732732175546019|2|4812127620|147|35.104380197732347|0|35|1037|-80.771677|164|35.066546|ENGLISH MUFFINS|0.0|7|THOMAS LITE MULTIGRAIN EM PP|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00048121276201|BREAKFAST|COMMERCIAL BAKERY|-80.732725|80.732734120956124|45|1
35.082768|121b47af8507ed97e981a7f1bb61d2153865fb2f|6.38|2014-12-28 18:22:00|80.732732175546019|2|4227200504|147|35.104380197732347|0|35|1201|-80.771677|33|35.066546|RTS CANNED|0.0|1|AMY'S ORG SP BLACK BEAN VEG|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00042272005048|SOUP|G1 GROCERY|-80.732725|80.732734120956124|45|2
35.082768|a6ccf24531229f6c91303ebbe1c1f420de5aafa9|6.38|2014-10-04 19:48:00|80.732732175546019|2|4227200504|147|35.10438019902076|0|35|1201|-80.7007|33|35.06858|RTS CANNED|0.0|1|AMY'S ORG SP BLACK BEAN VEG|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00042272005048|SOUP|G1 GROCERY|-80.732725|80.732725074728819|273|2
35.082768|396be8f376acf764a226967e4457897ee610fd6a|6.38|2014-11-23 15:30:00|80.732732175546019|2|4227200504|147|35.10438019902076|0|35|1201|-80.7007|33|35.06858|RTS CANNED|0.0|1|AMY'S ORG SP BLACK BEAN VEG|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00042272005048|SOUP|G1 GROCERY|-80.732725|80.732725074728819|273|2
35.082768|7215247c03d12f67b5b6e10b7aabb0b53b418585|5.98|2015-03-03 18:59:00|80.732732175546019|2|4227200504|147|35.104380197732347|0|35|1201|-80.771677|33|35.066546|RTS CANNED|0.0|1|AMY'S ORG SP BLACK BEAN VEG|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00042272005048|SOUP|G1 GROCERY|-80.732725|80.732734120956124|45|2
35.082768|0b88c4c77ee58f969362f976c7082e61235bd6d5|5.98|2015-02-16 18:07:00|80.732732175546019|2|4227200504|147|35.104380197732347|0|35|1201|-80.771677|33|35.066546|RTS CANNED|0.0|1|AMY'S ORG SP BLACK BEAN VEG|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00042272005048|SOUP|G1 GROCERY|-80.732725|80.732734120956124|45|2
35.082768|3d1e0e90f68ce25f58f3fc0b6fe5ee84727748fd|5.98|2015-01-24 19:46:00|1.4091206135396188|2|4227200504|147|0.6123098123133061|0|47|1201|-80.732725|33|35.082768|RTS CANNED|0.0|1|AMY'S ORG SP BLACK BEAN VEG|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|0.61242566243833529|00042272005048|SOUP|G1 GROCERY|-80.732725|1.409051865357139|147|2
35.082768|cfd57e2c3d4f4bd51ddfd7f8abfd2b7f6a21912f|6.38|2014-10-12 19:34:00|80.732732175546019|2|4227200504|147|35.104380197732347|0|35|1201|-80.771677|33|35.066546|RTS CANNED|0.0|1|AMY'S ORG SP BLACK BEAN VEG|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00042272005048|SOUP|G1 GROCERY|-80.732725|80.732734120956124|45|2
35.082768|a86329c070280c421127d206328a58cde6335f90|5.98|2015-02-25 19:25:00|80.732732175546019|2|4227200504|147|35.104380197732347|0|35|1201|-80.771677|33|35.066546|RTS CANNED|0.0|1|AMY'S ORG SP BLACK BEAN VEG|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00042272005048|SOUP|G1 GROCERY|-80.732725|80.732734120956124|45|2
35.082768|731443428539df71ddbe73e682739e809ec0a2aa|6.38|2015-01-05 18:40:00|80.732732175546019|2|4227200504|147|35.104380197732347|0|35|1201|-80.771677|33|35.066546|RTS CANNED|0.0|1|AMY'S ORG SP BLACK BEAN VEG|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00042272005048|SOUP|G1 GROCERY|-80.732725|80.732734120956124|45|2
35.082768|9b66d54095a2f7b28579a6f0e1fb9fde6cd1d5eb|1.59|2015-03-08 17:05:00|80.732732175546019|2|4650073332|147|35.104380197732347|0|35|393|-80.771677|68|35.066546|NFS-AIR FRESHENERS|0.0|1|GLADE AEROSOL LAVENDR VANILLA|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00046500733345|FRESHENERS/DEODORIZERS|G1 GROCERY|-80.732725|80.732734120956124|45|1
35.082768|d8486c8e6edd96b0a41a45010fa6657984f22b88|3.89|2014-12-20 17:20:00|1.4091206135396188|2|2100012277|147|0.6123098123133061|0|47|320|-80.732725|53|35.082768|COTTAGE CHEESE|0.0|3|BREAKSTONE 2% COTTAGE CHEESE|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|0.61242566243833529|00021000123544|CULTURES|DAIRY|-80.732725|1.409051865357139|147|1
35.082768|7f718eb917327ddd2b17dbdbe175c98b5f93c15d|7.78|2014-10-11 12:19:00|80.732732175546019|2|2200001530|147|35.104380197732347|0|35|45|-80.771677|7|35.066546|PEG GUM|1.0|1|ORBIT SPEARMINT BOTTLE|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00022000015297|CANDY|G1 GROCERY|-80.732725|80.732734120956124|45|2
35.082768|bd8eb1eae6f90e011062c564bc551c0c14cf06c0|9.99|2014-10-17 18:55:00|1.4091206135396188|2|7103800044|147|0.6123098123133061|0|47|66|-80.732725|10|35.082768|GROUND CAN|2.0|1|CHOCK FULL O'NUTS GOURM ROAST|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|0.61242566243833529|00071038011740|COFFEE|G1 GROCERY|-80.732725|1.409051865357139|147|1
35.082768|635751140adaf71cb458d77d88045fa315855a0e|7.98|2014-11-15 14:42:00|1.4091206135396188|2|20405400000|147|0.6123098123133061|0|47|504|-80.732725|64|35.082768|FRESH BERRIES|1.99|4|RED RASPBERRIES 6 OZ|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|0.61242566243833529|00715756100019|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|2
35.082768|500b40c33e5d50562593da6661e42cf6a7d28472|3.99|2014-11-03 18:25:00|1.4091206135396188|2|20405400000|147|0.6123098123133061|0|47|504|-80.732725|64|35.082768|FRESH BERRIES|1.49|4|RED RASPBERRIES 6 OZ|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|0.61242566243833529|00715756100019|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|1
35.082768|1eb251cb3d00611bad27d77e5641d7fd9e0b6c53|3.4|2014-09-13 16:55:00|1.4091206135396188|2||147|0.6123098123133061|0|47|501|-80.732725|64|35.082768|FRESH PEARS|0.51|4|BARTLETT PEARS|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|0.61242566243833529|00204409000009|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|1
35.082768|78ea09db3b6e398b2f6c3883b590bfffd902403e|6.99|2014-10-19 17:13:00|80.732732175546019|2|7027710518|147|35.104380197732347|0|35|2020|-80.771677|505|35.066546|CHEESE SPECIALTIES|0.0|6|ATHENOS FETA TRADITIONAL CHUNK|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00070277105180|SPECIALTY CHEESE|DELI|-80.732725|80.732734120956124|45|1
35.082768|053602d77fd06f9b998a97d04df215b94095ebbf|2.19|2014-11-17 19:00:00|1.4091206135396188|2|7203608066|147|0.6123098123133061|0|47|1220|-80.732725|275|35.082768|PASTA SC PREMIUM|0.0|1|HTO PASTA SC TOM BASIL|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|0.61242566243833529|00072036080660|PASTA SAUCES|G1 GROCERY|-80.732725|1.409051865357139|147|1
35.082768|5234fe9660f76f195136ad897132e45e54857c1c|16.02|2015-02-11 11:33:00|80.732732175546019|2|20436500000|147|35.104380194112174|0|35|562|-80.80146|64|35.17739|FRESH CUT FRUIT|0.0|4|VEG TRAY MISC. BY POUND|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00204365000006|FRESH PRODUCE|PRODUCE|-80.732725|80.732742802445514|208|1
35.082768|41c0afc9951a579368f3681f82b58fc9e6580537|7.7|2015-01-16 22:48:00|1.4091206135396188|2|4812127620|147|0.6123098123133061|0|47|1037|-80.732725|164|35.082768|ENGLISH MUFFINS|1.93|7|THOMAS 100% WHEAT ENG MUFN PP|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|0.61242566243833529|00048121184070|BREAKFAST|COMMERCIAL BAKERY|-80.732725|1.409051865357139|147|2
35.082768|fead686881fe007e1da8b2d58e74461db1776d1e|4.99|2015-01-17 15:09:00|1.4091206135396188|2|61611202795|147|0.6123098123133061|0|47|581|-80.732725|136|35.082768|FRESH SALSA|0.0|4|WHOLLY GUACAMOL CLASSIC 16OZ|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|0.61242566243833529|00616112027950|OTHER MERCHANDISE|PRODUCE|-80.732725|1.409051865357139|147|1
35.082768|22e6c24e0b908943fddf93a9bdd37c5ee4a9c9a6|3.49|2015-02-08 18:23:00|80.732732175546019|2|3800001611|147|35.104380197732347|0|35|61|-80.771677|9|35.066546|RTE CEREAL ADULT|0.0|1|KELLOGG SPECIAL K 12 OZ BOX|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00038000016110|CEREAL|G1 GROCERY|-80.732725|80.732734120956124|45|1
35.082768|9f38c115fc7765aa8ed97dcc3bc812cb1af96330|3.39|2015-01-05 15:41:00|80.732732175546019|2|1862770327|147|35.104380197732347|0|35|61|-80.771677|9|35.066546|RTE CEREAL ADULT|0.0|1|KASHI GO LEAN CRUNCH|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00018627703273|CEREAL|G1 GROCERY|-80.732725|80.732734120956124|45|1
35.082768|f62ac4e0b3ea82c05f563c69303b1f9f3e4d4321|4.99|2015-02-06 17:12:00|1.4091206135396188|2|2531711100|147|0.6123098123133061|0|47|845|-80.732725|100|35.082768|NATURAL/ORGANIC BACON|0.0|19|APPLEGATE GOOD MORNING BACON|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|0.61242566243833529|00025317111003|BACON|CASE READY MEATS|-80.732725|1.409051865357139|147|1
35.082768|effde319eeda401dd18f9b9ca6cfcc52152dfba2|2.5|2014-12-05 18:00:00|80.732732175546019|2|7203652034|147|35.10438019902076|0|35|74|-80.7007|9|35.06858|RTE CEREAL ALL FAMILY|0.53|1|HT CER CORN FLAKES|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00072036520340|CEREAL|G1 GROCERY|-80.732725|80.732725074728819|273|1
35.082768|4fa581f58c4edae48244cea01ffab288321a84c9|2.5|2015-02-24 16:28:00|80.732732175546019|2|7203652034|147|35.10438019902076|0|35|74|-80.7007|9|35.06858|RTE CEREAL ALL FAMILY|0.53|1|HT CER CORN FLAKES|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00072036520340|CEREAL|G1 GROCERY|-80.732725|80.732725074728819|273|1
35.082768|84988f9ae544f00ddc844bd31e4836c47df4dfc2|2.69|2015-02-03 16:38:00|80.732732175546019|2|88491200620|147|35.104380197732347|0|35|74|-80.771677|9|35.066546|RTE CEREAL ALL FAMILY|0.0|1|POST HONEY GRAHAM OH'S|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00884912006202|CEREAL|G1 GROCERY|-80.732725|80.732734120956124|45|1
35.082768|d6057b565f40c4cee71758dce677313bf9d2fcee|4.89|2015-02-12 16:19:00|80.732732175546019|2|1600027529|147|35.104380197732347|0|35|61|-80.771677|9|35.066546|RTE CEREAL ADULT|0.0|1|GM RAISIN NUT BRAN|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00016000275294|CEREAL|G1 GROCERY|-80.732725|80.732734120956124|45|1
35.082768|a30bec5a2c0af27ee8b7a1314eadf3e1f16489bb|4.89|2015-02-21 12:11:00|80.732732175546019|2|1600027529|147|35.104380197732347|0|35|61|-80.771677|9|35.066546|RTE CEREAL ADULT|0.0|1|GM RAISIN NUT BRAN|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00016000275294|CEREAL|G1 GROCERY|-80.732725|80.732734120956124|45|1
35.082768|b79c960bb5d70a28ebc993971c646d714ee42309|4.29|2015-01-23 18:59:00|1.4091206135396188|2|3000006119|147|0.6123098123133061|0|47|74|-80.732725|9|35.082768|RTE CEREAL ALL FAMILY|0.0|1|QUAKER ORIGINAL LIFE|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|0.61242566243833529|00030000061190|CEREAL|G1 GROCERY|-80.732725|1.409051865357139|147|1
35.082768|a281b4e45e84f3a3062b59da77dde077fe745e63|4.29|2015-02-16 10:08:00|80.732732175546019|2|3000006119|147|35.104380197732347|0|35|74|-80.771677|9|35.066546|RTE CEREAL ALL FAMILY|0.0|1|QUAKER ORIGINAL LIFE|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00030000061190|CEREAL|G1 GROCERY|-80.732725|80.732734120956124|45|1
35.082768|5460075ddeeec635cf7a1603127b8679d23d5291|3.67|2014-12-14 19:32:00|80.732732175546019|2|7203655019|147|35.104380197732347|0|35|332|-80.771677|52|35.066546|STRING/SNACK|0.0|3|HT LIGHT STRING CHEESE|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00072036705136|CHEESE|DAIRY|-80.732725|80.732734120956124|45|1
35.082768|e13abc0ce92457e3b100107f0e86cf0b84fd011d|3.99|2014-10-01 18:27:00|80.732732175546019|2|7203663995|147|35.104380197732347|0|35|342|-80.771677|57|35.066546|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00072036631282|MILK|DAIRY|-80.732725|80.732734120956124|45|1
35.082768|511fdec5e012032a56a4b29ec0a77d1e3332d264|3.49|2015-02-19 21:00:00|80.732732175546019|2|7203663995|147|35.104380197732347|0|35|342|-80.771677|57|35.066546|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00072036631282|MILK|DAIRY|-80.732725|80.732734120956124|45|1
35.082768|e9c200e4939bea54a8843fb515faffbd65912a1d|3.99|2014-12-09 12:17:00|80.732732175546019|2|7203663995|147|35.104380196506291|0|35|342|-80.770346|57|35.052812|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00072036631282|MILK|DAIRY|-80.732725|80.732737741718609|40|1
35.082768|761048034c89c3e93aa7d0a5d666ce6ff78b5330|3.99|2014-12-19 20:34:00|80.732732175546019|2|7203663995|147|35.104380197732347|0|35|342|-80.771677|57|35.066546|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00072036631282|MILK|DAIRY|-80.732725|80.732734120956124|45|1
35.082768|c49d8bc9aabebbbacd1bf3455282277613da46cf|3.95|2014-12-15 13:14:00|80.732732175546019|2|7203663995|147|35.104380197732347|0|35|342|-80.771677|57|35.066546|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00072036631282|MILK|DAIRY|-80.732725|80.732734120956124|45|1
35.082768|05dce9343ad3e009ab425a76f6403540da0520c6|3.99|2014-10-03 18:35:00|80.732732175546019|2|7203663995|147|35.104380197732347|0|35|342|-80.771677|57|35.066546|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00072036631282|MILK|DAIRY|-80.732725|80.732734120956124|45|1
35.082768|dd069c69c89bc38062610c16edc52cfa0558c085|3.99|2014-09-16 19:07:00|80.732732175546019|2|7203663995|147|35.104380197732347|0|35|342|-80.771677|57|35.066546|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00072036631282|MILK|DAIRY|-80.732725|80.732734120956124|45|1
35.082768|fd3c64cf29f8f378a90d4bac9da36db22b9bb013|3.99|2014-11-29 18:11:00|1.4091206135396188|2|7203663995|147|0.6123098123133061|0|47|342|-80.732725|57|35.082768|FRESH MILK|1.52|3|HARRIS TEETER FF SKIM MILK|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|0.61242566243833529|00072036631282|MILK|DAIRY|-80.732725|1.409051865357139|147|1
35.082768|96851560cc9311ea87b794266efc81668721e147|3.99|2015-02-24 12:03:00|80.732732175546019|2|4740064972|147|35.104380197982927|0|35|3941|-80.825175|1075|35.152722|SHAVING CREAM MEN-GEL|1.0|17|MACH3 GEL SHAV PREP EXT CMFRT|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00047400650046|SHAVING NEEDS/MEN HAIR|HBC|-80.732725|80.732733186123582|160|1
35.082768|e939365d0e8342fbb1021f3758f5a5d2d40faa43|1.99|2015-02-13 18:21:00|80.732732175546019|2|1130010497|147|35.104380197732347|0|35|727|-80.771677|7|35.066546|SEASONAL CANDY-SINGLE FAC|0.74|1|I/O(V15)BRACH SM CONV HEARTS|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00011300104978|CANDY|G1 GROCERY|-80.732725|80.732734120956124|45|1
35.082768|e84eb04304970e3c07391e20582d232e58b44976|6.43|2014-10-13 15:48:00|80.732732175546019|2||147|35.104380197732347|0|35|503|-80.771677|64|35.066546|FRESH GRAPES|3.23|4|RED GRAPES, SEEDLESS|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00204635000002|FRESH PRODUCE|PRODUCE|-80.732725|80.732734120956124|45|1
35.082768|a74e492fb56a8b296fd2f379d25efaa859c657f1|2.67|2014-09-23 13:11:00|80.732732175546019|2|7203670794|147|35.104380197982927|0|35|388|-80.825175|66|35.152722|NFS-DISHWASH PWDR/LIQUID|0.0|1|YH DISHWASHER RINSE AID|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00072036707949|DETERGENTS|G1 GROCERY|-80.732725|80.732733186123582|160|1
35.082768|53bc28fc84697e12cd24a7c3e2420abfd339dbbd|5.57|2014-10-02 19:42:00|80.732732175546019|2|7203698580|147|35.104380196506291|0|35|66|-80.770346|10|35.052812|GROUND CAN|0.0|1|HT CLASSIC  ROAST COFFEE CAN|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00072036985804|COFFEE|G1 GROCERY|-80.732725|80.732737741718609|40|1
35.082768|c575dae5a4bd728cf539ee9bae9fb3dcaf756852|4.69|2014-09-20 15:36:00|80.732732175546019|2|7756712130|147|35.104380197732347|0|35|251|-80.771677|43|35.066546|NON-DAIRY NOVELTIES|0.0|5|POPSICLE SF ORANGE/CHRY/GRAPE|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00077567022950|FROZEN NOVELTIES|FROZEN|-80.732725|80.732734120956124|45|1
35.082768|9f71bd8f279f606a83437e91d8cb209295ebd575|4.9|2014-12-06 14:11:00|80.732732175546019|2|5100013279|147|35.104380197732347|0|35|214|-80.771677|33|35.066546|BROTH|0.0|1|SWANSON BROTH LOW SODIUM BEEF|3091f82159b99f0be79187a7ca0f8b7b2e4983a0|1.4933507607483785|35.101032182271901|00051000142962|SOUP|G1 GROCERY|-80.732725|80.732734120956124|45|2
35.333742|a85060bd4c9a50b16f7c0cfb190ae54b3b630972|3.49|2014-09-13 16:39:00|1.4102725052409182|4|1410007712|472|0.6166901349502063|0|1|1253|-80.814133|12|35.333742|ALL OTHER COOKIES|0.0|1|PF CRISPY COOKIES TAHOE|31f7e97b17f1a12abf0b342ce8fce3986c1ae494|1.3324475206560855|0.61833652052202714|00014100075226|COOKIES|G1 GROCERY|-80.814133|1.4104727029946025|472|1
35.333742|6faaefc6bf4573511a5d9d5db7131a5780bfb0af|5.99|2015-01-07 17:41:00|80.780380710856576|4|8500001581|472|35.353025560413023|0|48|9943|-80.764523|885|35.341927|NFS POP RIESLING|0.0|13|BAREFOOT RIESLING|31f7e97b17f1a12abf0b342ce8fce3986c1ae494|1.3324475206560855|35.351085445956379|00085000015810|POPULAR (4-$7.99)|WINE|-80.814133|80.814140341324034|220|1
35.667941|57b6a42ba8e7fba2e661b42074e2c7e4045ef126|2.89|2015-03-08 16:25:00|1.4057311447477159|3|7203655029|178|0.6225230078570788|0|52|331|-80.497332|52|35.667941|NATURAL SLICED|0.92|3|HT SWISS 2% SLICES CHEESE|32561fbb6668f5ad61b499570320235161445336|4.58838341412873|0.6209993146566879|00072036983954|CHEESE|DAIRY|-80.497332|1.4049434824709919|178|1
35.667941|1b338960be15fa366fa131973af2b02acff9c841|3.39|2015-02-18 19:21:00|1.4057311447477159|3|3800031829|178|0.6225230078570788|0|52|74|-80.497332|9|35.667941|RTE CEREAL ALL FAMILY|0.89|1|KELL MIN WH LIL BITES ORIG|32561fbb6668f5ad61b499570320235161445336|4.58838341412873|0.6209993146566879|00038000596827|CEREAL|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|f8a8cc6c0b34d6d0173abf1056c5db8752076d9e|5.78|2015-02-28 20:18:00|80.497482303704658|3|3760007060|178|35.734345108575518|0|6|714|-80.605588|274|35.43259|MICROWAVE MEALS|0.89|1|DINTY MOORE CMPL BEEF STEW|32561fbb6668f5ad61b499570320235161445336|4.58838341412873|35.699188602026126|00037600070607|PREP FOODS DINNERS|G1 GROCERY|-80.497332|80.497572660638042|202|2
35.667941|bb4c4b6a43daa07c3f834ce91e24c0c2bd1a912e|3.79|2015-02-24 16:47:00|1.4057311447477159|3|7020055044|178|0.6225230078570788|0|52|580|-80.497332|136|35.667941|OTHER MERCH DRESSINGS|0.0|4|MARZ SIMPLY CAESAR DRESSING|32561fbb6668f5ad61b499570320235161445336|4.58838341412873|0.6209993146566879|00070200550469|OTHER MERCHANDISE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|3bfa51ae591936ff3ccbe78a6128b70cc10492dd|6.7|2015-02-24 16:41:00|1.4057311447477159|3|3700022205|178|0.6225230078570788|0|52|725|-80.497332|66|35.667941|NFS-DISHWASHING LIQUID|1.35|1|DAWN LIQ DISH ANTIBAC APPLE BL|32561fbb6668f5ad61b499570320235161445336|4.58838341412873|0.6209993146566879|00037000222026|DETERGENTS|G1 GROCERY|-80.497332|1.4049434824709919|178|2
35.667941|197dc9392a2b001c45b711b48f50017055437fcd|7.1|2015-02-19 18:51:00|1.4057311447477159|3|3800039125|178|0.6225230078570788|0|52|74|-80.497332|9|35.667941|RTE CEREAL ALL FAMILY|1.75|1|KELLOGG RICE KRISPIES 9|32561fbb6668f5ad61b499570320235161445336|4.58838341412873|0.6209993146566879|00038000318443|CEREAL|G1 GROCERY|-80.497332|1.4049434824709919|178|2
35.667941|9397966d285b4acd4cc53535def6be54ddb1cb95|3.29|2015-03-08 16:31:00|1.4057311447477159|3|78052632501|178|0.6225230078570788|0|52|1279|-80.497332|48|35.667941|SINGLE SERVE FLAVOR|0.97|5|CP 5 PIECES SHRIMP WONTON|32561fbb6668f5ad61b499570320235161445336|4.58838341412873|0.6209993146566879|00780526325015|FROZEN MEALS|FROZEN|-80.497332|1.4049434824709919|178|1
35.667941|a17651ba5bc639a048a1b2c678e7fd22037cd40d|1.39|2015-01-24 11:36:00|1.4057311447477159|3|5210076069|178|0.6225230078570788|0|52|80|-80.497332|34|35.667941|SEASONING PACKETS|0.39|1|MC G M BAJA CITRUS MARINADE|32561fbb6668f5ad61b499570320235161445336|4.58838341412873|0.6209993146566879|00052100351889|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|c744d8c83b2b14ed7d7b52538f0e399cfca46ddc|1.8|2015-02-19 19:02:00|1.4057311447477159|3|1862703000|178|0.6225230078570788|0|52|42|-80.497332|6|35.667941|GRANOLA/YOGURT BARS|0.0|1|KASHI BAR CHWY CHERRY DK CHOC|32561fbb6668f5ad61b499570320235161445336|4.58838341412873|0.6209993146566879|00018627030034|BREAKFAST FOODS|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.585842|930df6038cfc6a195560aa9ae9261e0e9bd4568e|4.0|2014-09-24 06:23:00|80.891462859624312|4|84115200732|99|35.65765599504018|0|45|1165|-80.764523|87|35.341927|NFS-FRESH CONSUMER BUNCH|0.0|9|BUNCH- 3/$12 DAISY BUNCHES|369558d4159423fb1830455f1367010032eb09eb|4.962183813555141|35.636605227883024|00841152007321|FLORAL|FLORAL|-80.875654|80.875832959396263|220|1
35.585842|675caf240616f212bb9f3f43a169a7b29caf2a4c|3.99|2014-12-31 18:50:00|80.891462859624312|4|4450097650|99|35.65765599504018|0|45|840|-80.764523|102|35.341927|TUBS|0.0|19|HF THIN SMOKED HAM|369558d4159423fb1830455f1367010032eb09eb|4.962183813555141|35.636605227883024|00044500976496|LUNCHMEATS|CASE READY MEATS|-80.875654|80.875832959396263|220|1
35.204336|72f32df0648e3143daa3835fba80a5220e288d62|4.99|2014-12-16 14:51:00|80.828402574597021|4|7203688143|61|35.214435120733839|0|8|561|-80.80146|64|35.17739|FR PROD ORGANIC PRODUCE|0.0|4|ORG HT SPRING MIX 11 OZ|38847650396225e5e4fdf503405be8408151c80a|0.6978248568085081|35.209978091326001|00072036881434|FRESH PRODUCE|PRODUCE|-80.844274|80.844275067692323|208|1
35.204336|ed0ebf485f36ecef1064d40a01b23c4216764cce|13.98|2015-02-19 19:53:00|80.828402574597021|4|4900002890|61|35.214435120733839|0|8|54|-80.80146|8|35.17739|DIET|3.49|23|COKE ZERO 12 OZ FRIDGEPACK CN|38847650396225e5e4fdf503405be8408151c80a|0.6978248568085081|35.209978091326001|00049000042559|CARBONATED BEVERAGES|BEVERAGE|-80.844274|80.844275067692323|208|2
35.204336|5255785b2b81d2614cfbfc2bec08416ddfae2843|9.99|2014-09-24 19:59:00|80.828402574597021|4|4113700387|61|35.214435120733839|0|8|386|-80.80146|65|35.17739|NFS-FIREPLACE LOGS|0.0|1|DURAFLAME STAX FIRELOGS|38847650396225e5e4fdf503405be8408151c80a|0.6978248568085081|35.209978091326001|00041137003878|CHARCOAL/LOGS/ACCESSORIES|G1 GROCERY|-80.844274|80.844275067692323|208|1
35.204336|cfb73cf19d70976089cfacdc5a96121326a8fc5f|6.79|2014-09-26 18:35:00|80.828402574597021|4|31031031805|61|35.214435120733839|0|8|4026|-80.80146|1080|35.17739|ORAL HYGI ORAL MEDICATN|0.0|17|ORAJEL MOUTH-AID (GEL)|38847650396225e5e4fdf503405be8408151c80a|0.6978248568085081|35.209978091326001|00310310318055|ORAL HYGIENE|HBC|-80.844274|80.844275067692323|208|1
35.204336|6061e822eba92a6cda5e7489b741078db6b49f1c|4.13|2014-10-27 11:49:00|80.828402574597021|4|20667200000|61|35.214435120733839|0|8|2019|-80.80146|505|35.17739|PRESSED COOKED CHEESE|0.0|6|JARLSBERG LITE (FC)|38847650396225e5e4fdf503405be8408151c80a|0.6978248568085081|35.209978091326001|00206672000007|SPECIALTY CHEESE|DELI|-80.844274|80.844275067692323|208|1
35.204336|076351e209eb2380cf9fdcdffec39d31ea64e110|3.69|2014-12-30 18:55:00|80.828402574597021|4|5150004815|61|35.214435120733839|0|8|1270|-80.80146|41|35.17739|SWEET BREAKFAST|0.0|5|SMUCKERS RED SUG WHL WHT STBRY|38847650396225e5e4fdf503405be8408151c80a|0.6978248568085081|35.209978091326001|00051500041383|BREAKFAST FOODS FROZEN|FROZEN|-80.844274|80.844275067692323|208|1
35.204336|5c306a7ff50fd65445ce8f470369b11d4c771d58|1.69|2015-01-01 13:07:00|80.828402574597021|4|4900000044|61|35.214435120733839|0|8|54|-80.80146|8|35.17739|DIET|0.0|23|CB COKE ZERO 20 OZ|38847650396225e5e4fdf503405be8408151c80a|0.6978248568085081|35.209978091326001|00049000040869|CARBONATED BEVERAGES|BEVERAGE|-80.844274|80.844275067692323|208|1
35.204336|623c616bf4f791d1345015d69552a437eb428356|5.33|2014-12-12 16:59:00|80.828402574597021|4||61|35.214435120733839|0|8|561|-80.80146|64|35.17739|FR PROD ORGANIC PRODUCE|1.5|4|ORG RED DEL APPLES|38847650396225e5e4fdf503405be8408151c80a|0.6978248568085081|35.209978091326001|00294016000004|FRESH PRODUCE|PRODUCE|-80.844274|80.844275067692323|208|1
35.204336|31342028eb067ade16b71f5110cd45f57ab40388|1.69|2015-01-30 19:07:00|80.828402574597021|4|1200000129|61|35.214435120733839|0|8|55|-80.80146|8|35.17739|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|38847650396225e5e4fdf503405be8408151c80a|0.6978248568085081|35.209978091326001|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.844274|80.844275067692323|208|1
35.204336|d8398c193c8d8ff52461eae0c15b5285281d9be7|8.99|2014-11-19 16:14:00|80.828402574597021|4|2188830231|61|35.214435120733839|0|8|4615|-80.80146|1215|35.17739|VITAMIN-MULTIPLE-ADULT|0.0|17|KIDS ONE CHEWABLE MULTIVITAMIN|38847650396225e5e4fdf503405be8408151c80a|0.6978248568085081|35.209978091326001|00021888302314|VITAMINS & SUPPLEMENTS|HBC|-80.844274|80.844275067692323|208|1
35.204336|7f58958ca4dc5b68dc63e06f80d5b7c90e59ea84|1.69|2014-10-15 12:00:00|80.828402574597021|4|4900000044|61|35.214435120733839|0|8|54|-80.80146|8|35.17739|DIET|0.0|23|CB DIET SPRITE ZERO20OZ|38847650396225e5e4fdf503405be8408151c80a|0.6978248568085081|35.209978091326001|00049000037197|CARBONATED BEVERAGES|BEVERAGE|-80.844274|80.844275067692323|208|1
35.318911|6acddcb4b58c424e918733d23db7109bff35c486|2.85|2014-10-12 13:43:00|1.4094857484078087|2|4112907700|167|0.616431285168843|0|26|1219|-80.780702|275|35.318911|PASTA SC CORE|0.85|1|CLASSICO SC ROASTED GARLIC|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00041129077825|PASTA SAUCES|G1 GROCERY|-80.780702|1.4098892219723687|167|1
35.318911|fe5ed4f30e216d3187ce5c4ddecc8b47c863e31d|12.99|2014-10-03 22:06:00|1.4094857484078087|2|4110080673|167|0.616431285168843|0|26|4379|-80.780702|1210|35.318911|ACID BLOCKER-SWALLOW|0.0|17|L ZEGERID|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00041100806734|STOMACH REMEDIES|HBC|-80.780702|1.4098892219723687|167|1
35.318911|e452cd12127b8cee8358980fafc33560d530557a|8.99|2014-12-04 12:49:00|1.4094857484078087|2|4132211080|167|0.616431285168843|0|26|293|-80.780702|48|35.318911|FROZEN SEAFOOD|3.0|5|SEAPAK SHRIMP SCAMPI|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00041322110800|FROZEN MEALS|FROZEN|-80.780702|1.4098892219723687|167|1
35.318911|3067e6343daed2d0db3e622d803b3eb421abbfe0|17.98|2015-02-04 14:13:00|1.4094857484078087|2|4132211080|167|0.616431285168843|0|26|293|-80.780702|48|35.318911|FROZEN SEAFOOD|7.98|5|SEAPAK SHRIMP SCAMPI|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00041322110800|FROZEN MEALS|FROZEN|-80.780702|1.4098892219723687|167|2
35.318911|f35b42410e827f8074ce187bfb464db08753b501|5.79|2014-11-16 16:04:00|1.4094857484078087|2|20165700000|167|0.616431285168843|0|26|297|-80.780702|49|35.318911|GROUND BEEF|1.29|2|HT GROUND BEEF CHUCK 80% LEAN|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00201657000003|BEEF|MEAT|-80.780702|1.4098892219723687|167|1
35.318911|06e94ed024974bd5d5daf32fd935a2b3df5f18ae|5.43|2014-10-02 17:30:00|1.4094857484078087|2|20165700000|167|0.616431285168843|0|26|297|-80.780702|49|35.318911|GROUND BEEF|0.6|2|HT GROUND BEEF CHUCK 80% LEAN|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00201657000003|BEEF|MEAT|-80.780702|1.4098892219723687|167|1
35.318911|ed972d79f3c4316aaca67e162546411a8e4417cb|2.45|2015-02-09 13:21:00|1.4094857484078087|2|5100013279|167|0.616431285168843|0|26|214|-80.780702|33|35.318911|BROTH|0.0|1|SWANSON BROTH LOW SOD CHICKEN|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00051000132796|SOUP|G1 GROCERY|-80.780702|1.4098892219723687|167|1
35.318911|9fed38576f9288cfe54762fa9f40404f8a5e0c8f|3.85|2014-12-28 11:11:00|1.4094857484078087|2|4812127620|167|0.616431285168843|0|26|1037|-80.780702|164|35.318911|ENGLISH MUFFINS|1.93|7|THOMAS HIGH FIBER PLAIN EM PP|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00048121181086|BREAKFAST|COMMERCIAL BAKERY|-80.780702|1.4098892219723687|167|1
35.318911|d52699e9a79ac5881e96303eb87598be78d18f4f|2.69|2014-09-21 19:26:00|1.4094857484078087|2|7203663996|167|0.616431285168843|0|26|342|-80.780702|57|35.318911|FRESH MILK|0.0|3|HARRIS TEETER WHOLE MILK|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00072036639967|MILK|DAIRY|-80.780702|1.4098892219723687|167|1
35.318911|3879578ff40e238eb99246deb27d81f5778ec1f4|2.29|2015-02-06 22:10:00|1.4094857484078087|2|7203663996|167|0.616431285168843|0|26|342|-80.780702|57|35.318911|FRESH MILK|0.0|3|HARRIS TEETER WHOLE MILK|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00072036639967|MILK|DAIRY|-80.780702|1.4098892219723687|167|1
35.318911|483fe76506f0f54c58afe0288d30c27b86ce8e22|2.49|2014-12-16 17:13:00|1.4094857484078087|2|7203663996|167|0.616431285168843|0|26|342|-80.780702|57|35.318911|FRESH MILK|0.0|3|HARRIS TEETER WHOLE MILK|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00072036639967|MILK|DAIRY|-80.780702|1.4098892219723687|167|1
35.318911|33aa31dcf202787a2a076d453d3e2839581ec4f4|2.29|2015-01-15 17:15:00|1.4094857484078087|2|7203663996|167|0.616431285168843|0|26|342|-80.780702|57|35.318911|FRESH MILK|0.0|3|HARRIS TEETER WHOLE MILK|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00072036639967|MILK|DAIRY|-80.780702|1.4098892219723687|167|1
35.318911|eebf96457e12198eadb36d9b7244dc39c7a51d38|1.67|2014-12-15 17:03:00|80.77969194620016|2|7203670564|167|35.330740396555015|0|20|416|-80.737839|71|35.297134|NFS-BLEACH|0.0|1|YH BLEACH|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|35.345012799095393|00072036705648|LAUNDRY SUPPLIES|G1 GROCERY|-80.780702|80.780702457814314|258|1
35.318911|57d317772c73d971080d25fe894138eb51d19248|2.69|2014-09-13 17:36:00|1.4094857484078087|2|7203663996|167|0.616431285168843|0|26|342|-80.780702|57|35.318911|FRESH MILK|0.0|3|HARRIS TEETER WHOLE MILK|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00072036639967|MILK|DAIRY|-80.780702|1.4098892219723687|167|1
35.318911|1ea494e18b02f46eb1a168014ff5642126658575|2.69|2014-09-17 18:31:00|80.77969194620016|2|7203663996|167|35.330740396555015|0|20|342|-80.737839|57|35.297134|FRESH MILK|0.0|3|HARRIS TEETER WHOLE MILK|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|35.345012799095393|00072036639967|MILK|DAIRY|-80.780702|80.780702457814314|258|1
35.318911|17e9e8ac0b4e9039775583dc59a78e20a32b6c13|2.59|2014-10-28 16:28:00|1.4094857484078087|2|7203663996|167|0.616431285168843|0|26|342|-80.780702|57|35.318911|FRESH MILK|0.0|3|HARRIS TEETER WHOLE MILK|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00072036639967|MILK|DAIRY|-80.780702|1.4098892219723687|167|1
35.318911|1a6512f79a93d1846314cadab4d6639e69b8a575|2.59|2014-11-22 10:11:00|1.4094857484078087|2|7203663996|167|0.616431285168843|0|26|342|-80.780702|57|35.318911|FRESH MILK|0.82|3|HARRIS TEETER WHOLE MILK|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00072036639967|MILK|DAIRY|-80.780702|1.4098892219723687|167|1
35.318911|2ca86593b1deab7818e9a0e068332cc4d942bea0|2.59|2014-11-07 15:59:00|1.4094857484078087|2|7203663996|167|0.616431285168843|0|26|342|-80.780702|57|35.318911|FRESH MILK|0.0|3|HARRIS TEETER WHOLE MILK|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00072036639967|MILK|DAIRY|-80.780702|1.4098892219723687|167|1
35.318911|7a03bc9e76bbe35d19f388ce2aa216c85e76d985|2.29|2015-01-08 13:12:00|1.4094857484078087|2|7203663996|167|0.616431285168843|0|26|342|-80.780702|57|35.318911|FRESH MILK|0.0|3|HARRIS TEETER WHOLE MILK|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00072036639967|MILK|DAIRY|-80.780702|1.4098892219723687|167|1
35.318911|f5adf279b09d2944f9ba8af8a5ce8f67039ff2dd|4.19|2015-02-19 16:11:00|1.4094857484078087|2|7203663089|167|0.616431285168843|0|26|345|-80.780702|57|35.318911|ORGANIC MILK|0.0|3|HTO ORGANIC CRTN WHOLE MILK|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00072036763860|MILK|DAIRY|-80.780702|1.4098892219723687|167|1
35.318911|5612b84db9575ffb5676349537c5c73bd33e0c42|4.79|2014-10-19 17:55:00|1.4094857484078087|2|76172098749|167|0.616431285168843|0|26|195|-80.780702|30|35.318911|SALAD & COOKING OIL|0.0|1|MAZOLA CORN OIL|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00761720987490|SHORTENING/OIL|G1 GROCERY|-80.780702|1.4098892219723687|167|1
35.318911|24bf066bfb00c5c68f57752547599eb854ac510e|1.89|2014-12-18 13:52:00|1.4094857484078087|2|5150020430|167|0.616431285168843|0|26|101|-80.780702|15|35.318911|FLOUR-ALL PURPOSE|0.0|1|PILLSBURY ALL PURPOSE FLOUR|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00051500204306|FLOUR|G1 GROCERY|-80.780702|1.4098892219723687|167|1
35.318911|c4af3e4195fd92306775fc2a7c751cb09dad76d5|8.35|2014-12-21 14:49:00|1.4094857484078087|2|76211188813|167|0.616431285168843|0|26|37|-80.780702|10|35.318911|PODS/CUPS/SINGLES|1.36|1|STARBUCKS HOUSE BLEND KCUP|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00762111888136|COFFEE|G1 GROCERY|-80.780702|1.4098892219723687|167|1
35.318911|a96dd3c2ad39f6203b61877ad13ad399b59d0056|4.23|2015-02-01 14:45:00|1.4094857484078087|2||167|0.616431285168843|0|26|529|-80.780702|64|35.318911|FRESH ASPARAGUS|2.12|4|GREEN  ASPARAGUS|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00204080000008|FRESH PRODUCE|PRODUCE|-80.780702|1.4098892219723687|167|1
35.318911|f38bb55eca1ad6c97ecaf7e8fd0ba0bfdd71336f|7.58|2014-12-19 15:15:00|1.4094857484078087|2|2100062503|167|0.616431285168843|0|26|318|-80.780702|52|35.318911|SHREDDED/GRATED CHEESE|1.29|3|KRAFT FINELY SHREDDED SHARP C|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00021000638741|CHEESE|DAIRY|-80.780702|1.4098892219723687|167|2
35.318911|b8c9568fe79d37910e8f326bd79c6e2f2ed12991|6.99|2015-01-21 21:09:00|80.77969194620016|2|7309102222|167|35.330740396555015|0|20|6901|-80.737839|1582|35.297134|DOG MEDICINES|0.0|18|VETSCRIPT ANITITCH SPRY DG/CT|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|35.345012799095393|00073091022220|PET NEEDS|GM|-80.780702|80.780702457814314|258|1
35.318911|b7bf802d25474528c61a7d58e5f7762aaf3d51c6|0.47|2015-02-05 16:00:00|1.4094857484078087|2|7248600220|167|0.616431285168843|0|26|11|-80.780702|2|35.318911|MUFFIN MIXES|0.0|1|JIFFY CORN MUFFIN MIX|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00072486002205|BAKING MIXES|G1 GROCERY|-80.780702|1.4098892219723687|167|1
35.318911|13849d05227b8b24c458786d99d0e0da3bd8ab1c|0.47|2014-11-01 10:43:00|80.77969194620016|2|7248600220|167|35.330740396560884|0|20|11|-80.814133|2|35.333742|MUFFIN MIXES|0.0|1|JIFFY CORN MUFFIN MIX|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|35.345012799095393|00072486002205|BAKING MIXES|G1 GROCERY|-80.780702|80.78070203228107|472|1
35.318911|aea52fd39eab89955f1134308b8d8f1ff7a8287f|15.98|2015-03-05 13:20:00|1.4094857484078087|2|20176400000|167|0.616431285168843|0|26|636|-80.780702|49|35.318911|MARINATED BEEF|0.0|2|HT RANCHER GARLIC PETITE TNDR|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00201764000002|BEEF|MEAT|-80.780702|1.4098892219723687|167|1
35.318911|cb6b18e96ec0b0d57ba16efc2440a7d6594a2f3a|1.34|2014-10-31 14:34:00|1.4094857484078087|2|7203653081|167|0.616431285168843|0|26|1275|-80.780702|50|35.318911|BOX VEG|0.34|5|HT CHOPPED SPINACH|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00072036530813|VEGETABLES-FROZEN|FROZEN|-80.780702|1.4098892219723687|167|1
35.318911|f9bc0afabf635bbb5d42a54847c88e2d569abd5f|1.34|2015-01-27 15:39:00|80.77969194620016|2|7203653081|167|35.330740396555015|0|20|1275|-80.737839|50|35.297134|BOX VEG|0.0|5|HT CHOPPED SPINACH|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|35.345012799095393|00072036530813|VEGETABLES-FROZEN|FROZEN|-80.780702|80.780702457814314|258|1
35.318911|2c9d191d2ec3f50d7d2cfbd6ff2d964d1739d5a6|18.99|2015-02-21 16:11:00|80.77969194620016|2|6574311526|167|35.330740396555015|0|20|3476|-80.737839|1040|35.297134|BRAND-PAUL MITCHELL|0.0|17|P MITCHELL T/TREE LAV MINT CND|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|35.345012799095393|00065743115268|PROFESSIONAL HAIR & SCALP CARE|HBC|-80.780702|80.780702457814314|258|1
35.318911|15d1a396cb0db1d3426712c3fb5dc794171abd17|4.19|2014-10-13 14:31:00|1.4094857484078087|2|4812127620|167|0.616431285168843|0|26|1037|-80.780702|164|35.318911|ENGLISH MUFFINS|2.09|7|THOMAS SEASONAL EM PP|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00048121221003|BREAKFAST|COMMERCIAL BAKERY|-80.780702|1.4098892219723687|167|1
35.318911|b772da0350d199d54da71f19e0bc99497f2723b7|2.89|2014-12-06 13:17:00|1.4094857484078087|2|7203663102|167|0.616431285168843|0|26|339|-80.780702|57|35.318911|EGGNOGS/DRINKS|0.89|3|I/O HARRIS TEETER EGG NOG|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00072036631022|MILK|DAIRY|-80.780702|1.4098892219723687|167|1
35.318911|b6ae8042926ea34abce2166ff56658902d4dbadc|2.19|2015-01-13 18:34:00|80.77969194620016|2|76857300210|167|35.330740396555015|0|20|544|-80.737839|64|35.297134|FRESH PRODUCE FRSH HERBS|0.0|4|PKG FRESH DILL|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|35.345012799095393|00768573002103|FRESH PRODUCE|PRODUCE|-80.780702|80.780702457814314|258|1
35.318911|2fefc26ea3fc8d2586cafc5bd44fef0840c73b92|4.49|2015-01-11 08:21:00|80.77969194620016|2|7203698586|167|35.33074039301804|0|20|66|-80.8955|10|35.4437|GROUND CAN|0.0|1|HT CLASSIC DECAF CAN COFFEE|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|35.345012799095393|00072036985866|COFFEE|G1 GROCERY|-80.780702|80.780713221322245|272|1
35.318911|39a6214dfc976b13ef1b5310ae8d36e7c3bfab59|3.29|2015-01-29 14:47:00|80.77969194620016|2|7225091171|167|35.330740396560884|0|20|1033|-80.814133|163|35.333742|HAMBURGER|0.0|7|NATOWN WHITEWHEAT HAMS|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|35.345012799095393|00072250911719|BUNS/ROLLS|COMMERCIAL BAKERY|-80.780702|80.78070203228107|472|1
35.318911|574bde94b64af7c6a98281aeca7035a186ad1fc9|13.98|2015-01-04 14:15:00|1.4094857484078087|2|3700013885|167|0.616431285168843|0|26|389|-80.780702|66|35.318911|NFS-LAUNDRY DETERGENTS|1.0|1|TIDE ULTRA STAIN RELEASE 46OZ|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00037000875864|DETERGENTS|G1 GROCERY|-80.780702|1.4098892219723687|167|2
35.318911|b6cb51cd1466b59a969f1d81ae7fb6b4fd04d792|5.99|2014-11-14 17:51:00|80.77969194620016|2|7203698286|167|35.330740396560884|0|20|3917|-80.814133|1075|35.333742|DISPOSABLE RAZOE-MEN|0.0|17|HT 6 BLADE DSPBL RAZOR MEN|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|35.345012799095393|00072036982865|SHAVING NEEDS/MEN HAIR|HBC|-80.780702|80.78070203228107|472|1
35.318911|6896695e4155f7ceca3be218c3401d2b91795614|7.99|2015-01-17 20:50:00|80.77969194620016|2|1820017993|167|35.33074039301804|0|20|458|-80.8955|82|35.4437|CRAFT BEER|0.0|16|SHOCK TOP SEASONAL 6PK|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|35.345012799095393|00018200179938|DOMESTIC BEER|BEER|-80.780702|80.780713221322245|272|1
35.318911|e507b4da7a074ccaa35240434ae3fa44a0a78e90|2.78|2015-01-01 09:27:00|80.77969194620016|2|2310034974|167|35.330740395982367|0|20|158|-80.764523|24|35.341927|NFS-DOG FOOD-WET|0.0|1|PEDIGREE PLUS HLTHY DIGESTION|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|35.345012799095393|00023100349732|PET FOOD/SUPPLIES|G1 GROCERY|-80.780702|80.78070653453473|220|2
35.318911|630cd5d632296c369d3bb43c3e31bd4d654fb30c|13.29|2014-12-22 18:15:00|80.77969194620016|2|3700013882|167|35.330740396560884|0|20|389|-80.814133|66|35.333742|NFS-LAUNDRY DETERGENTS|0.0|1|TIDE ORIGINAL 64LD|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|35.345012799095393|00037000138822|DETERGENTS|G1 GROCERY|-80.780702|80.78070203228107|472|1
35.318911|0329990ab1d090c4a1bff22fe4686f9e814a8847|3.34|2014-09-26 17:16:00|1.4094857484078087|2|3663201899|167|0.616431285168843|0|26|343|-80.780702|59|35.318911|PUDDINGS|0.67|3|CREAMERY CHERRY CHEESECAKE|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00036632018939|SNACKS/SPREADS/DIPS-DAIRY|DAIRY|-80.780702|1.4098892219723687|167|2
35.318911|5b30c3eb625b188cee17ec75ac5983450520c9b1|15.96|2015-02-01 08:07:00|80.77969194620016|2|3000005620|167|35.33074039301804|0|20|228|-80.8955|36|35.4437|TABLE SYRUP|5.96|1|AUNT JEMIMA ORIGINAL SYRUP|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|35.345012799095393|00030000059708|TABLE SYRUPS|G1 GROCERY|-80.780702|80.780713221322245|272|4
35.318911|04676d151204509c7a7ce3088fae3784bbdaa0e7|13.25|2015-01-12 19:12:00|1.4094857484078087|2|3700088211|167|0.616431285168843|0|26|426|-80.780702|72|35.318911|NFS-PAPER TOWELS|0.0|1|BOUNTY TOWEL 8 GIANT WHITE|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00037000882138|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.780702|1.4098892219723687|167|1
35.318911|9d80bc33e8143f0985b71193e3e9737e08b21c10|15.98|2015-02-21 08:44:00|80.77969194620016|2|2550000371|167|35.33074039301804|0|20|66|-80.8955|10|35.4437|GROUND CAN|0.0|1|FOLGERS CLASSIC DECAF CAN|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|35.345012799095393|00025500003719|COFFEE|G1 GROCERY|-80.780702|80.780713221322245|272|2
35.318911|e03cc3e53da4594d873f5423690c7eb605659b20|39.98|2014-09-21 08:20:00|80.77969194620016|2|3057614032|167|35.33074039301804|0|20|228|-80.8955|36|35.4437|TABLE SYRUP|0.0|1|ANDERSON'S PUR MAPL SYRUP 32OZ|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|35.345012799095393|00030576140329|TABLE SYRUPS|G1 GROCERY|-80.780702|80.780713221322245|272|2
35.318911|ca505340aeb61268ef89e98b5d07ed2cd2aa58a6|9.17|2014-09-21 08:23:00|80.77969194620016|2||167|35.33074039301804|0|20|502|-80.8955|64|35.4437|FRESH BANANAS|0.0|4|BANANAS, YELLOW|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|35.345012799095393|00204011000008|FRESH PRODUCE|PRODUCE|-80.780702|80.780713221322245|272|4
35.318911|cf798f14d830b11549bc347b08bcdefebf964898|0.85|2015-01-26 16:03:00|1.4094857484078087|2||167|0.616431285168843|0|26|502|-80.780702|64|35.318911|FRESH BANANAS|0.0|4|BANANAS, YELLOW|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00204011000008|FRESH PRODUCE|PRODUCE|-80.780702|1.4098892219723687|167|1
35.318911|3055fdfa3d3f496da50f33be6f0a3ef26cdf1234|6.99|2014-11-29 22:10:00|1.4094857484078087|2|7203698720|167|0.616431285168843|0|26|6899|-80.780702|1582|35.318911|DOG HOUSEBREAKING PADS|0.0|18|YP DELUXE PUPPY PADS-14CT|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00072036987204|PET NEEDS|GM|-80.780702|1.4098892219723687|167|1
35.318911|2608d62d9c33856df52b4b5025170c535ad54e84|6.99|2014-12-20 22:59:00|1.4094857484078087|2|7203698720|167|0.616431285168843|0|26|6899|-80.780702|1582|35.318911|DOG HOUSEBREAKING PADS|0.0|18|YP DELUXE PUPPY PADS-14CT|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00072036987204|PET NEEDS|GM|-80.780702|1.4098892219723687|167|1
35.318911|a30ac8c5d2a9041bdea005eeaa7de1be628f435d|5.29|2014-10-21 16:37:00|1.4094857484078087|2|7033060845|167|0.616431285168843|0|26|8727|-80.780702|1810|35.318911|LIGHTER|0.0|18|(JHK)(PPL)(FE) BIC SUR S LGHTR|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00070330608450|LIGHTERS|GM|-80.780702|1.4098892219723687|167|1
35.318911|834e714ef0c94b69bf21f672b3eb333b87674b2c|11.59|2015-01-04 01:15:00|1.4094857484078087|2|30573016940|167|0.616431285168843|0|26|4317|-80.780702|1205|35.318911|IBUPROFEN|0.0|17|ADVIL LIQUI-GELS  -16940|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00305730169400|PAIN RELIEF|HBC|-80.780702|1.4098892219723687|167|1
35.318911|247efaf3ab574fa7739bd8c53cbb4a780fcc722f|5.3|2015-01-26 16:11:00|1.4094857484078087|2|2100061223|167|0.616431285168843|0|26|316|-80.780702|52|35.318911|CREAM CHEESE|1.3|3|PHILLY CREAM CHEESE - BRICK|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00021000612239|CHEESE|DAIRY|-80.780702|1.4098892219723687|167|2
35.318911|816c41886beb4d788978b252b771933b5e801ad4|0.97|2015-01-01 14:50:00|80.77969194620016|2|7203698757|167|35.330740396560884|0|20|31|-80.814133|4|35.333742|NON CARBONATED WATER|0.0|1|HT DISTILLED WATER|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|35.345012799095393|00072036360601|BOTTLED WATER|G1 GROCERY|-80.780702|80.78070203228107|472|1
35.318911|e75c76ea1f23bb8af139f8169278f839ac0df42d|1.79|2015-01-24 18:03:00|1.4094857484078087|2|7203663220|167|0.616431285168843|0|26|330|-80.780702|55|35.318911|EGGS|0.0|3|HT GRADE A    LARGE EGGS|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|0.61471665291522548|00072036632203|EGGS FRESH|DAIRY|-80.780702|1.4098892219723687|167|1
35.318911|6402db00af52dc6f5ceb5124b49c096c3ec3ab31|10.88|2014-10-27 18:15:00|80.77969194620016|2|20596800000|167|35.330740395982367|0|20|1821|-80.764523|410|35.341927|BH TURKEY|0.0|6|BOARS HEAD CAJUN TURKEY|39ee9e1c3d548a25a6b249ece4145d908f926aa1|0.8173827353883971|35.345012799095393|00205968000004|BH MEAT|DELI|-80.780702|80.78070653453473|220|1
35.124987|8adae4bf5b62c22d471cc541528077e95c529b33|8.91|2014-12-10 19:23:00|1.4091206135396188|1|7203658035|157|0.6130466728702054|0|47|358|-80.709466|100|35.124987|REGULAR BACON|0.0|19|HT LOW SALT SLICED BACON|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00072036590237|BACON|CASE READY MEATS|-80.709466|1.4086459192264178|157|3
35.124987|66524f89a4fa3865d43051ebe5503877f6244092|3.35|2014-09-24 14:56:00|80.7095026033777|1|7203656080|157|35.139506220647377|0|51|318|-80.70901|52|35.17335|SHREDDED/GRATED CHEESE|0.0|3|HT NACHO TACO MEXICAN BLEND|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00072036560834|CHEESE|DAIRY|-80.709466|80.709474979800646|174|1
35.124987|29ba1180d7c25684a3285fb09164921f0651c3da|9.98|2015-01-08 14:44:00|1.4091206135396188|1|7203688080|157|0.6130466728702054|0|47|523|-80.709466|64|35.124987|FRESH POTATOES|2.49|4|HT YUKON GOLD 5 LB BAG|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00072036880802|FRESH PRODUCE|PRODUCE|-80.709466|1.4086459192264178|157|2
35.124987|827f650ec8d903cc37e6aa92cf780025f09c791d|14.97|2015-03-08 11:04:00|80.7095026033777|1|7418226981|157|35.139506220647377|0|51|722|-80.70901|73|35.17335|NFS-HAND SOAPS|4.47|1|SS HAND SOAP REFILL AQUARIUM|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00074182269852|PERSONAL SOAP/BATH ADDITIVES|G1 GROCERY|-80.709466|80.709474979800646|174|3
35.124987|afe52e75220302aedc3f33d61ccc73bec2241930|15.920000000000002|2015-01-22 14:39:00|1.4091206135396188|1|7418226981|157|0.6130466728702054|0|47|722|-80.709466|73|35.124987|NFS-HAND SOAPS|0.0|1|SS HAND SOAP REFILL AQUARIUM|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00074182269852|PERSONAL SOAP/BATH ADDITIVES|G1 GROCERY|-80.709466|1.4086459192264178|157|4
35.124987|d844b6c9600bc3de78e5d4708edec6a5351469a5|1.29|2015-02-27 19:30:00|1.4091206135396188|1|8379152001|157|0.6130466728702054|0|47|1981|-80.709466|480|35.124987|CHIPS|0.0|6|DIRTY POTATO CHIP BBQ|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00083791520049|DRY GOODS|DELI|-80.709466|1.4086459192264178|157|1
35.124987|fb6d1f7bda8f0a77fbf47f371fd8ab0dc8516fdf|2.68|2015-01-22 14:13:00|1.4091206135396188|1|8000000673|157|0.6130466728702054|0|47|190|-80.709466|29|35.124987|TUNA-CANNED|0.0|1|STARKIST TUNA CHUNK LIGHT|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00080000006738|SEAFOOD-CANNED|G1 GROCERY|-80.709466|1.4086459192264178|157|4
35.124987|fadb87048b2108e6e2346944d59b44f83b81e434|18.47|2014-11-03 17:59:00|80.7095026033777|1||157|35.139506222092137|0|51|500|-80.654118|64|35.123768|FRESH APPLES|6.94|4|HONEY CRISP APPLE|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00233283000003|FRESH PRODUCE|PRODUCE|-80.709466|80.709470232147311|473|1
35.124987|d9e4f26e6a169b02ee421e0e0a9fe86db58f4ffc|4.19|2014-10-20 18:50:00|1.4091206135396188|1|60308424372|157|0.6130466728702054|0|47|3606|-80.709466|1050|35.124987|SETTING LOTIONS|1.2|17|S/T FRUCTIS SMOOTHING MILK|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00603084260249|HAIR STYLING|HBC|-80.709466|1.4086459192264178|157|1
35.124987|a4d87061a53ff65f7b5ca2b0e464786c704c865e|15.98|2014-11-01 11:16:00|80.7095026033777|1|30521026958|157|35.139506222495768|0|51|3200|-80.739|1015|35.141204|HAND & BODY EXPERIENTIAL|4.0|17|VICL SPRAY COCOA LOTION|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00305210269637|HAND & BODY LOTION/SUN CARE|HBC|-80.709466|80.709466621902877|171|2
35.124987|6b3db02bbaf331fd00e050d247db55b631b90f99|16.38|2014-09-16 11:27:00|80.7095026033777|1|20896500000|157|35.139506222495768|0|51|977|-80.739|201|35.141204|FRESH HT CHICKEN|0.0|2|HT FRESH CHICKEN DRUMMETTES|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00208965000008|POULTRY|MEAT|-80.709466|80.709466621902877|171|6
35.124987|460d0c61cdd01e78bb2f1b424f3e22e76cfcee72|1.07|2015-02-21 11:47:00|1.4091206135396188|1||157|0.6130466728702054|0|47|522|-80.709466|64|35.124987|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00204664000004|FRESH PRODUCE|PRODUCE|-80.709466|1.4086459192264178|157|1
35.124987|c3b11c8c6fb89be2f08d296b47cbd2d481c486e4|8.59|2015-01-10 12:46:00|1.4091206135396188|1|7431207580|157|0.6130466728702054|0|47|4582|-80.709466|1215|35.124987|SPLMNT-WOMENS|0.0|17|NB HAIR SKIN AND NAILS|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00074312075803|VITAMINS & SUPPLEMENTS|HBC|-80.709466|1.4086459192264178|157|1
35.124987|7b629ab307d91759f9bd41dced4bd6df150dd2f3|5.78|2014-10-18 15:33:00|1.4091206135396188|1|8768400095|157|0.6130466728702054|0|47|121|-80.709466|20|35.124987|ASEPTIC JUICES|0.78|1|CAPRI SUN SPLASH COOLER 10PK|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00087684000977|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.709466|1.4086459192264178|157|2
35.124987|fc3909d4ebecd443f66e91e9eeee1115ddc57242|3.52|2015-01-10 12:14:00|1.4091206135396188|1|20196000000|157|0.6130466728702054|0|47|299|-80.709466|49|35.124987|ANGUS BEEF|0.44|2|ANGUS BF FLAT IRON STK CUSTOM|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00201960000004|BEEF|MEAT|-80.709466|1.4086459192264178|157|1
35.124987|9673137db0260cd9a8065dfb2c9b165c247ad08e|8.0|2014-12-21 16:38:00|80.7095026033777|1|4300000953|157|35.139506220647377|0|51|272|-80.70901|307|35.17335|TOPPINGS FROZEN|4.04|5|COOL WHIP WHIPPED TOPPING|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00043000009536|DESSERTS FROZEN|FROZEN|-80.709466|80.709474979800646|174|4
35.124987|11ef3c14ecb02cb227cdddc7fef2ae2b7479ca4c|9.38|2014-10-08 12:22:00|1.4091206135396188|1|4460030770|157|0.6130466728702054|0|47|416|-80.709466|71|35.124987|NFS-BLEACH|2.35|1|CLOROX BLEACH FRSH MEADOW CONC|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00044600307763|LAUNDRY SUPPLIES|G1 GROCERY|-80.709466|1.4086459192264178|157|2
35.124987|91f06941de59a9cd982c3d58306ae7cf1b10be90|5.98|2014-11-01 11:14:00|80.7095026033777|1|20894700000|157|35.139506222495768|0|51|977|-80.739|201|35.141204|FRESH HT CHICKEN|0.0|2|HT WHOLE CHICKEN|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00208947000002|POULTRY|MEAT|-80.709466|80.709466621902877|171|1
35.124987|0c0ada1ce11809d65b9823f821464d86763ef0a8|30.110000000000003|2015-01-22 17:36:00|1.4091206135396188|1|20894700000|157|0.6130466728702054|0|47|977|-80.709466|201|35.124987|FRESH HT CHICKEN|0.0|2|HT WHOLE CHICKEN|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00208947000002|POULTRY|MEAT|-80.709466|1.4086459192264178|157|12
35.124987|b540b806f272da8c58a4c6b58f947a363886b40c|9.49|2014-12-04 17:33:00|1.4091206135396188|1|2301290173|157|0.6130466728702054|0|47|1477|-80.709466|485|35.124987|SUSHI HYBRID|0.0|6|CRUNCHY DRAGON ROLL SP BR|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00023012901738|SUSHI|DELI|-80.709466|1.4086459192264178|157|1
35.124987|3eb08739cf8ecc801f3be8e36729d949cef49a84|3.5|2014-09-27 11:26:00|80.7095026033777|1|2920000212|157|35.139506222092137|0|51|149|-80.654118|23|35.123768|WHSE PASTA CORE|0.88|1|MUELLER ELBOW MACARONI|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00029200002133|PASTA|G1 GROCERY|-80.709466|80.709470232147311|473|2
35.124987|293989471f27f1c249e2a3715d23aedcc3359435|3.99|2014-10-04 15:44:00|1.4091206135396188|1|2500005542|157|0.6130466728702054|0|47|335|-80.709466|56|35.124987|ORANGE JUICE-REGRIGERATED|0.99|3|SIMPLY ORANGE ORIGINAL|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00025000055423|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.709466|1.4086459192264178|157|1
35.124987|8dcd152c191c182552a814eed713fc9dafac15dd|3.69|2015-03-01 11:01:00|80.7095026033777|1|2500005542|157|35.139506220647377|0|51|335|-80.70901|56|35.17335|ORANGE JUICE-REGRIGERATED|0.69|3|SIMPLY ORANGE ORIGINAL|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00025000055423|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.709466|80.709474979800646|174|1
35.124987|8b7efecc517e18698de3335e99c99dad098beb7b|11.99|2014-12-04 17:32:00|1.4091206135396188|1|2301286481|157|0.6130466728702054|0|47|1477|-80.709466|485|35.124987|SUSHI HYBRID|0.0|6|"CHEF SAMPLER ""A"""|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00023012864811|SUSHI|DELI|-80.709466|1.4086459192264178|157|1
35.124987|6c0869f48b38906f03837601bf86da62fc9f9d03|6.99|2015-02-07 10:38:00|1.4091206135396188|1|3700088234|157|0.6130466728702054|0|47|426|-80.709466|72|35.124987|NFS-PAPER TOWELS|0.0|1|BOUNTY TOWEL 2 SAS|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00037000882343|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.709466|1.4086459192264178|157|1
35.124987|d1d4ed06e4e5822708b84663e9ef764ea6f34a4f|3.29|2014-10-11 14:54:00|1.4091206135396188|1|3800031120|157|0.6130466728702054|0|47|44|-80.709466|6|35.124987|TOASTER PASTRIES-SHELF STABLE|0.79|1|KELL POPTART 12CT STRAWBERY|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00038000317200|BREAKFAST FOODS|G1 GROCERY|-80.709466|1.4086459192264178|157|1
35.124987|2a055536f04df0df59215b3a2c3172263d8b5d9e|22.14|2014-12-13 08:39:00|1.4091206135396188|1|3770032217|157|0.6130466728702054|0|47|423|-80.709466|72|35.124987|NFS-DISPOSE PLATES/BOWLS|3.84|1|CHINET LUNCH PLATE 8 3/4|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00037700323085|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.709466|1.4086459192264178|157|6
35.124987|a1b159452bc95b2054153bc28efac174ee4bda49|13.98|2014-12-06 09:20:00|1.4091206135396188|1|3700013885|157|0.6130466728702054|0|47|389|-80.709466|66|35.124987|NFS-LAUNDRY DETERGENTS|1.0|1|TIDE APRIL FRESH DOWNY HE 46OZ|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00037000874720|DETERGENTS|G1 GROCERY|-80.709466|1.4086459192264178|157|2
35.124987|6af897ab4fc9aa4ccad771bd0cd64449a29e6d53|7.95|2014-09-20 16:38:00|1.4091206135396188|1|3800031120|157|0.6130466728702054|0|47|44|-80.709466|6|35.124987|TOASTER PASTRIES-SHELF STABLE|0.0|1|KELL POPTART 12CT STRAWBERY|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00038000317200|BREAKFAST FOODS|G1 GROCERY|-80.709466|1.4086459192264178|157|3
35.124987|d487509a21788f844f20c59c25416fae280f8ab4|6.99|2015-01-03 11:38:00|1.4091206135396188|1|3700013885|157|0.6130466728702054|0|47|389|-80.709466|66|35.124987|NFS-LAUNDRY DETERGENTS|1.0|1|TIDE ULTRA STAIN RELEASE 46OZ|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00037000875864|DETERGENTS|G1 GROCERY|-80.709466|1.4086459192264178|157|1
35.124987|fc4826bbba040cf80642ad80a775f5a3fac293a6|9.98|2014-11-08 10:20:00|1.4091206135396188|1|4720015264|157|0.6130466728702054|0|47|312|-80.709466|51|35.124987|BUTTER|2.98|3|CHALLENGE SALTED BUTTER|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00047200152641|BUTTER & MARGARINE|DAIRY|-80.709466|1.4086459192264178|157|2
35.124987|cefee1119cc8eb9316ffaa4cd4934a9077a8ac37|2.99|2015-02-13 14:14:00|1.4091206135396188|1|4470036113|157|0.6130466728702054|0|47|659|-80.709466|103|35.124987|CHILDRENS LUNCH SNACKS|0.49|19|FUNPACK LUNCH TRKY/AMER STACK|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00044700006740|LUNCH SNACKS|CASE READY MEATS|-80.709466|1.4086459192264178|157|1
35.124987|d3a10a59050de3812c08d496cd9f030a596f5256|16.76|2014-11-14 12:23:00|80.7095026033777|1|5210007086|157|35.139506220346284|0|51|217|-80.732725|34|35.082768|EXTRACTS FOOD COLORING|5.04|1|E  MCCORMICK VANILLA EXTRACT|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00052100070865|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.709466|80.709475680354345|147|4
35.124987|eb33c95cda291fda70344402fe5e9be389158b11|2.99|2014-11-20 12:01:00|80.7095026033777|1|5190000001|157|35.139506222495768|0|51|362|-80.739|102|35.141204|PEPPERONIS|1.5|19|LOF CANADIAN BACON PEPPER|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00051900000027|LUNCHMEATS|CASE READY MEATS|-80.709466|80.709466621902877|171|1
35.124987|6f74389251b393fee4f6f93e0e664a62effd7449|8.38|2014-11-04 13:31:00|80.7095026033777|1|5210007086|157|35.139506220647377|0|51|217|-80.70901|34|35.17335|EXTRACTS FOOD COLORING|2.09|1|E  MCCORMICK VANILLA EXTRACT|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00052100070865|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.709466|80.709474979800646|174|2
35.124987|5869d47c154d6b8aab72bf3f4a8b19c0f75d0f2b|13.58|2014-12-20 09:58:00|1.4091206135396188|1|4900002890|157|0.6130466728702054|0|47|55|-80.709466|8|35.124987|REGULAR|6.79|23|FUZE ICE TEA LEMON 12 PK CAN|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00080793808694|CARBONATED BEVERAGES|BEVERAGE|-80.709466|1.4086459192264178|157|2
35.124987|493b935ecfe14389b8851ae666b0d7c0a4e87937|2.0|2015-02-02 11:06:00|80.7095026033777|1||157|35.139506222092137|0|51|565|-80.654118|64|35.123768|REDUCED PRODUCE|0.0|4|PRODUCE REWRAP BY CT|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00204845000007|FRESH PRODUCE|PRODUCE|-80.709466|80.709470232147311|473|2
35.124987|8d604e328ac479652de72282c438ea1470a17687|1.0|2015-01-30 12:27:00|80.7095026033777|1||157|35.139506218778173|0|51|565|-80.661096|64|35.172688|REDUCED PRODUCE|0.0|4|PRODUCE REWRAP BY CT|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00204845000007|FRESH PRODUCE|PRODUCE|-80.709466|80.709478719700101|474|1
35.124987|c821a0ee093ee24d2bf241a5bd47cf9adfc26cb1|14.2|2015-02-13 14:11:00|1.4091206135396188|1|3620001401|157|0.6130466728702054|0|47|1221|-80.709466|275|35.124987|PASTA SC VALUE|0.0|1|RAGU SC 45 OWS WITH MEAT|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00036200014110|PASTA SAUCES|G1 GROCERY|-80.709466|1.4086459192264178|157|4
35.124987|1747aa2afc3fb86c06780b6aad783a6bce9ec79d|4.29|2015-02-06 17:43:00|1.4091206135396188|1|2840015938|157|0.6130466728702054|0|47|201|-80.709466|31|35.124987|POTATO CHIPS|1.79|1|XXL RUFFLES SR CRM & ONION|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00028400159630|SNACKS|G1 GROCERY|-80.709466|1.4086459192264178|157|1
35.124987|86fab30bd08f2aa5a2d845da69462bc2f89e9324|10.58|2015-01-18 15:14:00|80.7095026033777|1|7104000015|157|35.139506222092137|0|51|332|-80.654118|52|35.123768|STRING/SNACK|2.6|3|POLLY-O-TWISTARELLAS|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00071040065311|CHEESE|DAIRY|-80.709466|80.709470232147311|473|2
35.124987|6c5f93d99be2828f24a542c39fdb0a11fd12a152|13.29|2015-01-31 11:03:00|1.4091206135396188|1|3700013882|157|0.6130466728702054|0|47|389|-80.709466|66|35.124987|NFS-LAUNDRY DETERGENTS|1.3|1|TIDE ORIGINAL 64LD|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00037000138822|DETERGENTS|G1 GROCERY|-80.709466|1.4086459192264178|157|1
35.124987|d12935ffdfa51e2c5f821d35aeadeef450aaea7f|6.98|2014-10-21 13:13:00|80.7095026033777|1|3600038587|157|35.139506220647377|0|51|426|-80.70901|72|35.17335|NFS-PAPER TOWELS|1.0|1|KLEENEX HAND TOWEL WHITE|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00036000385878|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.709466|80.709474979800646|174|2
35.124987|8f2440aa1369497e426d61c64ff4079347f4bd1f|4.29|2014-11-29 18:45:00|1.4091206135396188|1|2840016014|157|0.6130466728702054|0|47|201|-80.709466|31|35.124987|POTATO CHIPS|0.29|1|LAYS WAVY REGULAR|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00028400160209|SNACKS|G1 GROCERY|-80.709466|1.4086459192264178|157|1
35.124987|593c65452d9d25d3cbe19838a4f467c94d0b5c13|1.19|2015-03-03 13:41:00|80.7095026033777|1|7203698213|157|35.139506222092137|0|51|257|-80.654118|39|35.123768|TOMATOES|0.0|1|HT TOMATOES DICED FIRE RST GAR|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00072036982148|VEGETABLES-CAN/JAR|G1 GROCERY|-80.709466|80.709470232147311|473|1
35.124987|ef622cdfec53426719c5a7db7c35eb23f227c947|10.99|2014-09-16 14:50:00|80.7095026033777|1|7203683001|157|35.139506222092137|0|51|352|-80.654118|110|35.123768|IQF CHICKEN|3.01|19|HT 2.5 LB CHICKEN TENDR BRST|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00072036830029|FROZEN CASE MEAT|CASE READY MEATS|-80.709466|80.709470232147311|473|1
35.124987|480082621cfa69b22135eb711e6989144ca30eef|4.19|2015-01-11 11:26:00|80.7095026033777|1|38137003237|157|35.139506220647377|0|51|5182|-80.70901|1305|35.17335|BABY BATH PRODUCTS|1.69|17|JOHNSONS BABY WASH VAN-OATMEAL|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00381370040231|BABY HBC|HBC|-80.709466|80.709474979800646|174|1
35.124987|c718452081c858b0650ca2268daaff9c9dd64e20|4.29|2015-01-03 15:45:00|1.4091206135396188|1|2840016014|157|0.6130466728702054|0|47|201|-80.709466|31|35.124987|POTATO CHIPS|2.15|1|LAYS CLASSIC|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00028400160148|SNACKS|G1 GROCERY|-80.709466|1.4086459192264178|157|1
35.124987|03d9470a29b41acbada949447f8ea38bb284a236|1.75|2014-09-21 11:53:00|1.4091206135396188|1|3120001605|157|0.6130466728702054|0|47|106|-80.709466|16|35.124987|CRANBERRY SAUCE|0.0|1|OS CRANBERRY SC WHOLE|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00031200016034|FRUIT-CAN/JAR|G1 GROCERY|-80.709466|1.4086459192264178|157|1
35.124987|9f8fb17b47f4e08c960698f2d5a5580f891e1639|4.29|2014-10-03 13:22:00|1.4091206135396188|1|2840016014|157|0.6130466728702054|0|47|201|-80.709466|31|35.124987|POTATO CHIPS|2.15|1|LAYS CLASSIC|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00028400160148|SNACKS|G1 GROCERY|-80.709466|1.4086459192264178|157|1
35.124987|4133fd53b96878bdb0908a63e0473f4cb5f39238|2.19|2014-09-21 11:51:00|1.4091206135396188|1|4900005010|157|0.6130466728702054|0|47|55|-80.709466|8|35.124987|REGULAR|0.2|23|SPRITE  2 LITER|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00049000050158|CARBONATED BEVERAGES|BEVERAGE|-80.709466|1.4086459192264178|157|1
35.124987|1484d1b82412e630f397e759fd9a7d9932b683c5|2.99|2015-01-06 18:44:00|80.7095026033777|1|7127913204|157|35.139506222092137|0|51|555|-80.654118|64|35.123768|PACKAGED SALADS|0.0|4|F.E. FLAT LEAF SPINACH,PKG|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00071279132044|FRESH PRODUCE|PRODUCE|-80.709466|80.709470232147311|473|1
35.124987|75957b77cf008315d3c0063400a2a234600f30ab|5.99|2015-02-03 13:44:00|80.7095026033777|1|7203688103|157|35.139506220647377|0|51|562|-80.70901|64|35.17335|FRESH CUT FRUIT|0.0|4|HT WATERMELON CHUNKS 32OZ|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00072036881038|FRESH PRODUCE|PRODUCE|-80.709466|80.709474979800646|174|1
35.124987|153d73dde2f2dae1c213efdd026c840d06668099|5.88|2014-09-29 15:01:00|1.4091206135396188|1|74759930652|157|0.6130466728702054|0|47|62|-80.709466|7|35.124987|SPECIALTY BAR/BOX CHOCOLATE|0.0|1|GHIRADELLI DARK CHOC RASP SQ|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00747599306532|CANDY|G1 GROCERY|-80.709466|1.4086459192264178|157|4
35.124987|b5636440a9ede5c9e9177b323ce433da8559b0f9|7.9|2014-11-30 12:04:00|1.4091206135396188|1|4450097650|157|0.6130466728702054|0|47|840|-80.709466|102|35.124987|TUBS|0.0|19|HF BOLD TUSCAN TURKEY|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00044500329544|LUNCHMEATS|CASE READY MEATS|-80.709466|1.4086459192264178|157|2
35.124987|f6418d46b8af9474214e05d82fef3e078b41338e|5.3|2015-01-17 17:16:00|1.4091206135396188|1|8768400095|157|0.6130466728702054|0|47|121|-80.709466|20|35.124987|ASEPTIC JUICES|0.3|1|CAPRI SUN FRUIT PUNCH 10 PK|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00087684001073|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.709466|1.4086459192264178|157|2
35.124987|589f49c17aa8733ee172ae0e1be435b45ace3fa3|4.89|2014-09-22 12:49:00|1.4091206135396188|1|20337400000|157|0.6130466728702054|0|47|641|-80.709466|137|35.124987|PREMIUM PORK|2.23|2|PORK LOIN BNLS BUTTERFLY CHOPS|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00203382000006|PORK|MEAT|-80.709466|1.4086459192264178|157|1
35.124987|547fcc1b4efcc2d688db51348eb39ca27c304a99|2.85|2014-11-19 12:10:00|80.7095026033777|1|4400000055|157|35.139506222092137|0|51|88|-80.654118|13|35.123768|FLAKED SODA CRACKERS|0.35|1|NABISCO PREMIUMS|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00044000000578|CRACKERS|G1 GROCERY|-80.709466|80.709470232147311|473|1
35.124987|0b33b4cb3b82ef189d6a9210c0f3a744b7b9423f|4.29|2015-02-21 10:24:00|80.7095026033777|1|7590000542|157|35.139506220647377|0|51|1271|-80.70901|41|35.17335|PROTEIN BREAKFAST|2.3|5|B EVANS HARVEST BURRITO 6CT|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00075900007480|BREAKFAST FOODS FROZEN|FROZEN|-80.709466|80.709474979800646|174|1
35.124987|05972163abbeff8bf4c0bf04ce8311b4e57e05f6|2.57|2015-02-14 08:14:00|80.7095026033777|1|5150055003|157|35.139506220647377|0|51|228|-80.70901|36|35.17335|TABLE SYRUP|0.0|1|HUNGRY JACK BUTR PANCAKE SYRUP|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00051500550052|TABLE SYRUPS|G1 GROCERY|-80.709466|80.709474979800646|174|1
35.124987|60d5f610a2951231456711bde5f41b3d8e8e5745|4.49|2014-11-21 19:02:00|80.7095026033777|1|6843738350|157|35.139506186146114|0|51|46|-80.782849|7|35.372142|PKG CHOC|0.5|1|BROOKSDE GOJI RASPBRY|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00068437383509|CANDY|G1 GROCERY|-80.709466|80.709505730947626|122|1
35.124987|1a151dec56f8e9e95f6bd15e9b8e229fcfad9372|2.97|2015-01-24 11:51:00|80.7095026033777|1|7106801126|157|35.139506222092137|0|51|1277|-80.654118|279|35.123768|FROZEN SNACKS|0.0|5|STATE FAIR CLASSIC CORN DOGS|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00071068011260|FROZEN SANDWICH AND SNACKS|FROZEN|-80.709466|80.709470232147311|473|1
35.124987|9a034d7db57f359d2173095ef1451e1511313692|9.69|2014-11-16 12:50:00|80.7095026033777|1|3700086527|157|35.139506222495768|0|51|427|-80.739|72|35.141204|NFS-TOILET TISSUE|1.7|1|CHARMIN BATH SENSITIVE 6MR|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00037000857365|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.709466|80.709466621902877|171|1
35.124987|8510e09f9676f379ce63262f2a87741005b6cbdb|11.97|2014-09-22 14:31:00|1.4091206135396188|1|7203697777|157|0.6130466728702054|0|47|31|-80.709466|4|35.124987|NON CARBONATED WATER|3.1599999999999997|1|(U) HT PURIFIED WATER 24 PK|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00072036977779|BOTTLED WATER|G1 GROCERY|-80.709466|1.4086459192264178|157|3
35.124987|b18148d30533594d16289f44267b5f4d8010c292|1.29|2015-02-14 08:15:00|80.7095026033777|1|7203670688|157|35.139506220647377|0|51|4816|-80.70901|1235|35.17335|FIRST AID ADHESIVE BANDG|0.0|17|HT BUTTERFLY CLOSURE ADH STRIP|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00072036706881|FIRST AID|HBC|-80.709466|80.709474979800646|174|1
35.124987|f76e11b48a8dff442c85e26343e6b4243e7f6d98|1.19|2015-01-20 09:42:00|1.4091206135396188|1|4178900301|157|0.6130466728702054|0|47|1203|-80.709466|33|35.124987|RAMEN|0.19|1|MARUCHAN BOWL HOT SPICY SHRIMP|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00041789003035|SOUP|G1 GROCERY|-80.709466|1.4086459192264178|157|1
35.124987|fd3d9c7b633b7cb0a08dc88ff0dd135d5a20921f|3.59|2015-02-11 09:04:00|80.7095026033777|1|4000024906|157|35.139506220647377|0|51|46|-80.70901|7|35.17335|PKG CHOC|0.0|1|M&M DARK CHOC PEANUT|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00040000236153|CANDY|G1 GROCERY|-80.709466|80.709474979800646|174|1
35.124987|16eb5d13e14acebecbe2c4f711f6e394e131b7c5|0.97|2015-01-10 12:41:00|1.4091206135396188|1|4300020431|157|0.6130466728702054|0|47|94|-80.709466|14|35.124987|PUDDING MIXES|0.0|1|JELLO INST PUDDING LEMON|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00043000204405|DESSERTS/GELS/SYRUPS|G1 GROCERY|-80.709466|1.4086459192264178|157|1
35.124987|c5c99cd4374c445e4a2fabe36c64c4a01418bb96|6.49|2014-10-22 11:51:00|80.7095026033777|1|60308441449|157|35.139506220647377|0|51|3500|-80.70901|1045|35.17335|CONDITIONER-MID PRICE|1.5|17|S/T GARNR MARVELOUS OIL (DRY)|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00603084414499|HAIR & SCALP CARE|HBC|-80.709466|80.709474979800646|174|1
35.124987|b03ab7b562310f54892468963e231ca2f4f59a95|9.98|2014-12-03 12:34:00|80.7095026033777|1|6827493471|157|35.139506222495768|0|51|31|-80.739|4|35.141204|NON CARBONATED WATER|4.0|1|NESTLE PURE LIFE .5L 24PK|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00068274934711|BOTTLED WATER|G1 GROCERY|-80.709466|80.709466621902877|171|2
35.124987|99e47aff5f830afab635d105408aa749aa00e20c|8.58|2015-01-18 15:12:00|80.7095026033777|1|3663200827|157|35.139506222092137|0|51|276|-80.654118|45|35.123768|ICE MILK/SHERBET/YOGURT-FROZEN|0.0|5|DANNON OIKOS FZ YOGURT VANILLA|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00036632008275|ICE CREAM|FROZEN|-80.709466|80.709470232147311|473|2
35.124987|ff40e64e5120399c850e0829d847575b4f27445b|3.49|2015-03-03 20:21:00|80.7095026033777|1|7203663995|157|35.139506220647377|0|51|342|-80.70901|57|35.17335|FRESH MILK|0.0|3|HARRIS TEETER 2% MILK|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00072036639981|MILK|DAIRY|-80.709466|80.709474979800646|174|1
35.124987|d1a5cf95acd5f072400342c9240bef5346d31ebf|11.88|2014-10-20 18:54:00|1.4091206135396188|1|2100000718|157|0.6130466728702054|0|47|317|-80.709466|52|35.124987|CHUNK AND BAR CHEESE|0.0|3|CRACKER BARREL CC EXTRA SHARP|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|0.61242566243833529|00021000007189|CHEESE|DAIRY|-80.709466|1.4086459192264178|157|4
35.124987|b543b1e8cb3425e0c9e5d9847322fdcf04110540|95.91999999999999|2015-01-30 12:46:00|80.7095026033777|1|7203671254|157|35.139506220263463|0|51|62|-80.62331|7|35.140781|SPECIALTY BAR/BOX CHOCOLATE|88.0|1|I/O HTT ASSORTED CHOCOLATE BOX|3c754abc1012814f22aa2c758f021df14061bcc1|1.0032432124065245|35.154129163572591|00072036712547|CANDY|G1 GROCERY|-80.709466|80.709475864323025|39|8
35.318911|061595fb9e14b8633c9a5e1e3a0a3c6b19ae598a|2.27|2014-11-17 12:52:00|80.77969194620016|3|7203611029|167|35.335073702378473|0|20|55|-80.945176|8|35.323246|REGULAR|0.0|23|HT COLA 12PK|3fcd53e862e9df4614efff01106fcb6707f56b61|1.1168039773374832|35.345012799095393|00072036110299|CARBONATED BEVERAGES|BEVERAGE|-80.780702|80.780715890081439|166|1
35.318911|cbf4771ae5e9a00c12d0635fccd81819556c6fc3|4.79|2014-12-27 16:11:00|80.77969194620016|3|7203611029|167|35.335073702378473|0|20|55|-80.945176|8|35.323246|REGULAR|1.79|23|HT COLA 12PK|3fcd53e862e9df4614efff01106fcb6707f56b61|1.1168039773374832|35.345012799095393|00072036110299|CARBONATED BEVERAGES|BEVERAGE|-80.780702|80.780715890081439|166|1
35.318911|743baf64841f7fad464a2d291c31b7c8396427d0|2.27|2014-10-06 20:59:00|80.77969194620016|3|7203611029|167|35.335073702378473|0|20|55|-80.945176|8|35.323246|REGULAR|0.27|23|HT COLA 12PK|3fcd53e862e9df4614efff01106fcb6707f56b61|1.1168039773374832|35.345012799095393|00072036110299|CARBONATED BEVERAGES|BEVERAGE|-80.780702|80.780715890081439|166|1
35.318911|35ebc853e485b88ae4cc9130dfa691b9854c1faa|2.27|2014-11-30 12:32:00|80.77969194620016|3|7203611029|167|35.335073702378473|0|20|55|-80.945176|8|35.323246|REGULAR|0.0|23|HT COLA 12PK|3fcd53e862e9df4614efff01106fcb6707f56b61|1.1168039773374832|35.345012799095393|00072036110299|CARBONATED BEVERAGES|BEVERAGE|-80.780702|80.780715890081439|166|1
35.318911|13eda644b12e30428f02ea5e0b82aee0465b14f7|4.49|2015-03-08 19:54:00|80.77969194620016|3|7203688080|167|35.335073702378473|0|20|523|-80.945176|64|35.323246|FRESH POTATOES|0.99|4|HT YUKON GOLD 5 LB BAG|3fcd53e862e9df4614efff01106fcb6707f56b61|1.1168039773374832|35.345012799095393|00072036880802|FRESH PRODUCE|PRODUCE|-80.780702|80.780715890081439|166|1
35.318911|ede0727020daa7a4945972ba8b3f191cb4940633|1.69|2014-11-01 14:25:00|80.77969194620016|3|7203688040|167|35.335073702378473|0|20|561|-80.945176|64|35.323246|FR PROD ORGANIC PRODUCE|0.0|4|ORG HT BABY CARROTS 1LB BAG|3fcd53e862e9df4614efff01106fcb6707f56b61|1.1168039773374832|35.345012799095393|00072036880406|FRESH PRODUCE|PRODUCE|-80.780702|80.780715890081439|166|1
35.318911|4994729f8c085ad73578d3869d213569aba5ffe6|5.99|2014-12-07 13:07:00|80.77969194620016|3|7203688215|167|35.335073702378473|0|20|500|-80.945176|64|35.323246|FRESH APPLES|0.0|4|HT GALA APPLE 5LB|3fcd53e862e9df4614efff01106fcb6707f56b61|1.1168039773374832|35.345012799095393|00072036882158|FRESH PRODUCE|PRODUCE|-80.780702|80.780715890081439|166|1
35.318911|06b14e88adb2a55ea6e552f7de71f7f13d43ce1d|3.49|2014-10-16 19:53:00|80.77969194620016|3|4400004557|167|35.335073705560816|0|20|89|-80.764523|12|35.341927|GRAHAM CRACKERS|0.99|1|TEDDY GRAHAMS CHOCOLATE CHIP|3fcd53e862e9df4614efff01106fcb6707f56b61|1.1168039773374832|35.345012799095393|00044000005979|COOKIES|G1 GROCERY|-80.780702|80.7807081959443|220|1
35.318911|e208df1055cce09ad2da0ed0ac5e5cf05642fc1b|3.59|2014-09-28 13:36:00|80.77969194620016|3|4850002013|167|35.335073702378473|0|20|335|-80.945176|56|35.323246|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA PP HOMESTYLE|3fcd53e862e9df4614efff01106fcb6707f56b61|1.1168039773374832|35.345012799095393|00048500301395|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.780702|80.780715890081439|166|1
35.318911|aabf764cd3a6b57ed1b448b472aabde53ad87793|2.29|2015-02-23 13:29:00|80.77969194620016|3|7203608066|167|35.335073702378473|0|20|1220|-80.945176|275|35.323246|PASTA SC PREMIUM|0.0|1|HTO PASTA SC TOM BASIL|3fcd53e862e9df4614efff01106fcb6707f56b61|1.1168039773374832|35.345012799095393|00072036080660|PASTA SAUCES|G1 GROCERY|-80.780702|80.780715890081439|166|1
35.318911|e290f7f16c00647e1d6f9bff19775445fce8264b|4.89|2014-11-10 15:22:00|80.77969194620016|3|2190874331|167|35.335073702378473|0|20|61|-80.945176|9|35.323246|RTE CEREAL ADULT|0.0|1|CASCADIAN ORG CINNAMON CRUNCH|3fcd53e862e9df4614efff01106fcb6707f56b61|1.1168039773374832|35.345012799095393|00021908455563|CEREAL|G1 GROCERY|-80.780702|80.780715890081439|166|1
35.318911|ce81d90eb0b70bc22daa383f75dfc0315de2b9f0|5.27|2014-10-16 19:54:00|80.77969194620016|3||167|35.335073705560816|0|20|501|-80.764523|64|35.341927|FRESH PEARS|0.53|4|BARTLETT PEARS|3fcd53e862e9df4614efff01106fcb6707f56b61|1.1168039773374832|35.345012799095393|00204409000009|FRESH PRODUCE|PRODUCE|-80.780702|80.7807081959443|220|1
35.318911|4805ea9b3e806d1bf813043ebd6ce3bfeb2508db|5.79|2014-12-31 15:23:00|80.77969194620016|3|81655901009|167|35.335073705560816|0|20|429|-80.764523|73|35.341927|NFS-BAR SOAP|2.9|1|ZEST COCOA BUTTR&SHEA BAR SOAP|3fcd53e862e9df4614efff01106fcb6707f56b61|1.1168039773374832|35.345012799095393|00816559012513|PERSONAL SOAP/BATH ADDITIVES|G1 GROCERY|-80.780702|80.7807081959443|220|1
35.318911|5d9919c8041e2ee1a3a33cb8c4da8fcfe10c2463|1.69|2014-09-12 18:21:00|80.77969194620016|3|1200000159|167|35.335073706343273|0|20|31|-80.737839|4|35.297134|NON CARBONATED WATER|0.0|1|CB AQUAFINA WATER 20 OZ|3fcd53e862e9df4614efff01106fcb6707f56b61|1.1168039773374832|35.345012799095393|00012000001598|BOTTLED WATER|G1 GROCERY|-80.780702|80.780702625553033|258|1
35.318911|2d5750f67ac05c55969cc61144d7ede1a6a13574|7.98|2014-11-06 13:03:00|80.77969194620016|3|71279710059|167|35.335073702378473|0|20|335|-80.945176|56|35.323246|ORANGE JUICE-REGRIGERATED|0.99|3|INDIAN RIVER ORANGE JUICE|3fcd53e862e9df4614efff01106fcb6707f56b61|1.1168039773374832|35.345012799095393|00712797100596|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.780702|80.780715890081439|166|2
35.318911|50f7aa4f7f8fd0359d8d777279e7f1c4c6e00475|4.49|2014-12-20 10:13:00|80.77969194620016|3|71279710059|167|35.335073702378473|0|20|335|-80.945176|56|35.323246|ORANGE JUICE-REGRIGERATED|0.0|3|INDIAN RIVER ORANGE JUICE|3fcd53e862e9df4614efff01106fcb6707f56b61|1.1168039773374832|35.345012799095393|00712797100596|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.780702|80.780715890081439|166|1
35.318911|de7f6be0dd99def674c9004ae631acdce15ddb85|2.49|2015-01-16 22:55:00|80.77969194620016|3|7535511228|167|35.335073706343273|0|20|139|-80.737839|20|35.297134|REMAINING SHELF STABLE JUICES|0.0|1|HEALTHY BALANCE POME/BLUE/ACAI|3fcd53e862e9df4614efff01106fcb6707f56b61|1.1168039773374832|35.345012799095393|00075355111756|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.780702|80.780702625553033|258|1
35.318911|d7e7865610dae48976d6668ce5566f06077b754f|1.0|2014-11-21 17:42:00|80.77969194620016|3|4000000435|167|35.335073703699521|0|20|47|-80.86175|7|35.40953|REGISTER BARS|0.2|1|(FE)3-MUSKETEER BARS|3fcd53e862e9df4614efff01106fcb6707f56b61|1.1168039773374832|35.345012799095393|00040000422082|CANDY|G1 GROCERY|-80.780702|80.780713348112769|209|1
35.318911|d5c95c13df8375efc181b64b15fa377171db3570|3.89|2015-01-16 22:56:00|80.77969194620016|3|61126954602|167|35.335073706343273|0|20|97|-80.737839|8|35.297134|ENERGY DRINKS|0.0|23|CB RED BULL SF UPER SLEEK|3fcd53e862e9df4614efff01106fcb6707f56b61|1.1168039773374832|35.345012799095393|00611269546026|CARBONATED BEVERAGES|BEVERAGE|-80.780702|80.780702625553033|258|1
35.318911|5a0ed77a0696d4ed9858b8972bbb0189184b0b31|14.99|2015-01-16 22:55:00|80.77969194620016|3|7199031600|167|35.335073706343273|0|20|455|-80.737839|82|35.297134|DOMESTIC PREMIUM 12PK&>|0.0|16|COORS LIGHT 24PK 12OZ CAN|3fcd53e862e9df4614efff01106fcb6707f56b61|1.1168039773374832|35.345012799095393|00071990316006|DOMESTIC BEER|BEER|-80.780702|80.780702625553033|258|1
35.006282|f67798287888269e0e3de42c210117cfca025322|4.29|2014-11-06 11:14:00|1.4091206135396188|4|7373100241|60|0.6109748797816256|0|47|495|-80.562829|108|35.006282|NON REFRIGERATED|0.0|19|MISSION SUNDRIED TOMATO WRAP|42e25ccd5d3ad6d31455978ed9c8877c42d3d4df|10.180886772947384|0.61242566243833529|00073731002902|TORTILLAS|CASE READY MEATS|-80.562829|1.4060866207711706|60|1
35.006282|e8b4c3d2486375206d3a8c6e9e40ef1ea490caf7|6.99|2014-09-23 13:09:00|1.4091206135396188|4|61458362401|60|0.6109748797816256|0|47|663|-80.562829|154|35.006282|FISH FILLETS/STEAKS PKGD|0.0|12|WHOLE CLEANED SQUID|42e25ccd5d3ad6d31455978ed9c8877c42d3d4df|10.180886772947384|0.61242566243833529|00614583624012|FISH FILLETS/STEAKS|SEAFOOD|-80.562829|1.4060866207711706|60|1
35.006282|eb1f582ee6d1d086f0a4a77f75e5f04c66fbf4bf|24.18|2014-09-26 13:51:00|1.4091206135396188|4|20829200000|60|0.6109748797816256|0|47|660|-80.562829|154|35.006282|FISH FILLETS WILD CGHT|2.42|12|WC FRESH HADDOCK FILLETS (NO)|42e25ccd5d3ad6d31455978ed9c8877c42d3d4df|10.180886772947384|0.61242566243833529|00208292000009|FISH FILLETS/STEAKS|SEAFOOD|-80.562829|1.4060866207711706|60|1
35.006282|559bf805d1326585b5dcbfd9e55c5a128cef8021|13.29|2014-11-14 14:47:00|1.4091206135396188|4|20829200000|60|0.6109748797816256|0|47|660|-80.562829|154|35.006282|FISH FILLETS WILD CGHT|1.33|12|WC FRESH HADDOCK FILLETS (NO)|42e25ccd5d3ad6d31455978ed9c8877c42d3d4df|10.180886772947384|0.61242566243833529|00208292000009|FISH FILLETS/STEAKS|SEAFOOD|-80.562829|1.4060866207711706|60|1
35.006282|deb26ae20cc6fff3dcef25cd05d81c9b638770d0|2.99|2015-02-13 13:51:00|1.4091206135396188|4|3338322235|60|0.6109748797816256|0|47|504|-80.562829|64|35.006282|FRESH BERRIES|0.0|4|BLUEBERRIES PINT|42e25ccd5d3ad6d31455978ed9c8877c42d3d4df|10.180886772947384|0.61242566243833529|00033383222011|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|1
35.006282|783cc6f069e9b1f132c64896dd002161f18afe34|19.96|2014-12-24 09:48:00|1.4091206135396188|4|20931900000|60|0.6109748797816256|0|47|676|-80.562829|148|35.006282|TAILS|0.0|12|WC LOBSTER TAILS 2/3 OZ  (CA)|42e25ccd5d3ad6d31455978ed9c8877c42d3d4df|10.180886772947384|0.61242566243833529|00209319000002|LOBSTERS|SEAFOOD|-80.562829|1.4060866207711706|60|1
35.006282|e10be19eddfe92d62a830195913a47b2d3a765dc|2.89|2014-10-24 14:38:00|1.4091206135396188|4|7203695174|60|0.6109748797816256|0|47|1625|-80.562829|373|35.006282|FROZEN DOUGH (ROLLS)|0.0|14|FRESH KAISER ROLLS 4 CT.|42e25ccd5d3ad6d31455978ed9c8877c42d3d4df|10.180886772947384|0.61242566243833529|00072036951748|ROLLS|BAKERY|-80.562829|1.4060866207711706|60|1
35.297134|6defd07ee01c8aa42046ba0cd49cd7df512e24e4|3.49|2014-12-27 21:19:00|1.4094857484078087|4|7203671181|258|0.6160512048176361|0|26|252|-80.737839|45|35.297134|PREMIUM ICE CREAM|0.49|5|HT RASPBERRY SHERBET|439c7f21faa78a615cc53a154488a9b45b19fded|1.369106876849274|0.61471665291522548|00072036711830|ICE CREAM|FROZEN|-80.737839|1.409141121495086|258|1
35.096737|4df0102a60ddd7d29b6b40b382a47f57256f27d1|2.85|2015-02-12 08:53:00|80.782094729586973|2|1920002522|30|35.112280194021089|0|27|404|-80.826724|69|35.195689|NFS-TOILET BOWL CLEANERS|0.0|1|LYSOL TOILET CLEANER CLING GEL|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00019200768788|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.78468|80.784695950319431|412|1
35.096737|3bf30e0d6c87beeb61099bc037e58e27cb19b118|4.99|2014-11-09 12:42:00|80.782094729586973|2|2840015297|30|35.112280194021089|0|27|204|-80.826724|31|35.195689|TORTILLA CHIPS|1.0|1|DORITOS NACHO CHEES PARTY SIZE|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00028400152976|SNACKS|G1 GROCERY|-80.78468|80.784695950319431|412|1
35.096737|8e319a3426a6e0870a27c232cf40c5ddbb6b7869|3.25|2014-11-23 14:56:00|80.782094729586973|2|3120020007|30|35.11228019496712|0|27|130|-80.80146|20|35.17739|CRANBERRY JUICE/DRINKS-SHELF|0.0|1|OSPRAY CRANBERRY JUICE|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00031200200075|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.78468|80.784694507674686|208|1
35.096737|132cc5aa5a0f6f960252f134b0e304451caa9878|2.5|2015-02-01 11:54:00|80.782094729586973|2|7203697755|30|35.11228019496712|0|27|74|-80.80146|9|35.17739|RTE CEREAL ALL FAMILY|0.71|1|HT CER CRISPY RICE|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00072036978509|CEREAL|G1 GROCERY|-80.78468|80.784694507674686|208|1
35.096737|b1279b4a8e072eafb480bfa0449fec2b287c5492|3.29|2015-01-11 15:33:00|80.782094729586973|2|7203688004|30|35.112280194021089|0|27|527|-80.826724|64|35.195689|FRESH CARROTS|0.0|4|HT BABY CARROTS 2LB BAG|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00072036880048|FRESH PRODUCE|PRODUCE|-80.78468|80.784695950319431|412|1
35.096737|c0b501641901d5d93d2745d40c8bc5630606df82|11.96|2014-12-24 09:22:00|80.782094729586973|2|3915310140|30|35.112280194021089|0|27|214|-80.826724|33|35.195689|BROTH|0.49|1|RACHAEL RAY CHCK LOW SOD STOCK|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00039153101449|SOUP|G1 GROCERY|-80.78468|80.784695950319431|412|4
35.096737|7a048e0b9c1a8dbeffc33423ea769ede225b56ea|5.98|2014-12-23 20:17:00|80.782094729586973|2|3915310140|30|35.112280194021089|0|27|214|-80.826724|33|35.195689|BROTH|0.98|1|RACHAEL RAY CHCK LOW SOD STOCK|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00039153101449|SOUP|G1 GROCERY|-80.78468|80.784695950319431|412|2
35.096737|5f6cc3bd9e10cbdb0557f2b03cba5588eaecee58|4.69|2015-01-17 16:37:00|80.782094729586973|2|5210000236|30|35.112280194021089|0|27|1245|-80.826724|34|35.195689|SINGLE SPICES|0.0|1|MC CREAM OF TARTAR|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00052100002361|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.78468|80.784695950319431|412|1
35.096737|096aca354714ad395a7e367c3bb87669aa543603|3.29|2014-09-15 11:06:00|80.782094729586973|2|61144334026|30|35.112280194021089|0|27|214|-80.826724|33|35.195689|BROTH|0.0|1|KITCHEN BASICS STOCK CHICKEN|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00611443340013|SOUP|G1 GROCERY|-80.78468|80.784695950319431|412|1
35.096737|6331b64f61a2691e99f814227521ae8335db4b11|1.69|2015-01-30 19:14:00|80.782094729586973|2|3660207290|30|35.112280194021089|0|27|4207|-80.826724|1200|35.195689|COUGH DROP-ADULT|0.0|17|RICOLA ECH. HONEY LEMN -30146|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00036602301467|COUGH/COLD/SINUS|HBC|-80.78468|80.784695950319431|412|1
35.096737|4b614616c7ddeb91fade2916b74cf7a91ad52bbe|1.27|2014-12-06 11:52:00|80.782094729586973|2|7203603051|30|35.112280197337974|0|27|29|-80.85013|3|35.175855|REMAINING BAKING SUPPLIES|0.0|1|HT BAKING POWDER|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00072036030511|BAKING SUPPLIES|G1 GROCERY|-80.78468|80.78469001773837|218|1
35.096737|da8f71b7af69da0cd498995a0556f6bd76fa4f09|27.99|2015-03-04 12:55:00|80.782094729586973|2|31284354120|30|35.112280194021089|0|27|4451|-80.826724|1210|35.195689|PROBIOTICS|0.0|17|PHILLIPS COLON HEALTH CAPS|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00312843541207|STOMACH REMEDIES|HBC|-80.78468|80.784695950319431|412|1
35.096737|8b5bacf093bcdc06dd125d4a2e3888410c603ce8|25.810000000000002|2014-10-12 15:57:00|80.782094729586973|2|20899100000|30|35.112280194021089|0|27|1421|-80.826724|201|35.195689|SMART CHICKEN VEGETABLE FED|0.0|2|SMART CHICKEN BREAST TENDERS|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00208991000003|POULTRY|MEAT|-80.78468|80.784695950319431|412|2
35.096737|1f7bf175bfd347e4340a33e04f9aad371f746de8|25.98|2015-02-16 15:07:00|80.782094729586973|2|7203695587|30|35.112280194021089|0|27|1707|-80.826724|387|35.195689|MESSAGE|6.0|14|12 INCH MESSAGE COOKIE|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00072036955876|COOKIES|BAKERY|-80.78468|80.784695950319431|412|2
35.096737|6cac2e6995d67f6759a0dd9101af0348d8139d82|3.0|2014-09-20 16:33:00|80.782094729586973|2|7203688157|30|35.112280194021089|0|27|556|-80.826724|64|35.195689|PACKAGED VEGETABLES|0.0|4|HT RV BABY ZUCCHINI SQUASH|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00072036881571|FRESH PRODUCE|PRODUCE|-80.78468|80.784695950319431|412|1
35.096737|c614f357b03310e3166802adb975adca17807614|3.79|2015-02-15 15:53:00|80.782094729586973|2|4950800600|30|35.112280194021089|0|27|1981|-80.826724|480|35.195689|CHIPS|0.0|6|MINI CHEDDAR PRETZEL CRISPS|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00049508002178|DRY GOODS|DELI|-80.78468|80.784695950319431|412|1
35.096737|b593cbfccb2d448ad29ff1346f619b4f6bb7b40b|4.76|2014-10-19 12:56:00|80.782094729586973|2|3940001747|30|35.112280194021089|0|27|242|-80.826724|39|35.195689|CANNED BEANS|0.19|1|BUSH BEAN RS DK KIDNEY|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00039400017301|VEGETABLES-CAN/JAR|G1 GROCERY|-80.78468|80.784695950319431|412|4
35.096737|29fb52e04655505cf890bfdc80f0272b225db1a8|8.89|2014-11-08 14:35:00|80.782094729586973|2|1410009655|30|35.112280194021089|0|27|87|-80.826724|13|35.195689|CHEESE CRACKERS|0.9|1|PF BULK GOLDFISH CHEDDAR|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00014100096559|CRACKERS|G1 GROCERY|-80.78468|80.784695950319431|412|1
35.096737|98fca5b5212ca1a25a05fded969164e97f073801|10.99|2014-10-18 16:35:00|80.782094729586973|2|74052210083|30|35.112280194021089|0|27|458|-80.826724|82|35.195689|CRAFT BEER|0.0|16|BELL'S 2 HEARTED ALE 6PK|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00740522100832|DOMESTIC BEER|BEER|-80.78468|80.784695950319431|412|1
35.096737|608f5a0ffd69e36a5b4055a22f2ca1e4f6013843|2.99|2015-02-16 08:47:00|80.782094729586973|2|7027223202|30|35.112280194021089|0|27|323|-80.826724|57|35.195689|TOPPINGS-REFRIGERATED|0.49|3|REDDI WIP EXTRA CREAMY|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00070272232034|MILK|DAIRY|-80.78468|80.784695950319431|412|1
35.096737|3c2557993ed7063205e572092830e573912c6480|7.99|2015-03-08 19:21:00|80.782094729586973|2|7027710518|30|35.112280194021089|0|27|2020|-80.826724|505|35.195689|CHEESE SPECIALTIES|0.0|6|ATHENOS FETA TRADITIONAL CHUNK|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00070277105180|SPECIALTY CHEESE|DELI|-80.78468|80.784695950319431|412|1
35.096737|a3cb416210d623e18c403ac409da6a6e4fad3c84|16.99|2015-02-01 15:46:00|80.782094729586973|2|18195400004|30|35.112280194021089|0|27|459|-80.826724|83|35.195689|IMPORT BEER|0.0|16|PERONI 12PK|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00181954000046|IMPORT BEER|BEER|-80.78468|80.784695950319431|412|1
35.096737|1bde11297b892ff896d627779f59675876d58705|4.59|2015-01-20 19:32:00|80.782094729586973|2|1862729292|30|35.112280199382489|0|27|1278|-80.85753|48|35.116638|SINGLE SERVE NUTRITIONAL|0.0|5|KASHI PESTO PASTA PRIMAVERA|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00018627292906|FROZEN MEALS|FROZEN|-80.78468|80.784682322579258|204|1
35.096737|2fc878d0336ae3b836e6098f20dae3a7b7e7dad2|4.29|2014-09-19 17:37:00|80.782094729586973|2|2840015636|30|35.11228019496712|0|27|204|-80.80146|31|35.17739|TORTILLA CHIPS|0.0|1|DORTIOS NACHO CHEESE|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00028400156363|SNACKS|G1 GROCERY|-80.78468|80.784694507674686|208|1
35.096737|1f8da969c57f6272ccf86a3f981866a8722a068e|3.79|2014-11-27 10:49:00|80.782094729586973|2|2500005542|30|35.112280194021089|0|27|335|-80.826724|56|35.195689|ORANGE JUICE-REGRIGERATED|0.0|3|SIMPLY ORANGE ORIGINAL|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00025000055423|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.78468|80.784695950319431|412|1
35.096737|c2c1186d748fa1a4525d13cb5220f507ac171940|8.49|2015-01-25 18:21:00|80.782094729586973|2|2737140002|30|35.112280194021089|0|27|5864|-80.826724|1538|35.195689|STERNO FUEL|0.0|18|7OZ STERNO 2PK COOKING FUEL|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00027371400024|KITCHEN GADGETS|GM|-80.78468|80.784695950319431|412|1
35.096737|d8e5de9e143fd28c8cb3e2b2a0e62e32db228057|4.99|2014-12-14 16:30:00|80.782094729586973|2|7203695160|30|35.112280194021089|0|27|1937|-80.826724|465|35.195689|COLD PREP FOODS ENTREES|0.0|6|PEPPERONI & CHEESE CALZONE|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00072036951601|COLD PREPARED FOODS|DELI|-80.78468|80.784695950319431|412|1
35.096737|a9efe02a1b4bbed1a4110f3b54cb7ff1964706a6|1.99|2014-11-09 12:44:00|80.782094729586973|2||30|35.112280194021089|0|27|274|-80.826724|44|35.195689|ICE|0.0|5|HT BAGGED ICE|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00072036480118|ICE|FROZEN|-80.78468|80.784695950319431|412|1
35.096737|63a1e8aaa5c659c224cfd19665950bc5d2813f06|8.95|2015-01-26 19:06:00|80.782094729586973|2|20690000000|30|35.112280194021089|0|27|2027|-80.826724|510|35.195689|SOMETHING CLASSIC|0.0|6|SOMETHING CLASSIC SOUPS|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00206900000007|SOMETHING CLASSIC|DELI|-80.78468|80.784695950319431|412|1
35.096737|315ad1438b60de0e14b01e53bf985307f89322df|2.79|2014-12-23 11:13:00|80.782094729586973|2|4400004833|30|35.112280194021089|0|27|27|-80.826724|3|35.195689|PIE & PASTRY SHELLS|0.3|1|NABISCO OREO PIE CRUST|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00044000048341|BAKING SUPPLIES|G1 GROCERY|-80.78468|80.784695950319431|412|1
35.096737|c4624f81bae27ad0223a149e2a950d5cfd2cceb7|2.99|2015-02-07 17:54:00|80.782094729586973|2|1800000338|30|35.112280194021089|0|27|1268|-80.826724|54|35.195689|BAGELS AND MUFFINS|0.0|3|PILLSBURY READY PIZZA CRUST|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00018000003389|DOUGH PRODUCTS|DAIRY|-80.78468|80.784695950319431|412|1
35.096737|527033d6ae2e58dd8ebc48e94a596bd187618ee3|2.34|2014-11-14 21:20:00|80.782094729586973|2||30|35.112280194021089|0|27|562|-80.826724|64|35.195689|FRESH CUT FRUIT|0.0|4|(SEEDLESS) WATERMELON CHUNKS|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00204485000009|FRESH PRODUCE|PRODUCE|-80.78468|80.784695950319431|412|1
35.096737|4b3065ce365af3c93a17eb03858e7846b0abaf2c|10.99|2014-11-26 12:48:00|80.782094729586973|2|78535701280|30|35.112280194021089|0|27|37|-80.826724|10|35.195689|PODS/CUPS/SINGLES|5.5|1|PEET'S 10CT BRAZIL MINAS NATUR|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00785357012653|COFFEE|G1 GROCERY|-80.78468|80.784695950319431|412|1
35.096737|e22e6a96a1d7b50918f4863a0949c6afaf426c93|6.0|2015-02-08 09:45:00|80.782094729586973|2|812|30|35.11228019496712|0|27|1639|-80.80146|377|35.17739|BULK (DONUTS)|0.0|14|NEW BULK DONUT CODE|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00000000008120|DONUTS|BAKERY|-80.78468|80.784694507674686|208|6
35.096737|e67bc94d5fbdb9825def35becb01eaa485084e0e|13.99|2014-11-24 17:52:00|80.782094729586973|2|8378322200|30|35.112280191914941|0|27|458|-80.850065|82|35.030252|CRAFT BEER|0.0|16|SIERRA NEVADA PALE ALE 12PK|442203e01a20a083b6bb6f5490a95092f8f74667|1.0739975498726126|35.102887530186244|00083783222005|DOMESTIC BEER|BEER|-80.78468|80.784698767950715|470|1
35.603432|a5ab7a4ccfebd68c635d84971f599f054bc3cc69|9.99|2015-01-18 17:26:00|80.891462859624312|4|4740012602|274|35.624652118127379|0|45|3917|-80.875654|1075|35.585842|DISPOSABLE RAZOE-MEN|2.0|17|GOODNEWS DISP RAZORS REGULAR|4798faeef2bb5f29d5463ff10993062955a83acf|1.4662589243268478|35.636605227883024|00047400125988|SHAVING NEEDS/MEN HAIR|HBC|-80.895009|80.895011453123558|99|1
35.603432|41a675ab7223fcb1f7f541d0c712211afd114b36|8.99|2015-01-29 16:06:00|80.891462859624312|4|7203688111|274|35.624652118127379|0|45|583|-80.875654|136|35.585842|NUTS|0.0|4|HT SLICED NATURAL ALMONDS,TRAY|4798faeef2bb5f29d5463ff10993062955a83acf|1.4662589243268478|35.636605227883024|00072036881113|OTHER MERCHANDISE|PRODUCE|-80.895009|80.895011453123558|99|1
35.603432|d8f28349a7e3958c301599cd7387ddbc741072f1|2.69|2014-09-24 17:12:00|80.891462859624312|4|7203663996|274|35.624652118127379|0|45|342|-80.875654|57|35.585842|FRESH MILK|0.0|3|HARRIS TEETER 2%   MILK|4798faeef2bb5f29d5463ff10993062955a83acf|1.4662589243268478|35.636605227883024|00072036639998|MILK|DAIRY|-80.895009|80.895011453123558|99|1
35.603432|ba57abb5c60ace2ba8c6dd57e67027ab8f2804fa|13.98|2014-11-24 18:36:00|80.891462859624312|4|76108880069|274|35.624652118127379|0|45|1939|-80.875654|465|35.585842|COLD PREP FOODS SIDES|0.0|6|MASHED POTATOES|4798faeef2bb5f29d5463ff10993062955a83acf|1.4662589243268478|35.636605227883024|00761088800691|COLD PREPARED FOODS|DELI|-80.895009|80.895011453123558|99|2
35.603432|dc676d7dbdacc81cea68b43b1420fb42889dd53b|1.2|2014-10-05 20:52:00|80.891462859624312|4|89470001004|274|35.624652118127379|0|45|685|-80.875654|61|35.585842|GREEK|0.0|3|CHOBANI NF BLUBERRY|4798faeef2bb5f29d5463ff10993062955a83acf|1.4662589243268478|35.636605227883024|00894700010052|YOGURT|DAIRY|-80.895009|80.895011453123558|99|1
35.603432|f5fbb43464faa8bd60b62383b1c091b8295998c9|2.55|2014-12-21 18:31:00|80.891462859624312|4|7203663996|274|35.624652118127379|0|45|342|-80.875654|57|35.585842|FRESH MILK|0.0|3|HARRIS TEETER 2%   MILK|4798faeef2bb5f29d5463ff10993062955a83acf|1.4662589243268478|35.636605227883024|00072036639998|MILK|DAIRY|-80.895009|80.895011453123558|99|1
35.603432|be99fbd526cf05fe6124f6a8944b1c9133ca3cbe|2.99|2014-11-10 17:44:00|80.891462859624312|4|4082202224|274|35.624652118127379|0|45|581|-80.875654|136|35.585842|FRESH SALSA|0.0|4|SABRA GUACAMOLE CLASSIC|4798faeef2bb5f29d5463ff10993062955a83acf|1.4662589243268478|35.636605227883024|00040822022248|OTHER MERCHANDISE|PRODUCE|-80.895009|80.895011453123558|99|1
35.603432|89a55066bba411dfd53cedd8ed91d3fd342915ee|3.74|2014-12-07 13:15:00|80.891462859624312|4|7203620120|274|35.624652118127379|0|45|139|-80.875654|20|35.585842|REMAINING SHELF STABLE JUICES|0.0|1|HT RECONSTITUTED LEMON JUICE|4798faeef2bb5f29d5463ff10993062955a83acf|1.4662589243268478|35.636605227883024|00072036201201|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.895009|80.895011453123558|99|2
35.116638|918d5cb4095bc7173daf48da7b35b6566b768cfd|8.98|2014-09-18 14:19:00|80.856688219393845|1|71575620002|204|35.131248911135707|0|15|504|-80.824767|64|35.116751|FRESH BERRIES|1.0|4|STRAWBERRIES 1LB CLAM|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00715756200023|FRESH PRODUCE|PRODUCE|-80.85753|80.857532666903609|294|2
35.116638|bbba43f4c5e3e28325df699672d62e0d16f18c7e|12.01|2014-12-20 13:45:00|1.4091206135396188|1||204|0.6129009553309565|0|47|561|-80.85753|64|35.116638|FR PROD ORGANIC PRODUCE|1.51|4|ORG HH BUNCH TOMATOES|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00294664000005|FRESH PRODUCE|PRODUCE|-80.85753|1.4112301235300906|204|1
35.116638|b94f644d7d34c329f2151e51ad0953c05e4632da|9.98|2015-03-08 09:11:00|1.4091206135396188|1|71575620002|204|0.6129009553309565|0|47|504|-80.85753|64|35.116638|FRESH BERRIES|4.98|4|STRAWBERRIES 1LB CLAM|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00715756200023|FRESH PRODUCE|PRODUCE|-80.85753|1.4112301235300906|204|2
35.116638|45ac049a2242ee138586818740cd5e81cd17eaae|3.99|2015-03-02 05:20:00|1.4091206135396188|1|85281048712|204|0.6129009553309565|0|47|330|-80.85753|55|35.116638|EGGS|0.0|3|LOL ALL NAT XL BROWN EGGS|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00852810487126|EGGS FRESH|DAIRY|-80.85753|1.4112301235300906|204|1
35.116638|76a22fee3ec9cfaf093afef3ab2d2ca2e1d99505|3.99|2014-12-29 16:19:00|80.856688219393845|1|3338324028|204|35.131248911135707|0|15|504|-80.824767|64|35.116751|FRESH BERRIES|0.99|4|BLACKBERRIES 6 OZ|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00891700002087|FRESH PRODUCE|PRODUCE|-80.85753|80.857532666903609|294|1
35.116638|7426273cbdb69141be47b9f9f30081d9165c8440|0.99|2014-11-10 18:12:00|80.856688219393845|1||204|35.13124890930947|0|15|540|-80.825175|64|35.152722|FRESH CELERY|0.0|4|COO CELERY (RPC) 24'S|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00204070000001|FRESH PRODUCE|PRODUCE|-80.85753|80.857539321200392|160|1
35.116638|e1be7dfb672afb5f668e2808a449cc0cb57c9f44|20.99|2014-11-26 16:42:00|1.4091206135396188|1|8751292795|204|0.6129009553309565|0|47|9964|-80.85753|887|35.116638|NFS-S/PREM-PINOT NOIR|0.0|13|RODNEY STRONG RR PINOT NOIR|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00087512927957|SUPER PREMIUM ($11-$14.99)|WINE|-80.85753|1.4112301235300906|204|1
35.116638|9122937d3e2a1525bc2321d647b7fc064b537884|20.99|2015-01-11 16:12:00|1.4091206135396188|1|8751292795|204|0.6129009553309565|0|47|9964|-80.85753|887|35.116638|NFS-S/PREM-PINOT NOIR|0.0|13|RODNEY STRONG RR PINOT NOIR|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00087512927957|SUPER PREMIUM ($11-$14.99)|WINE|-80.85753|1.4112301235300906|204|1
35.116638|2368d619aba51f9f7be37f8935e3eedb9e5780b2|6.98|2015-02-25 10:17:00|80.856688219393845|1|20455000000|204|35.13124890930947|0|15|542|-80.825175|64|35.152722|FRESH VEGETABLES REMAIN|0.0|4|BRUSSEL SPROUTS 1LB (RPC)|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00094922577160|FRESH PRODUCE|PRODUCE|-80.85753|80.857539321200392|160|2
35.116638|7492eec1fdfe255a3df6b3df5ad5442c5a32b49d|20.99|2014-11-22 16:07:00|1.4091206135396188|1|8751292795|204|0.6129009553309565|0|47|9964|-80.85753|887|35.116638|NFS-S/PREM-PINOT NOIR|0.0|13|RODNEY STRONG RR PINOT NOIR|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00087512927957|SUPER PREMIUM ($11-$14.99)|WINE|-80.85753|1.4112301235300906|204|1
35.116638|5989ae8b425f5ece05bcc021935801a1f4166d2f|3.49|2015-01-11 16:08:00|1.4091206135396188|1|20455000000|204|0.6129009553309565|0|47|542|-80.85753|64|35.116638|FRESH VEGETABLES REMAIN|0.0|4|BRUSSEL SPROUTS 1LB (RPC)|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00094922577160|FRESH PRODUCE|PRODUCE|-80.85753|1.4112301235300906|204|1
35.116638|7393f893c932977fb06dd7154e83f0ed0c856638|3.49|2015-02-05 20:01:00|80.856688219393845|1|7797508005|204|35.131248908216527|0|15|202|-80.85013|31|35.175855|PRETZELS|0.3|1|SOH SOURDOUGH HARD PRETZEL|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00077975080030|SNACKS|G1 GROCERY|-80.85753|80.857541602840982|218|1
35.116638|eb7354b1a707d2d9709cc105965d1a474b8364b7|7.49|2014-10-14 14:38:00|1.4091206135396188|1|7490836026|204|0.6129009553309565|0|47|1220|-80.85753|275|35.116638|PASTA SC PREMIUM|1.5|1|DELGROSSO SC MARINARA|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00074908360269|PASTA SAUCES|G1 GROCERY|-80.85753|1.4112301235300906|204|1
35.116638|ced1ccefd39eabf562383deeaab43aac887602a2|2.89|2014-12-12 12:51:00|1.4091206135396188|1|2409407012|204|0.6129009553309565|0|47|151|-80.85753|23|35.116638|DSD PASTA CORE|0.0|1|DE CECCO FETTUCCINE # 6|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00024094070060|PASTA|G1 GROCERY|-80.85753|1.4112301235300906|204|1
35.116638|56685e015c94d8c3b58ebb61e4e32020ddcb63aa|12.4|2014-10-09 21:33:00|80.856688219393845|1|2920000212|204|35.131248909433786|0|15|149|-80.849471|23|35.161696|WHSE PASTA CORE|0.0|1|MUELLER POT SZ SPAGHETTI|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00029200907964|PASTA|G1 GROCERY|-80.85753|80.857539025206648|35|8
35.116638|a5a796b5890e5736c05c5f64d67b27f5ba0e3651|4.99|2014-10-27 16:49:00|1.4091206135396188|1|2301290130|204|0.6129009553309565|0|47|1477|-80.85753|485|35.116638|SUSHI HYBRID|0.0|6|CALIFORNIA ROLL SP|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00023012901301|SUSHI|DELI|-80.85753|1.4112301235300906|204|1
35.116638|607c3ec9799be538ec5bf6ec638a845e78849e71|5.99|2014-11-08 08:05:00|1.4091206135396188|1|2301290165|204|0.6129009553309565|0|47|1477|-80.85753|485|35.116638|SUSHI HYBRID|0.0|6|VEGETABLE COMBO SP BRN RICE|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00023012901653|SUSHI|DELI|-80.85753|1.4112301235300906|204|1
35.116638|b57f659042b32f31d68a7fda8eccd2dbcf445ee8|3.99|2014-10-22 13:44:00|1.4091206135396188|1|1410007111|204|0.6129009553309565|0|47|1038|-80.85753|164|35.116638|SWIRL/TOASTING|0.0|7|PEP CINNAMON BREAD 16 OZ  PP|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00014100070610|BREAKFAST|COMMERCIAL BAKERY|-80.85753|1.4112301235300906|204|1
35.116638|0db9993f662cf60fa3fabee234e163d60eb0b876|2.69|2014-12-02 05:53:00|1.4091206135396188|1|1600026460|204|0.6129009553309565|0|47|42|-80.85753|6|35.116638|GRANOLA/YOGURT BARS|0.0|1|NV BAR CRN HONEY OATS|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00016000264601|BREAKFAST FOODS|G1 GROCERY|-80.85753|1.4112301235300906|204|1
35.116638|7b418d73d6a28fbb04a4f6d1d4b273b846b50a75|3.19|2015-02-20 11:29:00|80.856688219393845|1|74759961274|204|35.13124890439326|0|15|16|-80.844274|3|35.204336|BAKING CHOCOLATE/CHIPS/MORSELS|0.0|1|GHIRADELLI 60% BITTRSWEET CHIP|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00747599612749|BAKING SUPPLIES|G1 GROCERY|-80.85753|80.857547367555895|61|1
35.116638|5aabb9dca33ff7f46df19c14bd73a42bae9922f0|20.96|2014-09-21 17:47:00|80.856688219393845|1|20895300000|204|35.13124890439326|0|15|977|-80.844274|201|35.204336|FRESH HT CHICKEN|4.52|2|HT FRESH BNLS CHICKEN BREAST|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00208953000003|POULTRY|MEAT|-80.85753|80.857547367555895|61|2
35.116638|67a91a32459d590270f152f279f175d2ec7e41bf|10.23|2015-01-25 18:37:00|80.856688219393845|1|20895300000|204|35.131248909433786|0|15|977|-80.849471|201|35.161696|FRESH HT CHICKEN|0.0|2|HT FRESH BNLS CHICKEN BREAST|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00208953000003|POULTRY|MEAT|-80.85753|80.857539025206648|35|1
35.116638|d0d1b815d685ed061d758e1532795fe355d2eb14|3.29|2014-09-13 13:14:00|1.4091206135396188|1|71536440037|204|0.6129009553309565|0|47|71|-80.85753|11|35.116638|GROC CONDIMENTS MARINADE|0.0|1|D WRLD HRBR MARINADE SRIRACHA|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00715364400372|CONDIMENTS|G1 GROCERY|-80.85753|1.4112301235300906|204|1
35.116638|48c8e3b9fb86e64a51aa76059e69161bd30f2c23|2.99|2015-02-27 17:33:00|80.856688219393845|1|81204900640|204|35.131248911135707|0|15|504|-80.824767|64|35.116751|FRESH BERRIES|0.0|4|BLUEBERRIES 6 OZ|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00761635203906|FRESH PRODUCE|PRODUCE|-80.85753|80.857532666903609|294|1
35.116638|126f0824febfcf84210afc514c2b7c42c8cad71f|4.69|2015-01-05 16:13:00|80.856688219393845|1|1600043779|204|35.131248911135707|0|15|1433|-80.824767|9|35.116751|GRANOLA|0.0|1|NV PROTEIN GRANOLA OATS HONEY|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00016000437791|CEREAL|G1 GROCERY|-80.85753|80.857532666903609|294|1
35.116638|64f842d6aba8dd21b79a5735859586a290e9306c|2.89|2014-11-24 05:55:00|1.4091206135396188|1|1760004370|204|0.6129009553309565|0|47|247|-80.85753|39|35.116638|VEGETABLES-FLANKER|1.1|1|MARTINDALE SWEET POTATOES CUT|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00017600043702|VEGETABLES-CAN/JAR|G1 GROCERY|-80.85753|1.4112301235300906|204|1
35.116638|2afac534fb2f25518eba563e75b657df0dfd27e4|4.69|2014-11-09 17:27:00|80.856688219393845|1|1600043779|204|35.131248911135707|0|15|1433|-80.824767|9|35.116751|GRANOLA|0.0|1|NV PROTEIN GRANOLA OATS HONEY|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00016000437791|CEREAL|G1 GROCERY|-80.85753|80.857532666903609|294|1
35.116638|4754168c4aef19691d20a084fa9ca8b8d9088be9|2.99|2014-12-03 18:10:00|1.4091206135396188|1|20443000000|204|0.6129009553309565|0|47|510|-80.85753|64|35.116638|FRESH PINEAPPLE|0.0|4|GOLD PINEAPPLES|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00643126072003|FRESH PRODUCE|PRODUCE|-80.85753|1.4112301235300906|204|1
35.116638|7e9b17fdab0d1e1aa33874a8db959bd3bf514811|29.97|2014-11-23 15:45:00|1.4091206135396188|1|83299201011|204|0.6129009553309565|0|47|4237|-80.85753|1200|35.116638|MEDICATED LIP CARE|0.0|17|I/O EOS LP BLM RR COLL 3PK|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00832992010114|COUGH/COLD/SINUS|HBC|-80.85753|1.4112301235300906|204|3
35.116638|da6d2930a0f6bb159085580c851c5fc596b574c9|4.49|2015-02-03 19:39:00|80.856688219393845|1|7116915895|204|35.13124890439326|0|15|734|-80.844274|3|35.204336|NFS-CANDLES/BIRTHDAY SUP|0.0|1|CAKE MATE HAPPY BIRTHDAY CANDL|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00071169158956|BAKING SUPPLIES|G1 GROCERY|-80.85753|80.857547367555895|61|1
35.116638|1ad7f172aa429c950a375371d1459462cd43f16b|12.99|2014-11-26 11:48:00|80.856688219393845|1|7023666334|204|35.13124890930947|0|15|1153|-80.825175|87|35.152722|NFS-FRESH CUT ARRANGE|0.0|9|PETITE EXPRESSION ARR.|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00070236663348|FLORAL|FLORAL|-80.85753|80.857539321200392|160|1
35.116638|f926a57210f36a148916bff743975af0695fc02d|4.99|2014-11-21 17:01:00|80.856688219393845|1|4950800823|204|35.131248909433786|0|15|1980|-80.849471|480|35.161696|CHOCOLATES|1.0|6|DARK CHOC PRETZEL CRISPS|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00049508008231|DRY GOODS|DELI|-80.85753|80.857539025206648|35|1
35.116638|953182a08b180d5b760f17fd4aee23ac23258334|7.99|2014-09-30 07:44:00|80.856688219393845|1|68954408301|204|35.131248908216527|0|15|685|-80.85013|61|35.175855|GREEK|0.0|3|FAGE TOTAL 2%|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00689544083023|YOGURT|DAIRY|-80.85753|80.857541602840982|218|1
35.116638|4e86ac37111e61d728af3ba28fd5a51246ad5367|7.98|2014-11-15 10:06:00|80.856688219393845|1|20405400000|204|35.131248911135707|0|15|504|-80.824767|64|35.116751|FRESH BERRIES|2.0|4|RED RASPBERRIES 6 OZ|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00715756100019|FRESH PRODUCE|PRODUCE|-80.85753|80.857532666903609|294|2
35.116638|5df18787fd2213bba9f95b1869074112bbe092cc|5.99|2014-10-13 11:35:00|80.856688219393845|1|76108880156|204|35.131248911135707|0|15|1939|-80.824767|465|35.116751|COLD PREP FOODS SIDES|0.0|6|MACARONI & CHEESE FAMILY SIZE|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00761088801568|COLD PREPARED FOODS|DELI|-80.85753|80.857532666903609|294|1
35.116638|b3d7ba50397920d9aab74f4f9da5b63b9936e5e2|11.97|2014-09-28 18:18:00|80.856688219393845|1|20405400000|204|35.131248911135707|0|15|504|-80.824767|64|35.116751|FRESH BERRIES|6.970000000000001|4|RED RASPBERRIES 6 OZ|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00715756100019|FRESH PRODUCE|PRODUCE|-80.85753|80.857532666903609|294|3
35.116638|91eba45dee8b73e8926d3c79810fe0873f625724|7.98|2015-01-29 12:33:00|80.856688219393845|1|20405400000|204|35.13124890930947|0|15|504|-80.825175|64|35.152722|FRESH BERRIES|0.0|4|RED RASPBERRIES 6 OZ|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00715756100019|FRESH PRODUCE|PRODUCE|-80.85753|80.857539321200392|160|2
35.116638|7a031c5f0415f604acf51e7af26cd896454d0512|15.96|2014-11-05 11:32:00|80.856688219393845|1|20405400000|204|35.13124890930947|0|15|504|-80.825175|64|35.152722|FRESH BERRIES|7.470000000000001|4|RED RASPBERRIES 6 OZ|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00715756100019|FRESH PRODUCE|PRODUCE|-80.85753|80.857539321200392|160|4
35.116638|7780f9783c4625037182692b2341529949c356e8|3.99|2015-02-09 17:31:00|80.856688219393845|1|20405400000|204|35.131248909433786|0|15|504|-80.849471|64|35.161696|FRESH BERRIES|0.0|4|RED RASPBERRIES 6 OZ|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00715756100019|FRESH PRODUCE|PRODUCE|-80.85753|80.857539025206648|35|1
35.116638|03a0907ad4a2c8037b5202c47a1d51054c83149c|4.07|2014-12-03 12:18:00|1.4091206135396188|1||204|0.6129009553309565|0|47|561|-80.85753|64|35.116638|FR PROD ORGANIC PRODUCE|0.0|4|COO ORG ROMA TOMATOES|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00294087000002|FRESH PRODUCE|PRODUCE|-80.85753|1.4112301235300906|204|1
35.116638|0b876d79f33bda0a3badcc6f046b9ffeea9e8d5f|7.98|2015-01-03 12:58:00|1.4091206135396188|1|20405400000|204|0.6129009553309565|0|47|504|-80.85753|64|35.116638|FRESH BERRIES|0.0|4|RED RASPBERRIES 6 OZ|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00715756100019|FRESH PRODUCE|PRODUCE|-80.85753|1.4112301235300906|204|2
35.116638|e196f5ebd301290971015a9b85e544e4022abdec|5.99|2014-09-28 16:58:00|1.4091206135396188|1|76108880156|204|0.6129009553309565|0|47|1939|-80.85753|465|35.116638|COLD PREP FOODS SIDES|1.0|6|MACARONI & CHEESE FAMILY SIZE|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00761088801568|COLD PREPARED FOODS|DELI|-80.85753|1.4112301235300906|204|1
35.116638|b8e4f6fca9408a9b3cff12874b0bc77a26d50892|15.96|2014-11-16 14:08:00|1.4091206135396188|1|20405400000|204|0.6129009553309565|0|47|504|-80.85753|64|35.116638|FRESH BERRIES|1.99|4|RED RASPBERRIES 6 OZ|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00715756100019|FRESH PRODUCE|PRODUCE|-80.85753|1.4112301235300906|204|4
35.116638|69f4ffe33145aaf47fee16559d6458494e6c39c7|3.99|2014-10-20 17:22:00|80.856688219393845|1|20405400000|204|35.131248911135707|0|15|504|-80.824767|64|35.116751|FRESH BERRIES|2.32|4|RED RASPBERRIES 6 OZ|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00715756100019|FRESH PRODUCE|PRODUCE|-80.85753|80.857532666903609|294|1
35.116638|31f77baa8ebeaacee70d86e09bc8abaddf648365|4.59|2015-03-03 19:56:00|80.856688219393845|1|74236523295|204|35.131248911135707|0|15|1262|-80.824767|57|35.116751|HALF N HALF WHIPPING CREAM|0.6|3|HORIZON ORGANIC HALF&HALF|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00742365232954|MILK|DAIRY|-80.85753|80.857532666903609|294|1
35.116638|4ee813398293f244b893e743132667300c5b5a97|7.98|2014-09-13 19:34:00|1.4091206135396188|1|20405400000|204|0.6129009553309565|0|47|504|-80.85753|64|35.116638|FRESH BERRIES|1.98|4|RED RASPBERRIES 6 OZ|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00715756100019|FRESH PRODUCE|PRODUCE|-80.85753|1.4112301235300906|204|2
35.116638|cc1b2fd5a779bfacd10f62b4bd2863ffbd20ad6d|7.98|2015-01-20 20:09:00|80.856688219393845|1|20405400000|204|35.13124890439326|0|15|504|-80.844274|64|35.204336|FRESH BERRIES|0.0|4|RED RASPBERRIES 6 OZ|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00715756100019|FRESH PRODUCE|PRODUCE|-80.85753|80.857547367555895|61|2
35.116638|74ece516a8aa8b2f7ae8b45c7874a69377f20b65|7.98|2015-02-12 17:17:00|80.856688219393845|1|20405400000|204|35.13124890930947|0|15|504|-80.825175|64|35.152722|FRESH BERRIES|0.0|4|RED RASPBERRIES 6 OZ|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00715756100019|FRESH PRODUCE|PRODUCE|-80.85753|80.857539321200392|160|2
35.116638|ada4e67f16460cab1c5ae66ca4cc5643469193ba|37.98|2014-12-23 19:56:00|80.856688219393845|1|89293100034|204|35.13124890930947|0|15|9964|-80.825175|887|35.152722|NFS-S/PREM-PINOT NOIR|0.0|13|A TO Z PINOT NOIR|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00892931000347|SUPER PREMIUM ($11-$14.99)|WINE|-80.85753|80.857539321200392|160|2
35.116638|36710ca21b33381cd445a68ed69b036d10c316f7|39.98|2014-12-09 21:52:00|1.4091206135396188|1|84849602021|204|0.6129009553309565|0|47|6841|-80.85753|1576|35.116638|SWEAT PANTS/SHIRTS|20.0|18|I/O LADIES CABLE KNIT LEGGINGS|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00848496020214|FAMILY APPAREL|GM|-80.85753|1.4112301235300906|204|2
35.116638|ef9753dd273426eb6fedb5e1e017841085cdb3d6|3.87|2015-01-06 18:33:00|80.856688219393845|1|4800000245|204|35.13124890439326|0|15|190|-80.844274|29|35.204336|TUNA-CANNED|0.8699999999999999|1|COS TUNA CHUNK LIGHT|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00048000002457|SEAFOOD-CANNED|G1 GROCERY|-80.85753|80.857547367555895|61|3
35.116638|efab18d4799396ee9ce0e3a93c8fa9cf0d3f4ecd|4.69|2014-12-14 14:58:00|1.4091206135396188|1|5210000236|204|0.6129009553309565|0|47|1245|-80.85753|34|35.116638|SINGLE SPICES|1.41|1|MC CREAM OF TARTAR|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00052100002361|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.85753|1.4112301235300906|204|1
35.116638|c366617c5742c0ddb26647054fa603883df0c160|4.15|2014-12-31 19:36:00|80.856688219393845|1|4400000488|204|35.131248908216527|0|15|89|-80.85013|12|35.175855|GRAHAM CRACKERS|0.65|1|HONEYMAID GRAHAMS|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00044000004637|COOKIES|G1 GROCERY|-80.85753|80.857541602840982|218|1
35.116638|114f476e827d46753b7886ad7636ff601fe3fcf1|9.99|2015-02-14 16:22:00|80.856688219393845|1|4200044517|204|35.131248911135707|0|15|426|-80.824767|72|35.116751|NFS-PAPER TOWELS|1.0|1|BRAWNY 6 BIG ROLL PICK A SIZE|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00042000445177|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.85753|80.857532666903609|294|1
35.116638|8102150a91a95ac4358406a4b1e52c1c657bf898|14.38|2015-02-06 12:23:00|1.4091206135396188|1|3760035160|204|0.6129009553309565|0|47|845|-80.85753|100|35.116638|NATURAL/ORGANIC BACON|3.59|19|HORMEL NATURAL CHOICE BACON|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00037600445955|BACON|CASE READY MEATS|-80.85753|1.4112301235300906|204|2
35.116638|9b29bf84341f875900993ce6aceb69742e63f460|7.99|2015-01-24 15:04:00|1.4091206135396188|1|3760035160|204|0.6129009553309565|0|47|845|-80.85753|100|35.116638|NATURAL/ORGANIC BACON|0.0|19|HORMEL NATURAL CHOICE BACON|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00037600445955|BACON|CASE READY MEATS|-80.85753|1.4112301235300906|204|1
35.116638|1fc745190a6aaf47ca13c4e0e7350e65243da595|7.19|2015-02-18 11:24:00|80.856688219393845|1|3760035160|204|35.13124890930947|0|15|845|-80.825175|100|35.152722|NATURAL/ORGANIC BACON|0.0|19|HORMEL NATURAL CHOICE BACON|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00037600445955|BACON|CASE READY MEATS|-80.85753|80.857539321200392|160|1
35.116638|fcc4e0298bd57f5549933882a1675756aec5e0a7|3.38|2014-12-20 17:27:00|80.856688219393845|1|7203688003|204|35.131248911135707|0|15|527|-80.824767|64|35.116751|FRESH CARROTS|0.38|4|HT BABY CARROTS 1LB BAG|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00072036880031|FRESH PRODUCE|PRODUCE|-80.85753|80.857532666903609|294|2
35.116638|125f7c2f60a806705037bd12cf254204d7c5f9b4|1.69|2015-01-18 11:41:00|80.856688219393845|1|7203688003|204|35.131248911135707|0|15|527|-80.824767|64|35.116751|FRESH CARROTS|0.0|4|HT BABY CARROTS 1LB BAG|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00072036880031|FRESH PRODUCE|PRODUCE|-80.85753|80.857532666903609|294|1
35.116638|9f69419d4256a6885344211eea8cabe83636cd5f|1.69|2015-01-31 19:42:00|80.856688219393845|1|7203688003|204|35.131248909433786|0|15|527|-80.849471|64|35.161696|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00072036880031|FRESH PRODUCE|PRODUCE|-80.85753|80.857539025206648|35|1
35.116638|565cabcdf02a2e6b894a8e1bd820998438cceb98|3.38|2014-09-12 05:19:00|1.4091206135396188|1|7203688003|204|0.6129009553309565|0|47|527|-80.85753|64|35.116638|FRESH CARROTS|0.38|4|HT BABY CARROTS 1LB BAG|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00072036880031|FRESH PRODUCE|PRODUCE|-80.85753|1.4112301235300906|204|2
35.116638|4359c1ba0026537be192a38fff2f4f5ef157197a|1.69|2015-02-23 16:49:00|80.856688219393845|1|7203688003|204|35.131248909433786|0|15|527|-80.849471|64|35.161696|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00072036880031|FRESH PRODUCE|PRODUCE|-80.85753|80.857539025206648|35|1
35.116638|7df51234882e4b57b75768ac3af171c3d4fa9046|1.69|2014-10-15 18:34:00|80.856688219393845|1|7203688003|204|35.131248909433786|0|15|527|-80.849471|64|35.161696|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00072036880031|FRESH PRODUCE|PRODUCE|-80.85753|80.857539025206648|35|1
35.116638|2d464f5139513abb8c2a86fe03e618585315a5f1|1.69|2014-11-03 17:45:00|80.856688219393845|1|7203688003|204|35.131248909433786|0|15|527|-80.849471|64|35.161696|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00072036880031|FRESH PRODUCE|PRODUCE|-80.85753|80.857539025206648|35|1
35.116638|6771f3c70070bcb80e0cf709896d7d31ab494d5b|3.38|2014-12-08 16:47:00|80.856688219393845|1|7203688003|204|35.131248909433786|0|15|527|-80.849471|64|35.161696|FRESH CARROTS|0.38|4|HT BABY CARROTS 1LB BAG|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00072036880031|FRESH PRODUCE|PRODUCE|-80.85753|80.857539025206648|35|2
35.116638|569092baa3b6f02f08473b7691a5798dddb6e82e|1.69|2014-11-25 06:02:00|1.4091206135396188|1|7203688003|204|0.6129009553309565|0|47|527|-80.85753|64|35.116638|FRESH CARROTS|0.0|4|HT BABY CARROTS 1LB BAG|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00072036880031|FRESH PRODUCE|PRODUCE|-80.85753|1.4112301235300906|204|1
35.116638|e9f8fed6315fd47f51508c97d75ccce132aa3ff1|2.99|2014-11-10 19:12:00|80.856688219393845|1|3338365583|204|35.131248911135707|0|15|522|-80.824767|64|35.116751|FRESH TOMATOES|0.2|4|SWEET GRAPE TOMATO (PINT)|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00072036880284|FRESH PRODUCE|PRODUCE|-80.85753|80.857532666903609|294|1
35.116638|e8f833e91bed11f96ba8c2f3813047917693e9b3|4.49|2015-02-04 15:12:00|80.856688219393845|1|7203695649|204|35.131248911135707|0|15|1699|-80.824767|387|35.116751|EVERYDAY (COOKIES)|1.0|14|HT CHOCO, CHOCO FROSTED COOKIE|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00072036956514|COOKIES|BAKERY|-80.85753|80.857532666903609|294|1
35.116638|bc161559c44d13b236f33bbf3787c45fc6693ff6|4.0|2014-11-25 17:07:00|1.4091206135396188|1|65780295163|204|0.6129009553309565|0|47|1165|-80.85753|87|35.116638|NFS-FRESH CONSUMER BUNCH|0.0|9|BUNCH- ALSTROEMERIA   RIVERD|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00657802951636|FLORAL|FLORAL|-80.85753|1.4112301235300906|204|1
35.116638|fd4e8a0187ddd90060ebab045e346c8447e3e3cb|5.69|2014-09-23 12:44:00|80.856688219393845|1||204|35.131248911135707|0|15|523|-80.824767|64|35.116751|FRESH POTATOES|1.32|4|COO SWEET POTATOES, BULK|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00204091000004|FRESH PRODUCE|PRODUCE|-80.85753|80.857532666903609|294|1
35.116638|ef792291bdb145c738eea3e80000aef473b84083|3.04|2015-02-10 19:44:00|80.856688219393845|1||204|35.131248908216527|0|15|523|-80.85013|64|35.175855|FRESH POTATOES|0.31|4|COO SWEET POTATOES, BULK|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00204091000004|FRESH PRODUCE|PRODUCE|-80.85753|80.857541602840982|218|1
35.116638|a3de805ea055021d2113501b2f0b2b693536fa17|3.32|2014-11-04 13:10:00|1.4091206135396188|1||204|0.6129009553309565|0|47|523|-80.85753|64|35.116638|FRESH POTATOES|0.78|4|COO SWEET POTATOES, BULK|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00204091000004|FRESH PRODUCE|PRODUCE|-80.85753|1.4112301235300906|204|1
35.116638|3730bd830c6b971147dc2aaa8fe3dcdb0f0db683|21.98|2015-02-21 20:44:00|80.856688219393845|1|7017787949|204|35.13124890439326|0|15|1247|-80.844274|37|35.204336|SINGLES PODS CUPS TEA|6.0|1|TWININGS TEA KCUP CHAI LATTE|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00070177879495|TEA|G1 GROCERY|-80.85753|80.857547367555895|61|2
35.116638|851350b7541cac8df0e521181cd5cc0a06b1f38b|1.69|2014-12-26 08:25:00|80.856688219393845|1|4900000044|204|35.131248908216527|0|15|55|-80.85013|8|35.175855|REGULAR|0.0|23|CB COKE SINGLE 20 OZ.|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00049000000443|CARBONATED BEVERAGES|BEVERAGE|-80.85753|80.857541602840982|218|1
35.116638|a4128669bcd80d19012adf23d2f89723b2bedfed|1.69|2015-02-17 14:39:00|80.856688219393845|1|4900000044|204|35.13124890930947|0|15|55|-80.825175|8|35.152722|REGULAR|0.0|23|CB COKE SINGLE 20 OZ.|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00049000000443|CARBONATED BEVERAGES|BEVERAGE|-80.85753|80.857539321200392|160|1
35.116638|912f41ced1cccba6543c29269582c5d1b68545ea|2.4|2015-02-15 17:21:00|80.856688219393845|1|7047000100|204|35.131248911135707|0|15|687|-80.824767|61|35.116751|BLENDED|0.0|3|YOPLAIT RASPBERRY YOGURT|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00070470003016|YOGURT|DAIRY|-80.85753|80.857532666903609|294|4
35.116638|c01cf69c4ce8a70d6b72349eab52267bfa0d094b|1.67|2014-12-14 11:32:00|80.856688219393845|1|7046208251|204|35.131248908216527|0|15|53|-80.85013|7|35.175855|THEATER BOX|0.33|1|SOUR PATCH KIDS THEATER BOX|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00070462098358|CANDY|G1 GROCERY|-80.85753|80.857541602840982|218|1
35.116638|66187281dac7fb9e23a155c7258f3958c73eb546|3.49|2014-11-24 07:40:00|80.856688219393845|1|7146426040|204|35.131248908216527|0|15|577|-80.85013|136|35.175855|OTHER MERCH FR MSC JUICE|0.0|4|BOLTHOUSE PERF PROTEN VAN CHAI|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00071464260408|OTHER MERCHANDISE|PRODUCE|-80.85753|80.857541602840982|218|1
35.116638|99cae10685b9f79f04c8c0932ccf597360513a8b|4.99|2014-12-23 11:40:00|80.856688219393845|1|7146426060|204|35.131248908216527|0|15|577|-80.85013|136|35.175855|OTHER MERCH FR MSC JUICE|0.0|4|BOLTHOUSE BERRY BOOST|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00071464280604|OTHER MERCHANDISE|PRODUCE|-80.85753|80.857541602840982|218|1
35.116638|42535eabff199a36f765e17630ffe835bbc18760|4.99|2015-02-04 05:13:00|1.4091206135396188|1|7146426060|204|0.6129009553309565|0|47|577|-80.85753|136|35.116638|OTHER MERCH FR MSC JUICE|0.0|4|BOLTHOUSE PERFECTLY PROTEIN|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00071464260606|OTHER MERCHANDISE|PRODUCE|-80.85753|1.4112301235300906|204|1
35.116638|479631df2d0f0bbee9702ca7f0f5a8bd06be3047|7.29|2014-11-14 11:41:00|80.856688219393845|1|5210000234|204|35.13124890930947|0|15|1245|-80.825175|34|35.152722|SINGLE SPICES|2.19|1|MC WHOLE CLOVES|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00052100002347|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.85753|80.857539321200392|160|1
35.116638|3ac0f41baed60df6e9ea415a140b482af0db6a02|8.99|2014-11-26 20:10:00|80.856688219393845|1|4900003165|204|35.131248908216527|0|15|31|-80.85013|4|35.175855|NON CARBONATED WATER|4.5|1|DASANI .5 LITER 24 PK|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00049000031652|BOTTLED WATER|G1 GROCERY|-80.85753|80.857541602840982|218|1
35.116638|2e92c00bb016fe1d94aa554faf38f0df185f7a1e|2.39|2014-10-28 20:36:00|1.4091206135396188|1|5150055538|204|0.6129009553309565|0|47|8|-80.85753|2|35.116638|BROWNIE MIXES|1.2|1|PILLS MILK CHOCOLATE BROWNIE|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00051500555392|BAKING MIXES|G1 GROCERY|-80.85753|1.4112301235300906|204|1
35.116638|f468c0edd61461f479cec10737bc20bf8785acfa|7.98|2014-11-15 10:08:00|80.856688219393845|1|7203663995|204|35.131248911135707|0|15|342|-80.824767|57|35.116751|FRESH MILK|0.0|3|HARRIS TEETER 1% MILK|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00072036631275|MILK|DAIRY|-80.85753|80.857532666903609|294|2
35.116638|1656d0a172146a4078fa1b1d17406281adf90925|3.99|2014-09-14 20:54:00|80.856688219393845|1|3338300084|204|35.13124890930947|0|15|500|-80.825175|64|35.152722|FRESH APPLES|0.0|4|GOLD DEL APPLE 3LB BAG|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00072036880277|FRESH PRODUCE|PRODUCE|-80.85753|80.857539321200392|160|1
35.116638|477dfbd278bf639474d180b9ba21c180d7d63b07|3.79|2015-03-08 09:57:00|80.856688219393845|1|7203688014|204|35.13124890930947|0|15|581|-80.825175|136|35.152722|FRESH SALSA|0.0|4|HT FRESH MEDIUM SALSA|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00072036880222|OTHER MERCHANDISE|PRODUCE|-80.85753|80.857539321200392|160|1
35.116638|f47d02004557c8a2d002bee21a278f493616783c|8.07|2015-01-10 14:55:00|80.856688219393845|1|1800000401|204|35.131248908216527|0|15|327|-80.85013|54|35.175855|DINNER ROLLS-REFRIGERATED|0.0|3|PILLSBURY CRESCENT ROLLS|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00018000004010|DOUGH PRODUCTS|DAIRY|-80.85753|80.857541602840982|218|3
35.116638|4c3e9b3a43efe3cfcdd3d2f3ece1c78d72a02ed1|8.58|2015-01-10 10:37:00|80.856688219393845|1|2840015636|204|35.131248911135707|0|15|204|-80.824767|31|35.116751|TORTILLA CHIPS|2.15|1|DORTIOS NACHO CHEESE|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00028400156363|SNACKS|G1 GROCERY|-80.85753|80.857532666903609|294|2
35.116638|a90e6c850e291848707c1fb691906fce4274fbdc|3.69|2014-12-21 17:13:00|80.856688219393845|1|88491201424|204|35.131248911135707|0|15|74|-80.824767|9|35.116751|RTE CEREAL ALL FAMILY|0.0|1|POST HNY BUNCHES HONEY RSTD|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00884912014245|CEREAL|G1 GROCERY|-80.85753|80.857532666903609|294|1
35.116638|2fadcfbf1fb1babdceca7f4057e7fcfeb1d88e8b|3.19|2015-03-09 14:42:00|80.856688219393845|1|82951530146|204|35.131248911135707|0|15|205|-80.824767|31|35.116751|REMAINING SNACKS|0.0|1|SENSBL PORT VEG STRAW RS OLV O|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00829515302108|SNACKS|G1 GROCERY|-80.85753|80.857532666903609|294|1
35.116638|5656bc6461f2e6c70da25233a2618e1a1e7b3fd4|8.98|2014-12-21 17:55:00|1.4091206135396188|1|4078498500|204|0.6129009553309565|0|47|257|-80.85753|39|35.116638|TOMATOES|0.0|1|SAN MARZANO TOM DICED|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00040784987500|VEGETABLES-CAN/JAR|G1 GROCERY|-80.85753|1.4112301235300906|204|2
35.116638|eceb901290f5799c986f4dce8e30472a13a1f8e7|5.99|2015-02-25 15:52:00|1.4091206135396188|1|4667741050|204|0.6129009553309565|0|47|6142|-80.85753|1546|35.116638|BULB-COMPACT FLUORESCENTS|0.0|18|PHILIP ECOVANTAGE 29W CLEAR|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00046677410506|LIGHT BULBS/ELECTRICAL|GM|-80.85753|1.4112301235300906|204|1
35.116638|ea22b69532ae84dc14898af6c739d5a6b538b920|2.99|2014-11-22 17:00:00|80.856688219393845|1|4113700642|204|35.13124890930947|0|15|386|-80.825175|65|35.152722|NFS-FIREPLACE LOGS|0.49|1|DURAFLAME STIX FIRELIGHTERS|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00041137006428|CHARCOAL/LOGS/ACCESSORIES|G1 GROCERY|-80.85753|80.857539321200392|160|1
35.116638|db3e445d3a8dd310367dbf9519b6e2ecb568f14c|7.99|2014-12-12 15:47:00|1.4091206135396188|1|5170081049|204|0.6129009553309565|0|47|388|-80.85753|66|35.116638|NFS-DISHWASH PWDR/LIQUID|0.0|1|FINISH POWERBALL FRESH 32CT|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00051700810499|DETERGENTS|G1 GROCERY|-80.85753|1.4112301235300906|204|1
35.116638|88c3a1a5aa4a1bd97fde5c2e773e7ce6a278c7c0|0.56|2015-03-08 17:49:00|80.856688219393845|1||204|35.131248909433786|0|15|524|-80.849471|64|35.161696|FRESH PROD FRESH ONIONS|0.0|4|COO SHALLOTS, BULK|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00204662000006|FRESH PRODUCE|PRODUCE|-80.85753|80.857539025206648|35|1
35.116638|4eb76ca2fd3a3234a5bd64422405e59c9da0b8f4|5.94|2014-10-04 11:35:00|80.856688219393845|1||204|35.13124890930947|0|15|562|-80.825175|64|35.152722|FRESH CUT FRUIT|0.0|4|SLICED STRAWBERRIES BY/LB|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00204217000000|FRESH PRODUCE|PRODUCE|-80.85753|80.857539321200392|160|1
35.116638|91833752ea6cd83935f06b54dee97f46edc09dba|3.99|2014-12-19 18:43:00|80.856688219393845|1|3338324028|204|35.131248911135707|0|15|504|-80.824767|64|35.116751|FRESH BERRIES|2.32|4|BLACKBERRIES 5.6 OZ|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00761635202602|FRESH PRODUCE|PRODUCE|-80.85753|80.857532666903609|294|1
35.116638|2286180b959406dadfbcbf0f589ce57c6ddadbe4|3.99|2014-11-03 08:44:00|80.856688219393845|1|75166677005|204|35.131248911135707|0|15|522|-80.824767|64|35.116751|FRESH TOMATOES|0.0|4|NATURESWEET CHERUBS 10.5 OZ|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00751666770058|FRESH PRODUCE|PRODUCE|-80.85753|80.857532666903609|294|1
35.116638|137012f289d9dfa30dd75c37c64cc8855d64d765|10.98|2014-12-06 09:34:00|80.856688219393845|1|827411111|204|35.131248911135707|0|15|55|-80.824767|8|35.116751|REGULAR|3.0|23|REEDS EXTRA GINGER BREW|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00008274444445|CARBONATED BEVERAGES|BEVERAGE|-80.85753|80.857532666903609|294|2
35.116638|9449365c004267242ac9e68750a55644a1d959f3|7.38|2014-12-13 14:46:00|1.4091206135396188|1|1410007412|204|0.6129009553309565|0|47|1253|-80.85753|12|35.116638|ALL OTHER COOKIES|1.0|1|PF MILANO MILK CHOCOLATE|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00014100099970|COOKIES|G1 GROCERY|-80.85753|1.4112301235300906|204|2
35.116638|1d0337de2beb6472c1b083351e8ba9d6b28ae815|3.39|2014-09-27 18:26:00|80.856688219393845|1|5000000929|204|35.131248911135707|0|15|326|-80.824767|54|35.116751|COOKIES/BROWNIES-REFRIGERATED|0.39|3|I/O NES HALLOWEEN CHOC CHIP|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00050000009299|DOUGH PRODUCTS|DAIRY|-80.85753|80.857532666903609|294|1
35.116638|f6544beb13a7afb45642dd24f5f1b4123b4413c6|3.49|2014-10-09 06:46:00|1.4091206135396188|1|7797508005|204|0.6129009553309565|0|47|202|-80.85753|31|35.116638|PRETZELS|0.3|1|SOH SNAP PRETZEL|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00077975080078|SNACKS|G1 GROCERY|-80.85753|1.4112301235300906|204|1
35.116638|0f23418a8ef8ec4d512fe7c32e26a8d5dcfe6c0e|4.49|2015-01-07 13:33:00|1.4091206135396188|1|2301290007|204|0.6129009553309565|0|47|1483|-80.85753|485|35.116638|SUSHI ROLL AND WRAP|0.0|6|SUMMER ROLL|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00023012900076|SUSHI|DELI|-80.85753|1.4112301235300906|204|1
35.116638|ec7e258ebf7a42dce16384ad1b0de7a351388f7c|2.99|2014-11-21 15:20:00|1.4091206135396188|1|2560000786|204|0.6129009553309565|0|47|1045|-80.85753|173|35.116638|DONUTS|0.99|7|TSTYKAKE SUGAR BAG DNTS|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00025600007860|SWEET BAKED GOODS|COMMERCIAL BAKERY|-80.85753|1.4112301235300906|204|1
35.116638|fa94c46bde22079c396732c6c456fee835f6615d|2.99|2014-10-12 12:32:00|80.856688219393845|1|2560000786|204|35.131248908216527|0|15|1045|-80.85013|173|35.175855|DONUTS|0.99|7|TSTYKAKE SUGAR BAG DNTS|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00025600007860|SWEET BAKED GOODS|COMMERCIAL BAKERY|-80.85753|80.857541602840982|218|1
35.116638|02c0ca24cb04cec5aaf800d6e12ef84ff8677153|2.19|2014-10-17 17:20:00|80.856688219393845|1|4900005010|204|35.131248909433786|0|15|55|-80.849471|8|35.161696|REGULAR|0.2|23|SPRITE  2 LITER|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00049000050158|CARBONATED BEVERAGES|BEVERAGE|-80.85753|80.857539025206648|35|1
35.116638|ce4372f7aff65200295b3959565219badb89bd3f|9.99|2014-09-11 20:42:00|80.856688219393845|1|2301200017|204|35.13124890930947|0|15|1479|-80.825175|485|35.152722|SUSHI HYBRID SPECIALTY|0.0|6|SUSHI ULTIMATE|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00023012000172|SUSHI|DELI|-80.85753|80.857539321200392|160|1
35.116638|6d8368cc74d6f0994e69745f1cba655350972a1d|2.0|2015-01-18 16:31:00|1.4091206135396188|1|7203606031|204|0.6129009553309565|0|47|1146|-80.85753|229|35.116638|SYRUPS|0.0|1|HT CHOCOLATE FLAVOR SYRUP|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00072036060310|COCOAS CREAMERS SYRUPS|G1 GROCERY|-80.85753|1.4112301235300906|204|1
35.116638|d0716af4830cffbf88990707d245d9c85382546c|3.39|2015-01-02 16:56:00|1.4091206135396188|1|5000012734|204|0.6129009553309565|0|47|341|-80.85753|57|35.116638|CREAMERS|0.0|3|COFFEEMATE SF FRENCH VANILLA|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00050000848119|MILK|DAIRY|-80.85753|1.4112301235300906|204|1
35.116638|f16d21229cac60733b4a71615bbf67a4766a08e8|4.19|2015-01-15 08:41:00|80.856688219393845|1|5210007086|204|35.131248905565805|0|15|217|-80.80146|34|35.17739|EXTRACTS FOOD COLORING|0.0|1|E  MCCORMICK VANILLA EXTRACT|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00052100070865|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.85753|80.857545824451464|208|1
35.116638|a60f69703dc04e909f4df41f0d5191ae74e17e9e|2.99|2015-01-12 16:47:00|80.856688219393845|1|7203663104|204|35.131248909433786|0|15|364|-80.849471|55|35.161696|ORGANIC AND CF EGGS|0.0|3|HTN NEST GRADE A LARGE EGG BRO|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00072036631046|EGGS FRESH|DAIRY|-80.85753|80.857539025206648|35|1
35.116638|6eb35b14149434ad27796e260ba7f215161234d2|6.19|2014-10-03 19:42:00|80.856688219393845|1|2800021560|204|35.13124890439326|0|15|16|-80.844274|3|35.204336|BAKING CHOCOLATE/CHIPS/MORSELS|0.0|1|NESTLE SEMISWEET MORSELS|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00028000215606|BAKING SUPPLIES|G1 GROCERY|-80.85753|80.857547367555895|61|1
35.116638|8242d85b7477ecad04e3f5ebdd3407653e4b1b73|1.67|2014-11-11 14:21:00|1.4091206135396188|1|3120001605|204|0.6129009553309565|0|47|106|-80.85753|16|35.116638|CRANBERRY SAUCE|0.17|1|OS CRANBERRY SC WHOLE|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00031200016034|FRUIT-CAN/JAR|G1 GROCERY|-80.85753|1.4112301235300906|204|1
35.116638|2ff15ac6b77a90da159d28ced6efc58d7cd582d8|5.29|2014-10-06 16:27:00|80.856688219393845|1|7590000534|204|35.131248909433786|0|15|494|-80.849471|107|35.161696|HEAT & EAT SIDES|0.0|19|BOB EVANS FAMILY MASHED POTATO|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00075900005349|HEAT & EAT|CASE READY MEATS|-80.85753|80.857539025206648|35|1
35.116638|fd1523de91d15c356fe0a3ff7d518212a98bf6b6|5.69|2014-09-22 20:34:00|80.856688219393845|1|7756725423|204|35.131248911135707|0|15|252|-80.824767|45|35.116751|PREMIUM ICE CREAM|2.84|5|BREYERS CHOCOLATE I/C|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00077567254207|ICE CREAM|FROZEN|-80.85753|80.857532666903609|294|1
35.116638|f38de08de8f37761f61d988625ff5ca4a76d08b8|7.69|2014-10-23 14:13:00|1.4091206135396188|1|8087800550|204|0.6129009553309565|0|47|3503|-80.85753|1045|35.116638|CONDITIONER-PREMIUM|0.0|17|PANTENE CND DLY MOIS RENEWAL|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00080878171316|HAIR & SCALP CARE|HBC|-80.85753|1.4112301235300906|204|1
35.116638|3f18ffd190d4229b986776acf6635ff76c67953a|5.29|2015-02-10 17:59:00|80.856688219393845|1|7590000534|204|35.131248911135707|0|15|494|-80.824767|107|35.116751|HEAT & EAT SIDES|0.0|19|BOB EVANS FAMILY MASHED POTATO|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00075900005349|HEAT & EAT|CASE READY MEATS|-80.85753|80.857532666903609|294|1
35.116638|9845c3c909fbde32c58b671ed513c17f8ac483f3|3.99|2015-02-02 13:02:00|80.856688219393845|1|66559609901|204|35.131248908216527|0|15|326|-80.85013|54|35.175855|COOKIES/BROWNIES-REFRIGERATED|0.0|3|IMMACULATE BAKE CHOC CHUNK|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00665596099014|DOUGH PRODUCTS|DAIRY|-80.85753|80.857541602840982|218|1
35.116638|4ba6c1747bfe769c03a5cf4aea16fd365adda406|1.29|2015-01-28 15:15:00|1.4091206135396188|1|1657191030|204|0.6129009553309565|0|47|30|-80.85753|4|35.116638|CARBONATED WATER|0.29|1|SPARKLING ICE STRWBRY LEMONADE|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00016571950293|BOTTLED WATER|G1 GROCERY|-80.85753|1.4112301235300906|204|1
35.116638|235a3bc5d99fbcc26f888d52360446c23d2610db|6.79|2014-11-05 06:00:00|1.4091206135396188|1|4850001833|204|0.6129009553309565|0|47|335|-80.85753|56|35.116638|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA CALCIUM ORANGE JUICE|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00048500018309|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.85753|1.4112301235300906|204|1
35.116638|11f914a74076d4ace25baf3788346769eb0584f5|3.98|2014-11-13 17:34:00|1.4091206135396188|1|7203698370|204|0.6129009553309565|0|47|205|-80.85753|31|35.116638|REMAINING SNACKS|0.98|1|HT SNACK MIX CHEDDAR|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00072036983718|SNACKS|G1 GROCERY|-80.85753|1.4112301235300906|204|2
35.116638|c22c748ec7edfb7c79af7199ccabd9fe38eb117b|3.98|2014-11-13 15:48:00|1.4091206135396188|1|7203698370|204|0.6129009553309565|0|47|205|-80.85753|31|35.116638|REMAINING SNACKS|0.98|1|HT SNACK MIX CHEDDAR|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00072036983718|SNACKS|G1 GROCERY|-80.85753|1.4112301235300906|204|2
35.116638|9d51ff099b1cd2ea5424d3fe4d68c469b3ed9a49|4.98|2014-09-12 05:11:00|1.4091206135396188|1|7978412711|204|0.6129009553309565|0|47|6618|-80.85753|1564|35.116638|FILLER PAPER|0.0|18|COLLEGE RULE FILLER PAPER 150C|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00079784127111|SCHOOL & OFFICE SUPPLY|GM|-80.85753|1.4112301235300906|204|2
35.116638|be97842bbf0aaebf2b4ab51cd1115394aafd970f|2.49|2015-02-11 16:56:00|80.856688219393845|1|7316826748|204|35.131248911135707|0|15|6975|-80.824767|1600|35.116751|VALENTINE CARDS IMP|0.49|18|AVENGER ASSEMBLE VAL CARDS|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00073168267486|SEASONAL MERCHANDISE|GM|-80.85753|80.857532666903609|294|1
35.116638|6bde9a252de633016c07ac762f9b50947f9855c9|5.97|2014-10-09 20:51:00|1.4091206135396188|1|7203676359|204|0.6129009553309565|0|47|345|-80.85753|57|35.116638|ORGANIC MILK|0.0|3|HTO ORGANIC FF SKIM GAL|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00072036763624|MILK|DAIRY|-80.85753|1.4112301235300906|204|1
35.116638|b93dcd4f1a9595122a38ec3fe8a12ff2e3d5bcc3|13.16|2015-03-02 17:53:00|80.856688219393845|1|7203688004|204|35.131248911135707|0|15|527|-80.824767|64|35.116751|FRESH CARROTS|0.0|4|HT BABY CARROTS 2LB BAG|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00072036880048|FRESH PRODUCE|PRODUCE|-80.85753|80.857532666903609|294|4
35.116638|7d5f8b9355fa83b2e3d74ab036af0264e2f4e770|9.53|2014-11-01 18:45:00|80.856688219393845|1|20617400000|204|35.131248908216527|0|15|1832|-80.85013|415|35.175855|BH SLICING CHEESE|0.0|6|BOARS HEAD MANCHEGO CHEESE|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00206174000000|SLICING CHEESE|DELI|-80.85753|80.857541602840982|218|1
35.116638|142ec409108a35cd8f1593c2c84b2c2500b90459|18.99|2014-11-24 05:59:00|1.4091206135396188|1|4740030374|204|0.6129009553309565|0|47|3917|-80.85753|1075|35.116638|DISPOSABLE RAZOE-MEN|0.0|17|MACH3 DISPOSABLE RAZORS SENS|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00047400303744|SHAVING NEEDS/MEN HAIR|HBC|-80.85753|1.4112301235300906|204|1
35.116638|b2db05f635e1be3583976f58a4ffda736b64a0c0|0.6|2015-03-06 10:21:00|80.856688219393845|1|7047000100|204|35.131248905565805|0|15|687|-80.80146|61|35.17739|BLENDED|0.0|3|YOPLAIT ORG MIXED BERRY|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00070470003108|YOGURT|DAIRY|-80.85753|80.857545824451464|208|1
35.116638|2e89e3c72c0e96ee708edcd7a4ea6e8ed7c34071|3.39|2015-01-14 13:22:00|1.4091206135396188|1|5260305445|204|0.6129009553309565|0|47|214|-80.85753|33|35.116638|BROTH|0.0|1|PACIFIC ORG LS BEEF BROTH|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00052603054362|SOUP|G1 GROCERY|-80.85753|1.4112301235300906|204|1
35.116638|8d5f62327ca6de94a289ccf8b101840e3b203ad6|2.99|2014-10-31 17:01:00|80.856688219393845|1|2500005426|204|35.131248908216527|0|15|338|-80.85013|56|35.175855|OTHER FRUIT JUICES|0.99|3|SIMPLY LEMONADE|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00025000054266|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.85753|80.857541602840982|218|1
35.116638|eb55832da6a0d6aacd2bc3e01ee122f282aa34a7|7.99|2014-11-15 17:14:00|80.856688219393845|1|8834510005|204|35.131248909433786|0|15|459|-80.849471|83|35.161696|IMPORT BEER|0.0|16|NEWCASTLE BROWN 6PK 12OZ BTL|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00088345100050|IMPORT BEER|BEER|-80.85753|80.857539025206648|35|1
35.116638|48c8f3ca78fa4bba34a2ec6e1e461df388d2a6f8|3.99|2015-02-09 19:50:00|1.4091206135396188|1|9396600033|204|0.6129009553309565|0|47|1262|-80.85753|57|35.116638|HALF N HALF WHIPPING CREAM|0.0|3|ORGANIC VALLEY HALF & HALF|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00093966000337|MILK|DAIRY|-80.85753|1.4112301235300906|204|1
35.116638|831370329dd0449fcfc75ad825c5528a4fe6578b|3.49|2014-12-09 21:12:00|80.856688219393845|1|4319415976|204|35.131248911135707|0|15|3698|-80.824767|1060|35.116751|PONYTAIL HOLDER|1.0|17|SCUNCI 18PK L ND ELASTICS BRWN|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00043194167760|HAIR CARE ACCESSORIES|HBC|-80.85753|80.857532666903609|294|1
35.116638|d853a1ced631810449411ebfcac387e78211c835|11.98|2014-12-14 13:17:00|1.4091206135396188|1|2301200009|204|0.6129009553309565|0|47|1479|-80.85753|485|35.116638|SUSHI HYBRID SPECIALTY|0.0|6|WRAP DELIGHT|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00023012000097|SUSHI|DELI|-80.85753|1.4112301235300906|204|2
35.116638|58294929dd8cf374ac0444628ffe670f586d875a|17.98|2014-12-05 07:09:00|80.856688219393845|1|4460000228|204|35.131248911135707|0|15|724|-80.824767|69|35.116751|NFS-DRAIN CLEANER/OPENER|0.0|1|LIQUID PLUMR PROF STRENGTH|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00044600002286|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.85753|80.857532666903609|294|2
35.116638|c2a9f895ece97e49b5e07c9dc39975d3443bc1f1|8.99|2014-10-19 17:26:00|1.4091206135396188|1|4460000228|204|0.6129009553309565|0|47|724|-80.85753|69|35.116638|NFS-DRAIN CLEANER/OPENER|0.0|1|LIQUID PLUMR PROF STRENGTH|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00044600002286|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.85753|1.4112301235300906|204|1
35.116638|7295b22dd1133d1bbfe32faf7a3b811675dbaa94|5.79|2015-01-27 14:32:00|1.4091206135396188|1|7247000603|204|0.6129009553309565|0|47|1641|-80.85753|377|35.116638|PACKAGED DONUTS|0.0|14|K K 12 CT GLAZED DONUTS PP|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00072470006035|DONUTS|BAKERY|-80.85753|1.4112301235300906|204|1
35.116638|3bd2e7c50c0231fd680889bef0d76378ddda7a69|1.49|2015-02-26 18:39:00|80.856688219393845|1|2200001340|204|35.131248908216527|0|15|727|-80.85013|7|35.175855|SEASONAL CANDY-SINGLE FAC|0.75|1|I/O(E15)STARBRST ORG JLYBN SS|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00022000013408|CANDY|G1 GROCERY|-80.85753|80.857541602840982|218|1
35.116638|81da181500f0b48c568bd2aaed64dce1ef7887ce|4.69|2014-10-01 18:01:00|80.856688219393845|1|5100007620|204|35.13124890439326|0|15|264|-80.844274|307|35.204336|DESSERT CAKES FROZEN|0.0|5|PEP FARM COCONUT CAKE|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00051000076250|DESSERTS FROZEN|FROZEN|-80.85753|80.857547367555895|61|1
35.116638|8cb98097ca7e13daa4f0d058f429bf29553a447f|5.99|2014-11-19 18:51:00|80.856688219393845|1|20531100000|204|35.131248908216527|0|15|1935|-80.85013|465|35.175855|CHEF CASE|0.0|6|GRILLED FARM RAISED SALMON|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00205311000002|COLD PREPARED FOODS|DELI|-80.85753|80.857541602840982|218|1
35.116638|7b55c27eb507dad32629e615b5cece3b3fdd3789|4.0|2015-01-22 19:31:00|80.856688219393845|1|7203663118|204|35.131248910102755|0|15|1262|-80.816172|57|35.059823|HALF N HALF WHIPPING CREAM|0.0|3|HT HALF & HALF|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00072036632043|MILK|DAIRY|-80.85753|80.857537227236833|66|2
35.116638|897ac76a69ebece4490f8514749112741653c27a|7.99|2015-02-05 17:47:00|80.856688219393845|1|7203695310|204|35.131248911135707|0|15|1970|-80.824767|475|35.116751|COLD PRE-MADE|0.0|6|FIVE CHEESE PIZZA|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00072036953100|PIZZA|DELI|-80.85753|80.857532666903609|294|1
35.116638|9a747f6d4edcafdc559770cc622edff8a616b27a|9.99|2014-10-14 10:56:00|80.856688219393845|1|7203696996|204|35.13124890439326|0|15|751|-80.844274|87|35.204336|NFS-BOUQUETS|0.0|9|9.99 DUOCHROMATIC BQT  SS|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00072036969965|FLORAL|FLORAL|-80.85753|80.857547367555895|61|1
35.116638|c3db3f1e0890934d663ab62fdc8a1573907eac67|3.99|2015-02-14 08:13:00|80.856688219393845|1|4400002854|204|35.131248908216527|0|15|90|-80.85013|13|35.175855|SNACK CRACKERS|0.49|1|OREO RED VELVET LIMITED EDITN|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00044000039455|CRACKERS|G1 GROCERY|-80.85753|80.857541602840982|218|1
35.116638|84f6014f676feb3443a5b0c69bc6c35862f6bb36|17.99|2014-09-26 19:23:00|1.4091206135396188|1|75452700417|204|0.6129009553309565|0|47|458|-80.85753|82|35.116638|CRAFT BEER|0.0|16|NEW BELGIUM SHIFT 12PK CANS|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00754527004170|DOMESTIC BEER|BEER|-80.85753|1.4112301235300906|204|1
35.116638|7ef3c56dc32e01654c141b4c41578e070256becb|38.99|2014-12-18 13:33:00|80.856688219393845|1|8847398050|204|35.13124890930947|0|15|9976|-80.825175|888|35.152722|NFS-U/PREM-PINOT NOIR|0.0|13|SOKOL BLOSSER PINOT NOIR|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00088473980500|ULTRA PREMIUM ($15-$19.99)|WINE|-80.85753|80.857539321200392|160|1
35.116638|5fd113cd054241c6fc52f5a4f52b503ae128c3b9|6.79|2014-09-16 20:22:00|80.856688219393845|1|7064003404|204|35.131248908216527|0|15|252|-80.85013|45|35.175855|PREMIUM ICE CREAM|3.4|5|B BUNNY CHUNKY COOKIE DOUGH|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00070640034222|ICE CREAM|FROZEN|-80.85753|80.857541602840982|218|1
35.116638|3ce974148eb99e1f72d1074122d8ec643f7d0753|2.29|2014-10-21 16:26:00|80.856688219393845|1|7203609021|204|35.131248909433786|0|15|88|-80.849471|13|35.161696|FLAKED SODA CRACKERS|0.4|1|HARRIS TEETER SALTINES|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00072036090218|CRACKERS|G1 GROCERY|-80.85753|80.857539025206648|35|1
35.116638|e29ff5bfe01e2bb399359ef14036c63c6f2860ac|10.89|2014-10-02 21:50:00|1.4091206135396188|1|7119000601|204|0.6129009553309565|0|47|156|-80.85753|24|35.116638|NFS-DOG FOOD-DRY|0.0|1|RACH RAY NUTRSH BEEF&RCE DOGFD|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00071190006035|PET FOOD/SUPPLIES|G1 GROCERY|-80.85753|1.4112301235300906|204|1
35.116638|168a507c20752db2a10ed058e7e3d4d59f95b81d|4.39|2014-09-19 16:46:00|1.4091206135396188|1|6843738350|204|0.6129009553309565|0|47|46|-80.85753|7|35.116638|PKG CHOC|0.89|1|BROOKSDE POMEGRANATE|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|0.61242566243833529|00068437389082|CANDY|G1 GROCERY|-80.85753|1.4112301235300906|204|1
35.116638|53e6170cbb92c2b139c001dc3192b4ff78fa97a9|11.59|2014-11-06 11:45:00|80.856688219393845|1|30573016940|204|35.131248908216527|0|15|4317|-80.85013|1205|35.175855|IBUPROFEN|0.0|17|ADVIL LIQUI-GELS  -16940|49ab44a582fd49d1636fae85f3ec615080ba1694|1.0095786866403311|35.134355925261694|00305730169400|PAIN RELIEF|HBC|-80.85753|80.857541602840982|218|1
35.17739|75c61352a352d28fdf41b83b8f5fc9185df6ffb0|3.69|2014-09-29 13:11:00|80.801203185414451|2|5000012734|208|35.188908061373944|0|24|341|-80.826724|57|35.195689|CREAMERS|1.19|3|COFFEEMATE SF ITALIAN SWT CRM|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|35.194272495053255|00050000145782|MILK|DAIRY|-80.80146|80.801461070058423|412|1
35.17739|24d47fa581eb199d2dc34348508e742a2fdad2d0|4.49|2015-03-04 17:22:00|1.4094857484078087|2|4812127707|208|0.613961277758128|0|26|1036|-80.80146|164|35.17739|BREAKFAST BAGELS|2.25|7|THOMAS HNYWHEAT BGL 6CT PP|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|0.61471665291522548|00048121226152|BREAKFAST|COMMERCIAL BAKERY|-80.80146|1.4102515174184975|208|1
35.17739|ca17c06794eb35b9b0172898bd4face7f32837cd|4.75|2014-11-09 13:29:00|1.4094857484078087|2|4610000715|208|0.613961277758128|0|26|332|-80.80146|52|35.17739|STRING/SNACK|0.0|3|SARGENTO STRING CHS CALCIUM|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|0.61471665291522548|00046100007150|CHEESE|DAIRY|-80.80146|1.4102515174184975|208|1
35.17739|2d89b76ff661ff87f7c4a373fd79ec1c56b8a382|4.79|2014-10-13 11:49:00|1.4094857484078087|2|4610000715|208|0.613961277758128|0|26|332|-80.80146|52|35.17739|STRING/SNACK|0.8|3|SARGENTO STRING CHS CALCIUM|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|0.61471665291522548|00046100007150|CHEESE|DAIRY|-80.80146|1.4102515174184975|208|1
35.17739|a0aeb61a5809f6b29f07297489c36b332f7ae52b|2.65|2015-02-01 16:44:00|1.4094857484078087|2|4119640471|208|0.613961277758128|0|26|1201|-80.80146|33|35.17739|RTS CANNED|0.65|1|PROG LIGHT NE CLAM CHOWDER|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|0.61471665291522548|00041196452815|SOUP|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|b2aa1cc985526dcd2fb5a6d8e5dcc6fcf8d5a15d|8.85|2014-10-22 12:18:00|1.4094857484078087|2|2370002188|208|0.613961277758128|0|26|291|-80.80146|48|35.17739|FROZEN POUTLRY|0.0|5|TYSON PULLED CHICK BREAST|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|0.61471665291522548|00023700039644|FROZEN MEALS|FROZEN|-80.80146|1.4102515174184975|208|1
35.17739|84e4d9f9681a93eebbcf0feae7a5df890a10efd3|4.99|2014-12-14 12:20:00|1.4094857484078087|2|2410044068|208|0.613961277758128|0|26|87|-80.80146|13|35.17739|CHEESE CRACKERS|1.01|1|CHEEZ-IT SCRABBLE JUNIOR|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|0.61471665291522548|00024100789351|CRACKERS|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|a052ca082a6510957aeff14926aecfbbe17c4983|5.49|2015-02-23 12:52:00|1.4094857484078087|2|7346102108|208|0.613961277758128|0|26|291|-80.80146|48|35.17739|FROZEN POUTLRY|1.5|5|BARBER F.F. BROCCOLI & CHEESE|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|0.61471665291522548|00073461908758|FROZEN MEALS|FROZEN|-80.80146|1.4102515174184975|208|1
35.17739|bed1165b14fc3f5af12418514b48b86552f33121|6.49|2014-12-07 17:47:00|1.4094857484078087|2|8520000101|208|0.613961277758128|0|26|9922|-80.80146|880|35.17739|NFS-COOLERS|0.0|13|N/A SUTTER HOME FRE CHARDONNAY|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|0.61471665291522548|00085200001019|BEVERAGE|WINE|-80.80146|1.4102515174184975|208|1
35.17739|22c619490aa232415d1d8c80d9f2ac8080def682|3.89|2015-02-05 13:34:00|1.4094857484078087|2|7203695502|208|0.613961277758128|0|26|1693|-80.80146|385|35.17739|CROISSANTS|0.0|14|ARTISAN BUTTER CROISSANTS|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|0.61471665291522548|00072036955029|SWEET GOODS|BAKERY|-80.80146|1.4102515174184975|208|1
35.17739|f930a456bae8ebd363e8a9039d1bf5b5336c85c7|3.79|2014-12-28 16:51:00|80.801203185414451|2|4470000063|208|35.188908061085527|0|24|359|-80.85013|101|35.175855|MEAT WIENERS|0.0|19|OSCAR MAYER SELECTS TURKEY FRK|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|35.194272495053255|00044700007440|WIENERS|CASE READY MEATS|-80.80146|80.801463330337285|218|1
35.17739|07ced3186d75edbfffd27d0dc5948bcd999b2a5c|8.99|2014-12-24 14:45:00|80.801203185414451|2|7069002336|208|35.188908061373944|0|24|757|-80.826724|3|35.195689|BAKING NUTS|3.0|1|FISHER PECAN CHOPPED|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|35.194272495053255|00070690023368|BAKING SUPPLIES|G1 GROCERY|-80.80146|80.801461070058423|412|1
35.17739|cd28f0ef6658d8b5d951f24f357c45a43503ef37|5.79|2014-11-15 14:07:00|1.4094857484078087|2|7069002333|208|0.613961277758128|0|26|757|-80.80146|3|35.17739|BAKING NUTS|1.8|1|FISHER PECAN HALVES|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|0.61471665291522548|00070690023313|BAKING SUPPLIES|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|92a5009983a97a62637ce736732f62bb766fbc8e|2.9|2015-02-28 11:29:00|1.4094857484078087|2|7056097811|208|0.613961277758128|0|26|1272|-80.80146|50|35.17739|BAG VEG STEAM|0.22999999999999998|5|PCTSWT STEAM EDAMAME/SEA SALT|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|0.61471665291522548|00070560977715|VEGETABLES-FROZEN|FROZEN|-80.80146|1.4102515174184975|208|2
35.17739|e53af43d481e1296152a13ae5bc2f01f4347f7ba|3.99|2015-03-09 14:23:00|80.801203185414451|2|7047046118|208|35.188908061373944|0|24|682|-80.826724|61|35.195689|KIDS|0.0|3|YOPLAIT STRWBRY COTTN CNDY 8PK|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|35.194272495053255|00070470461182|YOGURT|DAIRY|-80.80146|80.801461070058423|412|1
35.17739|de94d59cd824951b68acc66976a5022534c663bd|4.99|2014-11-21 11:18:00|80.801203185414451|2|71575620002|208|35.188908060643925|0|24|504|-80.825175|64|35.152722|FRESH BERRIES|0.0|4|STRAWBERRIES 1LB CLAM|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|35.194272495053255|00033383200330|FRESH PRODUCE|PRODUCE|-80.80146|80.801465130273954|160|1
35.17739|1684ee10aec58c48f5ef4f5145b6551aa032c072|3.69|2014-09-14 17:24:00|1.4094857484078087|2|71514172928|208|0.613961277758128|0|26|330|-80.80146|55|35.17739|EGGS|1.69|3|EGGLAND BEST GRADE A EX-LG EGG|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|0.61471665291522548|00715141729283|EGGS FRESH|DAIRY|-80.80146|1.4102515174184975|208|1
35.17739|5838aae76f79a753f8085da0189130d70c1ff1b6|0.6|2014-10-26 17:34:00|1.4094857484078087|2||208|0.613961277758128|0|26|524|-80.80146|64|35.17739|FRESH PROD FRESH ONIONS|0.0|4|COO YELLOW ONIONS, LRG|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|0.61471665291522548|00204665000003|FRESH PRODUCE|PRODUCE|-80.80146|1.4102515174184975|208|1
35.17739|3048c3e2d82c1ce83e320173ee281690ddcc4b32|3.69|2015-03-04 17:19:00|1.4094857484078087|2|7940042833|208|0.613961277758128|0|26|3536|-80.80146|1045|35.17739|SHAMPOO-PREMIUM|0.0|17|SUAVE SA FIRM CONTRL SCULPTGEL|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|0.61471665291522548|00079400428332|HAIR & SCALP CARE|HBC|-80.80146|1.4102515174184975|208|1
35.17739|5e0b6f1ef72e5ec2b77ba38db0b231496e12946f|3.94|2014-12-04 16:43:00|1.4094857484078087|2|7203614993|208|0.613961277758128|0|26|105|-80.80146|16|35.17739|FRUIT CUPS AND GELS|0.0|1|HT 4PK FRT CUP MANDARIN|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|0.61471665291522548|00072036980564|FRUIT-CAN/JAR|G1 GROCERY|-80.80146|1.4102515174184975|208|2
35.17739|9db3c116f8c591fa548920b8eb9d9040723af0ec|3.94|2014-10-08 14:50:00|80.801203185414451|2|7203614993|208|35.188908060485694|0|24|105|-80.810056|16|35.219587|FRUIT CUPS AND GELS|0.0|1|HT 4PK FRT CUP MANDARIN|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|35.194272495053255|00072036980564|FRUIT-CAN/JAR|G1 GROCERY|-80.80146|80.801465637051834|401|2
35.17739|85ef7f9dc8a5fc33a021543ec83488c44e03ce92|1.49|2014-09-27 11:36:00|80.801203185414451|2|4400003211|208|35.188908061085527|0|24|1252|-80.85013|12|35.175855|LUNCH BOX COOKIES|0.49|1|NABISCO GO CUPS NUTTER BUTTER|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|35.194272495053255|00044000032104|COOKIES|G1 GROCERY|-80.80146|80.801463330337285|218|1
35.17739|475ceddd01ae73ebaaa57f1af4de4773ce91c40b|3.99|2015-03-07 16:23:00|1.4094857484078087|2|1600027534|208|0.613961277758128|0|26|81|-80.80146|9|35.17739|RTE CEREAL KIDS|0.0|1|GM LUCKY CHARMS  11.5OZ|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|0.61471665291522548|00016000275348|CEREAL|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|90210642e3dda9b5a77e38eaab004a4ac9ce23cd|3.69|2014-10-28 16:15:00|80.801203185414451|2|7374401050|208|35.188908061085527|0|24|1269|-80.85013|41|35.175855|BREAKFAST SYRUP CARRIER|0.0|5|MURRY'S FRENCH TOAST STICK|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|35.194272495053255|00073744010505|BREAKFAST FOODS FROZEN|FROZEN|-80.80146|80.801463330337285|218|1
35.17739|342319f8946435d0508425af5a3e934189b88036|2.45|2014-12-06 10:31:00|1.4094857484078087|2|7203663217|208|0.613961277758128|0|26|330|-80.80146|55|35.17739|EGGS|0.0|3|HT GRADE A LARGE EGGS 18 CT|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|0.61471665291522548|00072036632173|EGGS FRESH|DAIRY|-80.80146|1.4102515174184975|208|1
35.17739|6054c83d444be547a05494800ffea441849a2113|1.99|2015-03-06 16:45:00|80.801203185414451|2|7203688096|208|35.188908060572864|0|24|526|-80.849471|64|35.161696|FRESH MUSHROOMS|0.0|4|HT SLICED WHITE MUSHROOMS|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|35.194272495053255|00072036880963|FRESH PRODUCE|PRODUCE|-80.80146|80.80146536377697|35|1
35.17739|0d49834f768b905aae19371b20846cbeb67d279f|8.29|2014-11-25 12:02:00|1.4094857484078087|2|4110001511|208|0.613961277758128|0|26|4243|-80.80146|1200|35.17739|NASAL PRODUCT-ADULT|0.0|17|AFRIN NO-DRIP SINUS -01509|4e2ce5b1243237a9a7ddadae6384ba68af858795|0.795870228111187|0.61471665291522548|00041100015099|COUGH/COLD/SINUS|HBC|-80.80146|1.4102515174184975|208|1
35.341927|4a110db3fa55bd07d6c8972ef3a5ee9fc72a0b20|3.18|2014-11-16 13:40:00|80.780380710856576|3|7581037101|220|35.357990124905804|0|48|1217|-80.780702|273|35.318911|ASIAN MEAL KITS/MW|0.0|1|SAN J SOUP PKT WHITE MISO|518eb5df5f1341df7e8a1eb31b0de2691d963dd4|1.1099231942190217|35.351085445956379|00075810371015|ASIAN PREP. FOODS|G1 GROCERY|-80.764523|80.764529159517309|167|2
35.341927|2022d5feef1fa7df72033b1c2cc0d18eac6dfdaa|9.69|2014-10-19 11:28:00|1.4102725052409182|3|88133400051|220|0.6168329901494819|0|1|36|-80.764523|10|35.341927|PREMIUM GROUND|3.7|1|DUNKIN'D FRENCH VANILLA GROUND|518eb5df5f1341df7e8a1eb31b0de2691d963dd4|1.1099231942190217|0.61833652052202714|00881334000474|COFFEE|G1 GROCERY|-80.764523|1.4096068451526882|220|1
35.341927|4196aac0025bbd8708202beea95cc79c774a0ac7|1.69|2014-10-04 18:09:00|1.4102725052409182|3|7203688003|220|0.6168329901494819|0|1|527|-80.764523|64|35.341927|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|518eb5df5f1341df7e8a1eb31b0de2691d963dd4|1.1099231942190217|0.61833652052202714|00072036880031|FRESH PRODUCE|PRODUCE|-80.764523|1.4096068451526882|220|1
35.341927|5f54860225d57d1156135c80da52127271576f2c|2.69|2014-10-26 16:02:00|1.4102725052409182|3|5210007114|220|0.6168329901494819|0|1|1245|-80.764523|34|35.341927|SINGLE SPICES|0.0|1|MC PARSLEY FLAKES|518eb5df5f1341df7e8a1eb31b0de2691d963dd4|1.1099231942190217|0.61833652052202714|00052100071145|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.764523|1.4096068451526882|220|1
35.341927|25800ee56264cfe55aa6663e847040c9f2507010|3.79|2015-02-28 17:21:00|1.4102725052409182|3|7097800832|220|0.6168329901494819|0|1|899|-80.764523|205|35.341927|KOSHER FROZEN FOODS|0.4|5|KINERET COFFEE WHITENER|518eb5df5f1341df7e8a1eb31b0de2691d963dd4|1.1099231942190217|0.61833652052202714|00070978008322|FROZEN KOSHER|FROZEN|-80.764523|1.4096068451526882|220|1
35.341927|3e46989a7e536b602e51c8a4116c4a3a959e206a|7.58|2015-01-17 13:52:00|1.4102725052409182|3|7097800832|220|0.6168329901494819|0|1|899|-80.764523|205|35.341927|KOSHER FROZEN FOODS|0.8|5|KINERET COFFEE WHITENER|518eb5df5f1341df7e8a1eb31b0de2691d963dd4|1.1099231942190217|0.61833652052202714|00070978008322|FROZEN KOSHER|FROZEN|-80.764523|1.4096068451526882|220|2
35.341927|e470d7c804ab3c8070f245296f497e79650bdb57|3.49|2015-02-21 14:40:00|1.4102725052409182|3|7203683254|220|0.6168329901494819|0|1|362|-80.764523|102|35.341927|PEPPERONIS|0.52|19|HT TURKEY PEPPERONI|518eb5df5f1341df7e8a1eb31b0de2691d963dd4|1.1099231942190217|0.61833652052202714|00072036832559|LUNCHMEATS|CASE READY MEATS|-80.764523|1.4096068451526882|220|1
35.341927|954017e9697f5bea58e959dcd2ec166ac74d5795|4.99|2015-01-04 15:18:00|1.4102725052409182|3|7203688012|220|0.6168329901494819|0|1|531|-80.764523|64|35.341927|FRESH CORN|0.0|4|HT PACKAGED WHITE CORN|518eb5df5f1341df7e8a1eb31b0de2691d963dd4|1.1099231942190217|0.61833652052202714|00072036880123|FRESH PRODUCE|PRODUCE|-80.764523|1.4096068451526882|220|1
35.341927|125aa7e0d8fea31d995480e97b384ba7935adc9e|3.49|2015-02-16 15:48:00|1.4102725052409182|3|7203688136|220|0.6168329901494819|0|1|556|-80.764523|64|35.341927|PACKAGED VEGETABLES|0.0|4|HT CELERY STICKS, AQUA PACK|518eb5df5f1341df7e8a1eb31b0de2691d963dd4|1.1099231942190217|0.61833652052202714|00072036881366|FRESH PRODUCE|PRODUCE|-80.764523|1.4096068451526882|220|1
35.341927|577e58b7a9639757e2a22045ed9d8662399e10ec|3.15|2014-12-20 09:31:00|1.4102725052409182|3||220|0.6168329901494819|0|1|523|-80.764523|64|35.341927|FRESH POTATOES|1.95|4|COO SWEET POTATOES, BULK|518eb5df5f1341df7e8a1eb31b0de2691d963dd4|1.1099231942190217|0.61833652052202714|00204091000004|FRESH PRODUCE|PRODUCE|-80.764523|1.4096068451526882|220|1
35.341927|fbad16ce7bd2dee4703aae667510328f86bc4ae3|2.69|2015-01-20 18:27:00|1.4102725052409182|3||220|0.6168329901494819|0|1|523|-80.764523|64|35.341927|FRESH POTATOES|0.0|4|COO SWEET POTATOES, BULK|518eb5df5f1341df7e8a1eb31b0de2691d963dd4|1.1099231942190217|0.61833652052202714|00204091000004|FRESH PRODUCE|PRODUCE|-80.764523|1.4096068451526882|220|1
35.341927|3dad1bb2c3638b1b45800f3340a4e611763265ba|4.19|2015-01-31 17:23:00|1.4102725052409182|3|1920089341|220|0.6168329901494819|0|1|404|-80.764523|69|35.341927|NFS-TOILET BOWL CLEANERS|2.09|1|LYSOL NO MESS WAND-LAVENDER|518eb5df5f1341df7e8a1eb31b0de2691d963dd4|1.1099231942190217|0.61833652052202714|00019200893428|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.764523|1.4096068451526882|220|1
35.341927|c7c50146f6fb742070020ece14e4ac8cbf455444|3.49|2014-11-28 18:44:00|1.4102725052409182|3|64034401620|220|0.6168329901494819|0|1|556|-80.764523|64|35.341927|PACKAGED VEGETABLES|0.0|4|DICED CELERY/ONIONS|518eb5df5f1341df7e8a1eb31b0de2691d963dd4|1.1099231942190217|0.61833652052202714|00640344021523|FRESH PRODUCE|PRODUCE|-80.764523|1.4096068451526882|220|1
35.341927|714089002224a841bfebb6ac536fd70a7c1ef4c0|3.49|2015-01-10 16:21:00|1.4102725052409182|3|7203688133|220|0.6168329901494819|0|1|556|-80.764523|64|35.341927|PACKAGED VEGETABLES|0.0|4|HT FAJITA MIX|518eb5df5f1341df7e8a1eb31b0de2691d963dd4|1.1099231942190217|0.61833652052202714|00072036881335|FRESH PRODUCE|PRODUCE|-80.764523|1.4096068451526882|220|1
35.341927|1b4d036be0c8cf755e940858d4b7dae4a6f32c60|8.0|2014-11-03 17:07:00|1.4102725052409182|3|7203698753|220|0.6168329901494819|0|1|1272|-80.764523|50|35.341927|BAG VEG STEAM|4.0|5|HT RDY QUK BROCCOLI BLEND|518eb5df5f1341df7e8a1eb31b0de2691d963dd4|1.1099231942190217|0.61833652052202714|00072036987518|VEGETABLES-FROZEN|FROZEN|-80.764523|1.4096068451526882|220|4
35.341927|1bc784f6cdca1eff98b84ad3782e529c6dd7efb2|8.99|2014-12-14 17:20:00|1.4102725052409182|3|75703700002|220|0.6168329901494819|0|1|1513|-80.764523|66|35.341927|NFS-LAUNDRY DETERGENT PODS|3.0|1|OXICLEAN DETG FRESH SCENT|518eb5df5f1341df7e8a1eb31b0de2691d963dd4|1.1099231942190217|0.61833652052202714|00757037000113|DETERGENTS|G1 GROCERY|-80.764523|1.4096068451526882|220|1
35.341927|45ac6b39042f5d6c2ef61aaf1883a9e2cf61fe14|13.58|2014-10-27 16:44:00|1.4102725052409182|3|7800001180|220|0.6168329901494819|0|1|54|-80.764523|8|35.341927|DIET|3.4|23|CD DT GINGER ALE 12PK|518eb5df5f1341df7e8a1eb31b0de2691d963dd4|1.1099231942190217|0.61833652052202714|00078000148169|CARBONATED BEVERAGES|BEVERAGE|-80.764523|1.4096068451526882|220|2
35.341927|04a70a38bf9b26d532a3f279014f430a171c43da|14.549999999999999|2014-11-04 17:42:00|1.4102725052409182|3|7790011553|220|0.6168329901494819|0|1|361|-80.764523|105|35.341927|BREAKFAST SAUSAGE|1.51|19|JIMMY DEAN HOT SAUSAGE|518eb5df5f1341df7e8a1eb31b0de2691d963dd4|1.1099231942190217|0.61833652052202714|00077900115639|BREAKFAST SAUSAGE|CASE READY MEATS|-80.764523|1.4096068451526882|220|3
35.341927|bc7672bb613495af4d0a00530dc86f8f64e24a61|2.69|2015-02-23 18:49:00|1.4102725052409182|3|7203688023|220|0.6168329901494819|0|1|555|-80.764523|64|35.341927|PACKAGED SALADS|0.0|4|HT CURLY SPINACH,PKG|518eb5df5f1341df7e8a1eb31b0de2691d963dd4|1.1099231942190217|0.61833652052202714|00072036880239|FRESH PRODUCE|PRODUCE|-80.764523|1.4096068451526882|220|1
35.103409|f24553f03d2d86757883bb809992a44e7feb9ec5|9.49|2015-03-08 13:16:00|1.4132775322775095|2|5400011971|88|0.6126700657242101|0|58|427|-80.992182|72|35.103409|NFS-TOILET TISSUE|3.5|1|SCOTT 1000 WHITE 8 ROLL|535feb5d5170f703c8df0928885a1770380055e5|1.7961688315973723|0.61177642288969325|00054000119712|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|a65e3c7c8074a4392d417a6c3abbca175a142829|3.58|2014-11-02 16:05:00|1.4132775322775095|2|2000011274|88|0.6126700657242101|0|58|245|-80.992182|39|35.103409|VEGETABLES-CORE|0.0|1|GREEN GIANT CORN WHITE SHOEPEG|535feb5d5170f703c8df0928885a1770380055e5|1.7961688315973723|0.61177642288969325|00020000105468|VEGETABLES-CAN/JAR|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|323f9c64570f98d1beec54071834f8ea56ae5f8b|3.19|2014-10-25 15:38:00|1.4132775322775095|2|82951530146|88|0.6126700657242101|0|58|205|-80.992182|31|35.103409|REMAINING SNACKS|1.6|1|SENSBL STRAW CINNAMON APPLE|535feb5d5170f703c8df0928885a1770380055e5|1.7961688315973723|0.61177642288969325|00829515302818|SNACKS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|289363d469c24473fc205d3dc1ed027c5f591ad6|5.94|2014-09-13 12:17:00|1.4132775322775095|2|4173600180|88|0.6126700657242101|0|58|194|-80.992182|30|35.103409|OLIVE OIL|3.0|1|FILIPPO BERIO PURE OLIVE OIL|535feb5d5170f703c8df0928885a1770380055e5|1.7961688315973723|0.61177642288969325|00041736001800|SHORTENING/OIL|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|ef20bc0d81d2156bb76eab36c52b1bda1a30f172|1.99|2015-02-28 12:08:00|1.4132775322775095|2|7680828073|88|0.6126700657242101|0|58|149|-80.992182|23|35.103409|WHSE PASTA CORE|1.99|1|BARILLA PASTA ELBOWS|535feb5d5170f703c8df0928885a1770380055e5|1.7961688315973723|0.61177642288969325|00076808516135|PASTA|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|d8ca5ec5154ceb4d15e81589bb330d2a90b69980|4.98|2015-01-03 14:33:00|1.4132775322775095|2|20337700000|88|0.6126700657242101|0|58|641|-80.992182|137|35.103409|PREMIUM PORK|0.0|2|PORK LOIN CHOPS BNLS THIN|535feb5d5170f703c8df0928885a1770380055e5|1.7961688315973723|0.61177642288969325|00203377000004|PORK|MEAT|-80.992182|1.413580244274486|88|1
35.103409|a89def609151a1ebc23a2d64e3eea0486deb2343|1.49|2014-12-14 14:06:00|1.4132775322775095|2|7203653022|88|0.6126700657242101|0|58|1273|-80.992182|50|35.103409|BAG VEG NON STEAM|0.0|5|HT CUT OKRA|535feb5d5170f703c8df0928885a1770380055e5|1.7961688315973723|0.61177642288969325|00072036537522|VEGETABLES-FROZEN|FROZEN|-80.992182|1.413580244274486|88|1
35.103409|dbdb6dccfe738f3a47e46203032297784eeb5eb5|2.99|2015-01-31 17:40:00|1.4132775322775095|2|7027223202|88|0.6126700657242101|0|58|323|-80.992182|57|35.103409|TOPPINGS-REFRIGERATED|0.0|3|REDDI WIP EXTRA CREAMY|535feb5d5170f703c8df0928885a1770380055e5|1.7961688315973723|0.61177642288969325|00070272232034|MILK|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|17d41b77baeb5cef542ff5b9fb0b17786bca5ddb|2.99|2014-11-27 09:21:00|1.4132775322775095|2|2529360050|88|0.6126700657242101|0|58|339|-80.992182|57|35.103409|EGGNOGS/DRINKS|0.3|3|I/O SILK NOG|535feb5d5170f703c8df0928885a1770380055e5|1.7961688315973723|0.61177642288969325|00025293600508|MILK|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|0068e575392b1987d6375c9e768be2d36e2abd65|6.63|2014-12-17 14:01:00|1.4132775322775095|2|20896500000|88|0.6126700657242101|0|58|977|-80.992182|201|35.103409|FRESH HT CHICKEN|0.0|2|HT FRESH CHICKEN DRUMMETTES|535feb5d5170f703c8df0928885a1770380055e5|1.7961688315973723|0.61177642288969325|00208965000008|POULTRY|MEAT|-80.992182|1.413580244274486|88|2
35.103409|6e2c46becbebae68f2a8dd593d9a6bbce2961858|13.33|2014-09-25 17:20:00|1.4132775322775095|2|20557100000|88|0.6126700657242101|0|58|1820|-80.992182|410|35.103409|BH BEEF|0.0|6|BOARS HEAD LONDON BROIL|535feb5d5170f703c8df0928885a1770380055e5|1.7961688315973723|0.61177642288969325|00205571000002|BH MEAT|DELI|-80.992182|1.413580244274486|88|1
35.103409|47a530003b214ea3b0fdf71eec183ce76e871334|3.39|2014-09-17 12:38:00|1.4132775322775095|2|4610000107|88|0.6126700657242101|0|58|331|-80.992182|52|35.103409|NATURAL SLICED|0.0|3|SARGENTO EXTRA SHARP SLICE|535feb5d5170f703c8df0928885a1770380055e5|1.7961688315973723|0.61177642288969325|00046100002728|CHEESE|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|343fcdb31ab727b1742a219e3c74e93d0d895171|5.49|2014-10-14 17:54:00|1.4132775322775095|2|74016901887|88|0.6126700657242101|0|58|661|-80.992182|144|35.103409|MEAT CONDIMENTS MARINADE|1.5|2|PETER LUGER NEW YORK STEAK SAU|535feb5d5170f703c8df0928885a1770380055e5|1.7961688315973723|0.61177642288969325|00740169018873|CONDIMENTS|MEAT|-80.992182|1.413580244274486|88|1
35.103409|c324db4ceb749f9984e194d02be3b79edda2a536|27.26|2014-09-21 14:20:00|1.4132775322775095|2|20237100000|88|0.6126700657242101|0|58|299|-80.992182|49|35.103409|ANGUS BEEF|6.82|2|ANGUS BEEF ROUND LONDON BROIL|535feb5d5170f703c8df0928885a1770380055e5|1.7961688315973723|0.61177642288969325|00202371000003|BEEF|MEAT|-80.992182|1.413580244274486|88|2
35.103409|d480fea51035baca4a3c13a87a6917b85776a4a9|4.99|2014-11-15 19:09:00|1.4132775322775095|2|7529506050|88|0.6126700657242101|0|58|275|-80.992182|45|35.103409|SUPER PREMIUM ICE CREAM|0.0|5|FRONT PORCH CHOC ROCKER IC|535feb5d5170f703c8df0928885a1770380055e5|1.7961688315973723|0.61177642288969325|00075295060534|ICE CREAM|FROZEN|-80.992182|1.413580244274486|88|1
35.103409|68883cb9d0625cf33dfd421d24e24c89a163612e|9.99|2015-01-28 16:27:00|1.4132775322775095|2|84105802208|88|0.6126700657242101|0|58|3917|-80.992182|1075|35.103409|DISPOSABLE RAZOE-MEN|0.0|17|QUATTRO MENS DISP RAZOR SENS|535feb5d5170f703c8df0928885a1770380055e5|1.7961688315973723|0.61177642288969325|00841058022084|SHAVING NEEDS/MEN HAIR|HBC|-80.992182|1.413580244274486|88|1
35.103409|80b4ba4afb0cac9ab4c93016fc8166570da12cd5|4.99|2014-09-26 19:33:00|1.4132775322775095|2|7529506050|88|0.6126700657242101|0|58|275|-80.992182|45|35.103409|SUPER PREMIUM ICE CREAM|1.49|5|FRONT PORCH MTN MINT CHIP IC|535feb5d5170f703c8df0928885a1770380055e5|1.7961688315973723|0.61177642288969325|00075295060565|ICE CREAM|FROZEN|-80.992182|1.413580244274486|88|1
35.103409|5436f45110bae5f9ef796cb6c02d2dcecf623a86|0.99|2015-02-12 11:59:00|1.4132775322775095|2|7203695306|88|0.6126700657242101|0|58|1895|-80.992182|450|35.103409|TEA|0.0|6|FFM LEMONADE|535feb5d5170f703c8df0928885a1770380055e5|1.7961688315973723|0.61177642288969325|00072036953070|BEVERAGES|DELI|-80.992182|1.413580244274486|88|1
35.103409|7925a1e36c660cd2d9c8917cc7df6297960aba52|6.79|2014-10-25 20:24:00|1.4132775322775095|2|7064003404|88|0.6126700657242101|0|58|252|-80.992182|45|35.103409|PREMIUM ICE CREAM|2.81|5|B BUNNY PREM PISTACHIO ALMOND|535feb5d5170f703c8df0928885a1770380055e5|1.7961688315973723|0.61177642288969325|00070640034192|ICE CREAM|FROZEN|-80.992182|1.413580244274486|88|1
35.323246|57efbb9b9939d91eb544ecb8e54458dbc710d70c|3.56|2015-01-05 18:55:00|80.945255278477163|4||166|35.384513767490162|0|13|566|-80.810056|64|35.219587|SERVICE BAR|0.25|4|HT SPINACH DIP|5411c661151caf7f1dc9c2a2a3e2d2b95e6141db|4.23345523465759|35.37387923947206|00204376000002|FRESH PRODUCE|PRODUCE|-80.945176|80.945210921822735|401|1
35.40953|2852054eaeb9bcf33896ed7a144f34e67484a33e|3.19|2014-10-29 13:18:00|80.86161257435397|4|82951530146|209|35.439006824749661|0|36|205|-80.80146|31|35.17739|REMAINING SNACKS|1.59|1|SENSBL PORT VEG STRAW RS OLV O|5571da260daa6c3db0373fe42d37e188031f70c1|2.0367820653285995|35.472272108304431|00829515302108|SNACKS|G1 GROCERY|-80.86175|80.861827371454851|208|1
35.40953|790f9f396e478be49cc94b60903b57be217bba1c|3.89|2014-12-12 17:08:00|80.86161257435397|4|2100012277|209|35.439006798614464|0|36|320|-80.849471|53|35.161696|COTTAGE CHEESE|0.0|3|BREAKSTONE 2% COTTAGE CHEESE|5571da260daa6c3db0373fe42d37e188031f70c1|2.0367820653285995|35.472272108304431|00021000123544|CULTURES|DAIRY|-80.86175|80.861841140846906|35|1
35.40953|69cc7ddb5595dcc951d6d709ed1fd098892838f5|5.99|2015-01-06 21:11:00|80.86161257435397|4|2858800340|209|35.439006809025152|0|36|5846|-80.85013|1538|35.175855|KITCHEN GADGETS BARWARE|1.0|18|(JHK) WAITERS CORKSCREW|5571da260daa6c3db0373fe42d37e188031f70c1|2.0367820653285995|35.472272108304431|00028588003404|KITCHEN GADGETS|GM|-80.86175|80.861835920789972|218|1
35.40953|df6687985477ce367ebf5023ce828f336d170bb6|2.69|2015-01-31 20:34:00|80.86161257435397|4|70935100013|209|35.439006809025152|0|36|556|-80.85013|64|35.175855|PACKAGED VEGETABLES|0.0|4|APIO BROCCOLI & CARROTS|5571da260daa6c3db0373fe42d37e188031f70c1|2.0367820653285995|35.472272108304431|00709351000256|FRESH PRODUCE|PRODUCE|-80.86175|80.861835920789972|218|1
35.444064|f9ee3db6abcb8ad8caf4ce8e66d805d7e1a9dfa1|2.69|2014-09-30 17:33:00|1.4102725052409182|4|7203663996|121|0.6186156170875914|0|1|342|-80.995484|57|35.444064|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00072036631299|MILK|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|8ab17f99192145988fad59b1b73fed6435183161|2.69|2014-09-15 18:16:00|1.4102725052409182|4|7203663996|121|0.6186156170875914|0|1|342|-80.995484|57|35.444064|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00072036631299|MILK|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|443d4b270d1b538788aa02ac0b1127f604d3f686|2.29|2015-02-25 18:32:00|1.4102725052409182|4|7203663996|121|0.6186156170875914|0|1|342|-80.995484|57|35.444064|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00072036631299|MILK|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|1bd3f55faa280675fcad9f7fd666c1a67eef3607|2.59|2014-11-07 17:25:00|1.4102725052409182|4|7203663996|121|0.6186156170875914|0|1|342|-80.995484|57|35.444064|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00072036631299|MILK|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|65c8169de9562a9467529f9906a009cbd6561cdf|2.29|2015-01-15 17:48:00|1.4102725052409182|4|7203663996|121|0.6186156170875914|0|1|342|-80.995484|57|35.444064|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00072036631299|MILK|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|2c9f3283a3b417d0b8af79260443ef4d6d3f041e|1.95|2014-11-10 16:23:00|1.4102725052409182|4|930000011|121|0.6186156170875914|0|1|161|-80.995484|25|35.444064|PEPPERS|0.0|1|MT OLV JALAPENO DICED|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00009300000161|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|cb7fe010772c4efd027397c262c7b14bbd94447d|1.79|2014-10-29 19:17:00|1.4102725052409182|4|5100001047|121|0.6186156170875914|0|1|212|-80.995484|33|35.444064|CONDENSED SOUP|0.79|1|CAMP COND MINESTRONE|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00051000011411|SOUP|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|cca0d0c59f2a3766b35a0e9f2122c8d70bdef07b|4.78|2014-12-16 14:32:00|80.995508130988839|4|5100002379|121|35.465223180906619|1|40|173|-80.945176|27|35.323246|CANNED POULTRY|0.78|1|SWANSON CANNED CHICKEN 4.5 OZ|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|35.466476270328783|00051000023797|PREPARED FOODS-RTS|G1 GROCERY|-80.995484|80.995510625946551|166|2
35.444064|e0b666a9f4cc55fd0bf1bf7e5328c095ac10c52f|3.0|2014-10-21 10:47:00|1.4102725052409182|4||121|0.6186156170875914|0|1|531|-80.995484|64|35.444064|FRESH CORN|0.0|4|COO YELLOW CORN|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00204078000003|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|5
35.444064|f57f2692a0623b64ce12015ca44a42feb269c32c|3.25|2015-01-12 14:54:00|1.4102725052409182|4|7203656080|121|0.6186156170875914|0|1|318|-80.995484|52|35.444064|SHREDDED/GRATED CHEESE|0.0|3|HT SHRED MOZZARELLA CHEESE 2%|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00072036000194|CHEESE|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|579a1759954da8ea9472ca3ba086b6865e80a522|1.99|2014-10-16 13:13:00|1.4102725052409182|4|3900004504|121|0.6186156170875914|0|1|114|-80.995484|14|35.444064|PUMPKIN|0.0|1|LIBBY SOLID PACK PUMPKIN|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00039000045049|DESSERTS/GELS/SYRUPS|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|945e0c05dd14fb7252d9d2db4d25dff827f18eb3|1.29|2014-11-24 18:25:00|1.4102725052409182|4|3940001810|121|0.6186156170875914|0|1|242|-80.995484|39|35.444064|CANNED BEANS|0.29|1|BUSH BEAN MIXED|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00039400017707|VEGETABLES-CAN/JAR|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|ef5e55a19ef438432dad34536930908eef20bb27|3.19|2015-02-01 15:32:00|1.4102725052409182|4|5000062231|121|0.6186156170875914|0|1|326|-80.995484|54|35.444064|COOKIES/BROWNIES-REFRIGERATED|0.69|3|NESTLE WHT CHOC CHIP MACADAMIA|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00050000009237|DOUGH PRODUCTS|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|19c9f06795b5f2559a8c79ef8fd23ae2388cbc66|2.0|2015-02-12 18:43:00|1.4102725052409182|4|5100002549|121|0.6186156170875914|0|1|1221|-80.995484|275|35.444064|PASTA SC VALUE|0.33|1|PREGO SC TRADITIONAL|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00051000025494|PASTA SAUCES|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|2e62fff55fd34c091cad6d9aca1de13e8e818fec|2.99|2015-02-02 18:11:00|1.4102725052409182|4|1380004717|121|0.6186156170875914|0|1|1278|-80.995484|48|35.444064|SINGLE SERVE NUTRITIONAL|0.0|5|LC CAFE CLSSC PEPPERONI PIZZA|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00013800047175|FROZEN MEALS|FROZEN|-80.995484|1.413637875046387|121|1
35.444064|980c97a029eb7e6c0d9e98f3f5d527a3bb7d9fea|1.39|2015-01-31 12:27:00|1.4102725052409182|4|5210094269|121|0.6186156170875914|0|1|80|-80.995484|34|35.444064|SEASONING PACKETS|0.39|1|MC MILD CHILI SEASONING MIX|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00052100155203|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|3f4c192df6348859a9a7f208a64d927a3ad54114|3.99|2015-02-25 18:30:00|1.4102725052409182|4|7203602701|121|0.6186156170875914|0|1|1878|-80.995484|435|35.444064|HUMMUS|0.3|6|FFM ARTISAN RED PEPPER HUMMUS|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00072036027030|SALADS|DELI|-80.995484|1.413637875046387|121|1
35.444064|3b9f095cfb7ecfcc4da8ef6a56e1a60130b8e19f|3.99|2015-03-09 14:43:00|1.4102725052409182|4|6055600161|121|0.6186156170875914|0|1|556|-80.995484|64|35.444064|PACKAGED VEGETABLES|0.0|4|CUTBUTTERNUT SQUASH|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00640344020601|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|ff48e6fee199abaa2887099cd727990a2f5a2308|5.26|2014-11-03 18:20:00|1.4102725052409182|4||121|0.6186156170875914|0|1|500|-80.995484|64|35.444064|FRESH APPLES|1.09|4|HONEY CRISP APPLE|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00233283000003|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|2
35.444064|476731d9b118e77cb180e0d70fa99cc235edc05e|3.65|2014-09-29 18:48:00|1.4102725052409182|4|2529300098|121|0.6186156170875914|0|1|1265|-80.995484|57|35.444064|ALMOND MILK|0.65|3|SILK PURE ALMOND VANILLA LIGHT|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00025293002173|MILK|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|3d87b30b1387aa9dc7a265bc70f42d846a5c06c3|3.65|2014-09-19 21:51:00|1.4102725052409182|4|2529300098|121|0.6186156170875914|0|1|1265|-80.995484|57|35.444064|ALMOND MILK|0.65|3|SILK PURE ALMOND VANILLA LIGHT|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00025293002173|MILK|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|617b9668d3c7e1754f37ec3df9750a10f4e80339|3.49|2015-02-13 15:42:00|1.4102725052409182|4|72243011016|121|0.6186156170875914|0|1|577|-80.995484|136|35.444064|OTHER MERCH FR MSC JUICE|0.0|4|ORG. GT KOMBUCHA MANGO|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00722430500164|OTHER MERCHANDISE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|0c89eac206c566ec22e2c5b5fc75c685f2e53cdf|14.96|2015-02-09 18:32:00|1.4102725052409182|4|20893900000|121|0.6186156170875914|0|1|657|-80.995484|201|35.444064|STR MDE VALUE ADD POLTRY|3.74|2|SPINACH & FETA CHCKN BREAST|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00208939000003|POULTRY|MEAT|-80.995484|1.413637875046387|121|2
35.444064|44cc94fd8a2f83cc23be22302a24276b7fbebae0|3.0|2015-02-22 15:30:00|1.4102725052409182|4|68954408130|121|0.6186156170875914|0|1|685|-80.995484|61|35.444064|GREEK|0.0|3|FAGE 0% WITH HONEY|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00689544081258|YOGURT|DAIRY|-80.995484|1.413637875046387|121|2
35.444064|7241f2529b487deb9090d31a70b8d037e2c51860|3.49|2015-02-15 17:44:00|1.4102725052409182|4|7797508161|121|0.6186156170875914|0|1|204|-80.995484|31|35.444064|TORTILLA CHIPS|0.99|1|SOH RESTURNT STYLE TORTILLA CH|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00077975081785|SNACKS|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|93c292bb232f1b1634148c26bd37122d86b02197|4.19|2014-11-01 12:05:00|1.4102725052409182|4|76026300010|121|0.6186156170875914|0|1|213|-80.995484|33|35.444064|SOUP MIXES|0.0|1|BEAR CREEK SOUP MIX CHED BROCC|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00760263000260|SOUP|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|5fc3ed92145425abd4b8a807a176393d3f3abd50|8.19|2014-09-24 21:13:00|1.4102725052409182|4|2840000288|121|0.6186156170875914|0|1|205|-80.995484|31|35.444064|REMAINING SNACKS|1.2|1|FRITOLAY FLAVOR 20 CTN|58b76af1852e3ba1588792c9da0f3abe6d3de22f|1.4620490711339067|0.61833652052202714|00028400002899|SNACKS|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.006282|d7e83af8b2b0701b172775c376d5378b1b7cbfe1|6.99|2014-11-22 14:31:00|80.562862110758871|3|7468210906|60|35.08247195967833|0|21|128|-80.699686|20|35.000049|APPLE JUICE-SHELF|1.0|1|I/O KNUDSEN CIDER 96 OZ|59f0c7563315a7ba84ec1c492510a1cead89bae3|5.264543458012708|35.054042368968126|00074682109061|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.562829|80.562892779961274|249|1
35.006282|6ba7613752c4ac41e0be756479e71c9bfb197134|3.79|2014-11-16 11:47:00|80.562862110758871|3|7774529186|60|35.08247195967833|0|21|555|-80.699686|64|35.000049|PACKAGED SALADS|0.0|4|R.P. BISTRO CRANBERRY WALNUT|59f0c7563315a7ba84ec1c492510a1cead89bae3|5.264543458012708|35.054042368968126|00077745294131|FRESH PRODUCE|PRODUCE|-80.562829|80.562892779961274|249|1
35.006282|ad839bdc370191ff998655299de331b260dc3e3f|7.58|2014-12-13 18:13:00|80.562862110758871|3|7774529186|60|35.08247195967833|0|21|555|-80.699686|64|35.000049|PACKAGED SALADS|0.0|4|R.P. BISTRO CRANBERRY WALNUT|59f0c7563315a7ba84ec1c492510a1cead89bae3|5.264543458012708|35.054042368968126|00077745294131|FRESH PRODUCE|PRODUCE|-80.562829|80.562892779961274|249|2
35.006282|8a371b16415aa69e86154e13c96dd9441738c7cb|1.16|2015-01-18 11:17:00|1.4091206135396188|3||60|0.6109748797816256|0|47|565|-80.562829|64|35.006282|REDUCED PRODUCE|0.0|4|PRODUCE REWRAP BY LB|59f0c7563315a7ba84ec1c492510a1cead89bae3|5.264543458012708|0.61242566243833529|00204844000008|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|1
35.006282|272f67fd0f52aa78f80b81b3afb74463cc87ac4a|7.99|2014-12-20 16:56:00|80.562862110758871|3|4145810534|60|35.08247195967833|0|21|265|-80.699686|307|35.000049|FROZEN PIES|3.0|5|EDWARDS CHOC CREAM W/HERSHEY'S|59f0c7563315a7ba84ec1c492510a1cead89bae3|5.264543458012708|35.054042368968126|00041458105565|DESSERTS FROZEN|FROZEN|-80.562829|80.562892779961274|249|1
35.006282|3aad14fef9d878e1115ce993276619bc775222e6|7.99|2014-10-11 17:40:00|80.562862110758871|3|4145810534|60|35.08247195967833|0|21|265|-80.699686|307|35.000049|FROZEN PIES|0.0|5|EDWARDS CHOC CREAM W/HERSHEY'S|59f0c7563315a7ba84ec1c492510a1cead89bae3|5.264543458012708|35.054042368968126|00041458105565|DESSERTS FROZEN|FROZEN|-80.562829|80.562892779961274|249|1
35.006282|8e9e788f38c837ad6d9b64b083201e3c521948aa|83.91|2015-02-28 21:06:00|80.562862110758871|3|20324300000|60|35.08247195967833|0|21|641|-80.699686|137|35.000049|PREMIUM PORK|9.0|2|PORK BABY BACK RIBS|59f0c7563315a7ba84ec1c492510a1cead89bae3|5.264543458012708|35.054042368968126|00203243000008|PORK|MEAT|-80.562829|80.562892779961274|249|4
35.006282|2a4ad1eba15467649ed84875a6a6248e2ee7782d|46.93|2014-10-26 13:16:00|80.562862110758871|3|20324300000|60|35.08247195967833|0|21|641|-80.699686|137|35.000049|PREMIUM PORK|11.01|2|PORK BABY BACK RIBS|59f0c7563315a7ba84ec1c492510a1cead89bae3|5.264543458012708|35.054042368968126|00203243000008|PORK|MEAT|-80.562829|80.562892779961274|249|2
35.006282|ef33594f58cdaa887eee14224ea6b428b9d73d21|6.859999999999999|2014-09-20 19:25:00|80.562862110758871|3|20328700000|60|35.08247195967833|0|21|641|-80.699686|137|35.000049|PREMIUM PORK|3.6799999999999997|2|PORK LOIN RIB END CHOPS BNLS|59f0c7563315a7ba84ec1c492510a1cead89bae3|5.264543458012708|35.054042368968126|00203287000002|PORK|MEAT|-80.562829|80.562892779961274|249|2
35.006282|d72ac1b9dcbb8813e33fe4640496eb661f0b1eb1|1.87|2014-11-02 13:35:00|80.562862110758871|3|7203653024|60|35.08247195967833|0|21|1273|-80.699686|50|35.000049|BAG VEG NON STEAM|0.0|5|HT MINI CORN ON THE COB|59f0c7563315a7ba84ec1c492510a1cead89bae3|5.264543458012708|35.054042368968126|00072036530240|VEGETABLES-FROZEN|FROZEN|-80.562829|80.562892779961274|249|1
35.006282|eab15985f544767aba4e4dc711218888d3b19936|3.25|2014-12-06 15:18:00|80.562862110758871|3|7203656080|60|35.08247195967833|0|21|318|-80.699686|52|35.000049|SHREDDED/GRATED CHEESE|0.0|3|HT GOURMENT SHARP BLEND|59f0c7563315a7ba84ec1c492510a1cead89bae3|5.264543458012708|35.054042368968126|00072036600783|CHEESE|DAIRY|-80.562829|80.562892779961274|249|1
35.006282|2445d70e9e650dbdd5d0327146e5f0e24950cafc|27.15|2015-01-11 16:05:00|80.562862110758871|3|20137100000|60|35.08247195967833|0|21|296|-80.699686|49|35.000049|RANCHER BEEF|4.99|2|VALUE PK T-BONE STEAKS|59f0c7563315a7ba84ec1c492510a1cead89bae3|5.264543458012708|35.054042368968126|00201371000006|BEEF|MEAT|-80.562829|80.562892779961274|249|1
35.006282|4e7d800698e4bd21a34a96d0892734da924cda97|3.38|2014-12-31 19:03:00|80.562862110758871|3|73801577715|60|35.08247195967833|0|21|545|-80.699686|64|35.000049|FRESH SPROUTS|0.38|4|BLACK-EYED PEAS, PKG|59f0c7563315a7ba84ec1c492510a1cead89bae3|5.264543458012708|35.054042368968126|00738015777159|FRESH PRODUCE|PRODUCE|-80.562829|80.562892779961274|249|2
35.006282|c6ca0248b4773ed4fea1cf74df2a1e8b7b4e06db|4.98|2015-02-15 15:18:00|80.562862110758871|3|4801400748|60|35.08247195967833|0|21|727|-80.699686|7|35.000049|SEASONAL CANDY-SINGLE FAC|0.98|1|I/O(V15)LOTS OF HEARTS BOUQUET|59f0c7563315a7ba84ec1c492510a1cead89bae3|5.264543458012708|35.054042368968126|00048014009145|CANDY|G1 GROCERY|-80.562829|80.562892779961274|249|2
35.006282|05117a3bcd4e0b664253c7e0c67b02c6043a38d1|9.99|2015-02-14 15:08:00|80.562862110758871|3|78539157005|60|35.08247195967833|0|21|263|-80.699686|307|35.000049|CHEESECAKE FROZEN|0.0|5|BILTMORE VAN BEAN CHEESECAKE|59f0c7563315a7ba84ec1c492510a1cead89bae3|5.264543458012708|35.054042368968126|00785391570058|DESSERTS FROZEN|FROZEN|-80.562829|80.562892779961274|249|1
35.006282|750c66a7c0dc3e944ab4f976b10bb7b5bfe3b92b|6.49|2015-01-24 16:21:00|80.562862110758871|3|5000030302|60|35.08247195967833|0|21|144|-80.699686|229|35.000049|CEAMERS-POWDERED|0.0|1|COFFEE MATE KILO|59f0c7563315a7ba84ec1c492510a1cead89bae3|5.264543458012708|35.054042368968126|00050000303021|COCOAS CREAMERS SYRUPS|G1 GROCERY|-80.562829|80.562892779961274|249|1
35.006282|1920446cd0823220b15671963b1de240621581dc|4.49|2014-12-12 13:59:00|1.4091206135396188|3|7027710520|60|0.6109748797816256|0|47|2020|-80.562829|505|35.006282|CHEESE SPECIALTIES|1.0|6|ATHENOS FETA TRADITIONAL CRMBD|59f0c7563315a7ba84ec1c492510a1cead89bae3|5.264543458012708|0.61242566243833529|00070277105203|SPECIALTY CHEESE|DELI|-80.562829|1.4060866207711706|60|1
35.006282|e0920d202e39917b092f68691b5441cf2b50d37d|15.3|2015-02-07 18:47:00|80.562862110758871|3|76211120604|60|35.08247195967833|0|21|36|-80.699686|10|35.000049|PREMIUM GROUND|1.32|1|STARBUCKS BRKF BLND GRND COFFE|59f0c7563315a7ba84ec1c492510a1cead89bae3|5.264543458012708|35.054042368968126|00762111206251|COFFEE|G1 GROCERY|-80.562829|80.562892779961274|249|2
35.006282|50269ec5d4b447fa267d78526e061a7ba1b0fd99|23.509999999999998|2014-09-25 20:07:00|80.562862110758871|3|20120300000|60|35.082471977542603|0|21|296|-80.732725|49|35.082768|RANCHER BEEF|9.05|2|BEEF RIBEYE STEAK BONELESS|59f0c7563315a7ba84ec1c492510a1cead89bae3|5.264543458012708|35.054042368968126|00201203000006|BEEF|MEAT|-80.562829|80.562831582853661|147|2
35.006282|69ccd76f70c1a76d5cc29f999416f19501461127|1.79|2015-03-08 19:02:00|80.562862110758871|3|2430004107|60|35.08247195967833|0|21|1044|-80.699686|173|35.000049|SW BAKD GOOD SNACK CAKES|0.0|7|LD FUDGE BROWNIE|59f0c7563315a7ba84ec1c492510a1cead89bae3|5.264543458012708|35.054042368968126|00024300041259|SWEET BAKED GOODS|COMMERCIAL BAKERY|-80.562829|80.562892779961274|249|1
35.006282|9a76d91d63b716ecc2bc76353ff121f588fb0a9a|4.99|2014-09-14 17:02:00|1.4091206135396188|3|7203698713|60|0.6109748797816256|0|47|4353|-80.562829|1205|35.006282|SLEEPING AID|0.0|17|HT ACETAMINOPHEN PM CAPLETS|59f0c7563315a7ba84ec1c492510a1cead89bae3|5.264543458012708|0.61242566243833529|00072036987136|PAIN RELIEF|HBC|-80.562829|1.4060866207711706|60|1
35.667941|7a25237924762aae3f5acc6f1199cf8f68c8207c|1.49|2015-02-14 15:12:00|1.4057311447477159|unknown|7156799788|178|0.6225230078570788|0|52|727|-80.497332|7|35.667941|SEASONAL CANDY-SINGLE FAC|0.75|1|I/O(V15)MCKY MINNIE VAL EXCHNG|5b40cab7848d0e7c22c61a50eac9235ca49d4936|2.8532768562543076|0.6209993146566879|00071567997881|CANDY|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|e5f20decf382293ae895fdd8b0daf441663899c1|4.49|2015-03-08 15:54:00|1.4057311447477159|unknown|3000006442|178|0.6225230078570788|0|52|61|-80.497332|9|35.667941|RTE CEREAL ADULT|1.99|1|QUAKER OATMEAL SQ HONEY NUT|5b40cab7848d0e7c22c61a50eac9235ca49d4936|2.8532768562543076|0.6209993146566879|00030000313282|CEREAL|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|b95502e8910a15c094e6880c9e5a666b6f189b75|2.85|2015-03-05 12:35:00|1.4057311447477159|unknown|4400000055|178|0.6225230078570788|0|52|88|-80.497332|13|35.667941|FLAKED SODA CRACKERS|0.35|1|NABISCO PREMIUMS|5b40cab7848d0e7c22c61a50eac9235ca49d4936|2.8532768562543076|0.6209993146566879|00044000000578|CRACKERS|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|0f5a8ce70297f6ad44a223446cfd5e20ee622470|1.5|2015-03-04 14:46:00|1.4057311447477159|unknown|7203641160|178|0.6225230078570788|0|52|247|-80.497332|39|35.667941|VEGETABLES-FLANKER|0.0|1|HT MIXED VEGETABLES|5b40cab7848d0e7c22c61a50eac9235ca49d4936|2.8532768562543076|0.6209993146566879|00072036411709|VEGETABLES-CAN/JAR|G1 GROCERY|-80.497332|1.4049434824709919|178|2
35.667941|d241eed09d4b288f45d952dbceea7f517ce1731d|5.49|2015-02-22 17:36:00|1.4057311447477159|unknown|3700035762|178|0.6225230078570788|0|52|417|-80.497332|71|35.667941|NFS-FABRIC SOFTENERS|0.0|1|DOWNY LIQ FAB SOFT CLEAN BREEZ|5b40cab7848d0e7c22c61a50eac9235ca49d4936|2.8532768562543076|0.6209993146566879|00037000393009|LAUNDRY SUPPLIES|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.006282|90f7021ff08d3be8447c6e66fe532e94735c485b|1.69|2014-11-26 11:27:00|80.562862110758871|3|4900000463|60|35.040504021150888|0|21|55|-80.64817|8|35.04711|REGULAR|0.58|23|SPRITE GLASS SINGLE|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00049000047820|CARBONATED BEVERAGES|BEVERAGE|-80.562829|80.562830632871794|129|1
35.006282|37c4609f26872298ec2c681dfdd82fc0d3d780ef|2.99|2015-01-19 17:14:00|80.562862110758871|3|7203659032|60|35.040504021150888|0|21|321|-80.64817|53|35.04711|RICOTTA/FARMERS CHEESE|0.0|3|HT PART SKIM RICOTTA CHEESE|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00072036600370|CULTURES|DAIRY|-80.562829|80.562830632871794|129|1
35.006282|86fccda3f64ef894581516e8cb5ac045e25901dc|3.69|2015-01-28 17:19:00|80.562862110758871|3|7518500003|60|35.040504021150888|0|21|1033|-80.64817|163|35.04711|HAMBURGER|1.1|7|MARTIN'S POTATO SANDWICH ROLLS|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00075185000039|BUNS/ROLLS|COMMERCIAL BAKERY|-80.562829|80.562830632871794|129|1
35.006282|10f2a4044b1edce333cd03cc83bebc8953c14142|2.99|2015-02-01 16:34:00|80.562862110758871|3|7565604301|60|35.040503999375318|0|21|6821|-80.62331|1580|35.140781|J HOOK LAMI PROGRAM|0.0|18|WRESTLER STICKY FIGHTER|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00075656043015|J-HOOK|GM|-80.562829|80.562876170729723|39|1
35.006282|ea0f8d9c4fc2cab373775d88fe6f1cef1bd3fae9|4.99|2015-01-31 14:38:00|1.4091206135396188|3|7403006610|60|0.6109748797816256|0|47|332|-80.562829|52|35.006282|STRING/SNACK|1.99|3|SORRENTO CHEDDAR STICKSTERS|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|0.61242566243833529|00074030069207|CHEESE|DAIRY|-80.562829|1.4060866207711706|60|1
35.006282|5cab135be7cb251fbd38bba7b9cbc00f2a8459ed|9.99|2015-03-07 20:07:00|80.562862110758871|3|8143431530|60|35.040504021150888|0|21|9962|-80.64817|887|35.04711|NFS-PREM-SAUV/FUME'BLANC|0.0|13|CB-NOBILO SAUVIGNON BLANC|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00081434315304|SUPER PREMIUM ($11-$14.99)|WINE|-80.562829|80.562830632871794|129|1
35.006282|86475bd344d52abadb381008e8fe73cc0b72e19a|7.98|2014-10-21 13:19:00|80.562862110758871|3|7464100992|60|35.040504021150888|0|21|562|-80.64817|64|35.04711|FRESH CUT FRUIT|0.0|4|RED APPLE SLICES 14OZ|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00074641009920|FRESH PRODUCE|PRODUCE|-80.562829|80.562830632871794|129|2
35.006282|7424455d66b767d848f598ad7c943dade22a33c1|11.99|2014-10-30 19:45:00|80.562862110758871|3|8143431530|60|35.040503999375318|0|21|9962|-80.62331|887|35.140781|NFS-PREM-SAUV/FUME'BLANC|0.0|13|CB-NOBILO SAUVIGNON BLANC|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00081434315304|SUPER PREMIUM ($11-$14.99)|WINE|-80.562829|80.562876170729723|39|1
35.006282|18cb88dd520956d64f9f8b7a0c7cb5eb6a01f2b9|15.99|2014-12-06 19:25:00|80.562862110758871|3|8769200033|60|35.040504015557424|0|21|463|-80.709466|84|35.124987|HARD CIDER|0.0|16|ANGRY ORCHARD CRISP CIDER 12PK|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00087692000334|SPECIALTY|BEER|-80.562829|80.562852948591427|157|1
35.006282|58075d670dcbbe6b3c0e63a3fab6841c148cdef3|3.29|2014-09-30 20:15:00|80.562862110758871|3|4157009460|60|35.040503999375318|0|21|1148|-80.62331|21|35.140781|ALMONDS|0.0|1|BLUE DIAM ALM CARML MACCHIATO|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00041570094600|NUTS|G1 GROCERY|-80.562829|80.562876170729723|39|1
35.006282|74a85fc6536f0f9bfe321b0b034e8f6a3209748a|3.29|2014-12-19 19:14:00|80.562862110758871|3|4157009460|60|35.040504009909071|0|21|1148|-80.654118|21|35.123768|ALMONDS|1.0|1|BLUE DIAM ALM CARML MACCHIATO|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00041570094600|NUTS|G1 GROCERY|-80.562829|80.562862911720046|473|1
35.006282|fec13104060760871d000e950e924d06bffee388|3.29|2014-11-28 17:19:00|80.562862110758871|3|4157009460|60|35.040504021150888|0|21|1148|-80.64817|21|35.04711|ALMONDS|0.0|1|BLUE DIAM ALM CARML MACCHIATO|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00041570094600|NUTS|G1 GROCERY|-80.562829|80.562830632871794|129|1
35.006282|ceb4d437a4b2d5d1f9cb02372592df26649ed544|3.63|2015-02-15 21:01:00|80.562862110758871|3||60|35.040504021150888|0|21|523|-80.64817|64|35.04711|FRESH POTATOES|0.0|4|COO SWEET POTATOES, BULK|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00204091000004|FRESH PRODUCE|PRODUCE|-80.562829|80.562830632871794|129|1
35.006282|5100d3ee3f8aa72aeb7712d6563e2a48290e55ff|4.99|2014-11-01 22:29:00|80.562862110758871|3|2531711100|60|35.040503999375318|0|21|845|-80.62331|100|35.140781|NATURAL/ORGANIC BACON|1.49|19|APPLEGATE GOOD MORNING BACON|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00025317111003|BACON|CASE READY MEATS|-80.562829|80.562876170729723|39|1
35.006282|74ce19ea0bf7c59f75161a965f8a59e2e80f1faa|5.19|2015-02-25 19:37:00|80.562862110758871|3|74236526435|60|35.040504015557424|0|21|345|-80.709466|57|35.124987|ORGANIC MILK|0.0|3|HORIZON WHOLE  DHA|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00742365264474|MILK|DAIRY|-80.562829|80.562852948591427|157|1
35.006282|223fb17deeb22f38ad39fcc3bc76486f234e71c6|4.69|2014-10-19 19:18:00|80.562862110758871|3|7468309950|60|35.040504021150888|0|21|1220|-80.64817|275|35.04711|PASTA SC PREMIUM|1.7|1|EMERIL PASTA SC MARINARA|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00074683099460|PASTA SAUCES|G1 GROCERY|-80.562829|80.562830632871794|129|1
35.006282|2bb09d21031e924bd54d164047ef6805724bf9b8|3.49|2014-12-26 17:15:00|80.562862110758871|3|7203676172|60|35.040503999375318|0|21|92|-80.62331|13|35.140781|REMAINING CRACKERS|1.49|1|HTT VEGETABLE SNACK CRACKER|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00072036761705|CRACKERS|G1 GROCERY|-80.562829|80.562876170729723|39|1
35.006282|a261eb210adaf65d51db75475422ebe17e8a110e|4.8|2015-02-18 21:22:00|80.562862110758871|3|3663202717|60|35.040504021150888|0|21|685|-80.64817|61|35.04711|GREEK|0.0|3|DANNON OIKOS STRAWBERRY TRAD|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00036632032188|YOGURT|DAIRY|-80.562829|80.562830632871794|129|4
35.006282|cdad22814c90af15a554ef92a36e110043fe19e2|2.4|2015-02-08 15:22:00|80.562862110758871|3|3663202717|60|35.040503999375318|0|21|685|-80.62331|61|35.140781|GREEK|0.0|3|DANNON OIKOS STRAWBERRY TRAD|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00036632032188|YOGURT|DAIRY|-80.562829|80.562876170729723|39|2
35.006282|433a5ea4f5eefb527348285452382610eba68684|5.49|2015-01-02 22:00:00|80.562862110758871|3|2301290132|60|35.040504021150888|0|21|1477|-80.64817|485|35.04711|SUSHI HYBRID|0.0|6|SPICY CALIFORNIA ROLL SP|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00023012901325|SUSHI|DELI|-80.562829|80.562830632871794|129|1
35.006282|2736e848d66c39870455fd01af32b2127cc43d42|7.49|2015-01-07 20:53:00|80.562862110758871|3|87240800453|60|35.040503999375318|0|21|1226|-80.62331|107|35.140781|HEAT & EAT ENTREES|0.0|19|MAMA MANCINI'S BEEF MEATBALLS|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00872408004535|HEAT & EAT|CASE READY MEATS|-80.562829|80.562876170729723|39|1
35.006282|7ab88cbfca426afbf57dbbdc5e2b7bed183f105d|11.99|2014-09-10 20:26:00|80.562862110758871|3|2301286481|60|35.040504021150888|0|21|1477|-80.64817|485|35.04711|SUSHI HYBRID|0.0|6|"CHEF SAMPLER ""A"""|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00023012864811|SUSHI|DELI|-80.562829|80.562830632871794|129|1
35.006282|e8510a80045d4609448cb652dbc5dbdc668b5de7|11.99|2014-09-19 21:38:00|80.562862110758871|3|2301286481|60|35.040503999375318|0|21|1477|-80.62331|485|35.140781|SUSHI HYBRID|0.0|6|"CHEF SAMPLER ""A"""|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00023012864811|SUSHI|DELI|-80.562829|80.562876170729723|39|1
35.006282|04d114767f39bb6cf4dc1510892c6aed4af571a0|3.99|2014-10-23 08:46:00|1.4091206135396188|3|87606300201|60|0.6109748797816256|0|47|97|-80.562829|8|35.006282|ENERGY DRINKS|0.5|23|MUSCLE MILK CHOCOLATE|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|0.61242566243833529|00876063002011|CARBONATED BEVERAGES|BEVERAGE|-80.562829|1.4060866207711706|60|1
35.006282|f4aeaa45a162bc0959db2144c7926547e83506a8|3.99|2014-12-21 19:12:00|80.562862110758871|3|4470009219|60|35.040503999375318|0|21|498|-80.62331|111|35.140781|PICKLES & SAUERKRAUT|0.99|19|CLAUSSEN MINI PICKLES|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00044700091920|MISC. PACKAGED MEATS|CASE READY MEATS|-80.562829|80.562876170729723|39|1
35.006282|9f02b69329bb2a9d37ee39d54fac2321bcdf1115|6.69|2014-09-18 20:28:00|80.562862110758871|3|4138309070|60|35.040503999375318|0|21|1263|-80.62331|57|35.140781|GOOD FOR YOU MILK|0.7|3|100 LACTAID WHOLE MILK|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00041383090738|MILK|DAIRY|-80.562829|80.562876170729723|39|1
35.006282|a737d2b0d7e3e2eb0751692b665090447554b2e4|7.38|2014-12-24 13:07:00|80.562862110758871|3|2016922150|60|35.040504021150888|0|21|494|-80.64817|107|35.04711|HEAT & EAT SIDES|1.19|19|SIMPLY MASHED POTATOES|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00020169221504|HEAT & EAT|CASE READY MEATS|-80.562829|80.562830632871794|129|2
35.006282|658fe6af32ad380d9b5b8f2e687b6dd233f8297c|6.49|2014-10-09 20:37:00|80.562862110758871|3|2301290139|60|35.040503999375318|0|21|1477|-80.62331|485|35.140781|SUSHI HYBRID|0.0|6|SPICY SALMON ROLL SP|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00023012901394|SUSHI|DELI|-80.562829|80.562876170729723|39|1
35.006282|21340b731ad254a48339d06583b0edd9b8c4e214|3.1|2014-10-26 16:45:00|80.562862110758871|3|3700000445|60|35.040503999375318|0|21|725|-80.62331|66|35.140781|NFS-DISHWASHING LIQUID|0.55|1|DAWN LIQ DISH ORIGINAL 9OZ|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00037000004455|DETERGENTS|G1 GROCERY|-80.562829|80.562876170729723|39|2
35.006282|74609fd45d09cf8f94b148f617815179698ad146|9.38|2014-09-26 18:09:00|1.4091206135396188|3|81829001282|60|0.6109748797816256|0|47|685|-80.562829|61|35.006282|GREEK|1.4|3|CHOBANI KEY LIME BLEND 2% 4PK|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|0.61242566243833529|00818290012753|YOGURT|DAIRY|-80.562829|1.4060866207711706|60|2
35.006282|b7f26fc0198f2dd88b356109fedda2100337d6a4|6.27|2015-01-14 20:34:00|80.562862110758871|3|7203676359|60|35.040503999375318|0|21|345|-80.62331|57|35.140781|ORGANIC MILK|0.0|3|HTO ORGANIC 2% MILK GAL|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00072036763600|MILK|DAIRY|-80.562829|80.562876170729723|39|1
35.006282|384b184b5b20190a877fc4e7e77ab29476b3bb77|1.36|2014-10-15 17:22:00|80.562862110758871|3||60|35.040503999375318|0|21|502|-80.62331|64|35.140781|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00204011000008|FRESH PRODUCE|PRODUCE|-80.562829|80.562876170729723|39|1
35.006282|6adfa97f0e49721e0ad5a6a6045f02f7845441ed|12.99|2015-01-30 20:30:00|80.562862110758871|3|7231123012|60|35.040503999375318|0|21|459|-80.62331|83|35.140781|IMPORT BEER|0.0|16|DOS EQUIS SP LG 12PK 12OZ BTL|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00072311230124|IMPORT BEER|BEER|-80.562829|80.562876170729723|39|1
35.006282|febb3a4b1bafdd1536157bcb3bae0039ea1583f7|7.35|2014-11-12 20:44:00|80.562862110758871|3|4470002268|60|35.040503999375318|0|21|358|-80.62331|100|35.140781|REGULAR BACON|3.68|19|OSCAR MAYER THICK SLIC BACON|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00044700019900|BACON|CASE READY MEATS|-80.562829|80.562876170729723|39|1
35.006282|445e53a959ca07b2f248583e1c383025e2ed1993|1.36|2014-11-05 17:59:00|1.4091206135396188|3||60|0.6109748797816256|0|47|502|-80.562829|64|35.006282|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|0.61242566243833529|00204011000008|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|1
35.006282|75c19bd81c3673e7498bda690b0801e0113c0d3f|14.99|2015-02-21 22:05:00|80.562862110758871|3|8378337512|60|35.040504021150888|0|21|458|-80.64817|82|35.04711|CRAFT BEER|0.0|16|SIERRA PALE ALE 12PK BOTTLE|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00083783375121|DOMESTIC BEER|BEER|-80.562829|80.562830632871794|129|1
35.006282|c167bfccd14c55af12ef691d1574a095212ca395|8.99|2014-11-21 19:14:00|80.562862110758871|3|8834510151|60|35.040504015557424|0|21|463|-80.709466|84|35.124987|HARD CIDER|0.0|16|STRONGBOW GOLD CIDER 6PK BTL|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00088345101514|SPECIALTY|BEER|-80.562829|80.562852948591427|157|1
35.006282|7d2dc1d17a73945af5316425d7d72b9df0fdf6ed|8.99|2015-01-23 21:36:00|80.562862110758871|3|8130800043|60|35.040503999375318|0|21|9950|-80.62331|886|35.140781|NFS-PREM-SAUV/FUME'BLANC|0.0|13|CB-CUPCAKE SAUV BLANC|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00081308000435|PREMIUM ($8-$10.99)|WINE|-80.562829|80.562876170729723|39|1
35.006282|aee6f9e3a4ad47cde155f5807f6b6b4b27530952|8.99|2014-11-15 22:28:00|80.562862110758871|3|8858649895|60|35.040504015557424|0|21|9947|-80.709466|886|35.124987|NFS-PREM-CHARDONNAY|0.0|13|CB-COLUMBIA CRST GRN EST CHARD|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00088586498954|PREMIUM ($8-$10.99)|WINE|-80.562829|80.562852948591427|157|1
35.006282|424060d89ef2b13cad62da74cd4efccef17fd089|8.99|2015-02-24 10:38:00|80.562862110758871|3|7080004170|60|35.040504021150888|0|21|1489|-80.64817|100|35.04711|STACK PACK BACON|3.0|19|SMFD APPLEWOOD STACK BACON|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00070800041701|BACON|CASE READY MEATS|-80.562829|80.562830632871794|129|1
35.006282|e755cea9ab8188d37b158b591d1108f5705075a2|3.79|2014-11-04 19:07:00|80.562862110758871|3|4138309010|60|35.040503999375318|0|21|1263|-80.62331|57|35.140781|GOOD FOR YOU MILK|0.0|3|LACTAID 100 WHOLE MILK|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00041383090363|MILK|DAIRY|-80.562829|80.562876170729723|39|1
35.006282|f9abb1b000dcc1b29a8eeb817ac32f9196a9d8a4|4.29|2015-01-24 18:07:00|80.562862110758871|3|2840006399|60|35.040503999375318|0|21|204|-80.62331|31|35.140781|TORTILLA CHIPS|1.29|1|TOSTITOS SCOOPS 10 OZ|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00028400064088|SNACKS|G1 GROCERY|-80.562829|80.562876170729723|39|1
35.006282|a9608078e812d2f8edfed7248c53779a69ea9a18|14.99|2014-11-08 22:56:00|80.562862110758871|3|79603061493|60|35.040504017639627|0|21|458|-80.770346|82|35.052812|CRAFT BEER|0.0|16|KONA VARIETY 12PK BOTTLES|5c271f493833580d74445561ced557aa59f11240|2.3646590201096993|35.054042368968126|00796030614934|DOMESTIC BEER|BEER|-80.562829|80.562848000659855|40|1
34.977331|99880b7de23632938a69cf924af810acbbc357a1|1.0|2014-12-09 14:39:00|1.41290891556208|4|78352054321|149|0.6104695895098807|0|33|8598|-81.027334|1792|34.977331|NEWSPAPERS|0.0|18|DAILY  CHARLOTTE OBSERVER|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00783520543218|NEWSPAPERS|GM|-81.027334|1.4141937624131469|149|1
34.977331|a80c00329f9fcac6f2181053acfe6da5413460b4|1.0|2015-03-06 18:06:00|1.41290891556208|4|78352054321|149|0.6104695895098807|0|33|8598|-81.027334|1792|34.977331|NEWSPAPERS|0.0|18|DAILY  CHARLOTTE OBSERVER|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00783520543218|NEWSPAPERS|GM|-81.027334|1.4141937624131469|149|1
34.977331|8fe50e885c3131db1e825a2b89492683b7188803|1.0|2015-02-20 17:56:00|1.41290891556208|4|78352054321|149|0.6104695895098807|0|33|8598|-81.027334|1792|34.977331|NEWSPAPERS|0.0|18|DAILY  CHARLOTTE OBSERVER|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00783520543218|NEWSPAPERS|GM|-81.027334|1.4141937624131469|149|1
34.977331|1e49e8387d1058f9d9fb6ea13e99f19371a782bf|2.59|2015-01-06 00:09:00|1.41290891556208|4|79271600032|149|0.6104695895098807|0|33|398|-81.027334|69|34.977331|NFS-BATHROOM CLEANERS|0.0|1|CLEAN SHOWER DAILY SHOWER CLEA|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00792716000329|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|ddef2cde2749403c5ecd89ca72ee7691f4f21257|2.29|2014-09-16 16:59:00|1.41290891556208|4|7203695175|149|0.6104695895098807|0|33|1607|-81.027334|371|34.977331|FROZEN DOUGH (BREAD)|0.0|14|FRESH LRG FRENCH BREAD|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00072036951755|BREAD|BAKERY|-81.027334|1.4141937624131469|149|1
34.977331|a1c7b25b57b386eb0c8d32093ba3ac9d46a7f052|7.99|2014-12-19 00:06:00|1.41290891556208|4|84323700813|149|0.6104695895098807|0|33|670|-81.027334|146|34.977331|CRAB PACKAGED|0.0|12|CHICKEN OF THE SEA 8OZ  CLAW|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00843237008131|CRAB|SEAFOOD|-81.027334|1.4141937624131469|149|1
34.977331|d513492210b932232d14ce32c2cb8a9d56fc2bd6|4.99|2015-02-28 18:27:00|1.41290891556208|4|87604500400|149|0.6104695895098807|0|33|68|-81.027334|11|34.977331|BARBECUE SAUCES|0.0|1|GUY FIERI BBQ SC CAROLINA # 6|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00876045004002|CONDIMENTS|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|592ffa88e1b60fb029fef2467d8d1176bc0659ce|5.75|2014-10-07 13:21:00|1.41290891556208|4|20807400000|149|0.6104695895098807|0|33|648|-81.027334|154|34.977331|FISH FLTS/STK FARM RAISD|0.0|12|FRESH CATFISH FILLETS|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00208074000005|FISH FILLETS/STEAKS|SEAFOOD|-81.027334|1.4141937624131469|149|1
34.977331|ce978d6f2651ecd3aa5fcc574315e9e336ac0b9f|1.34|2014-10-13 17:10:00|1.41290891556208|4|7203627087|149|0.6104695895098807|0|33|158|-81.027334|24|34.977331|NFS-DOG FOOD-WET|0.0|1|HT YOURPET GRAVY LONDON GRILL|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00072036310439|PET FOOD/SUPPLIES|G1 GROCERY|-81.027334|1.4141937624131469|149|2
34.977331|9858166c2ed937b0e73742daa6fb5b68a2d4476e|2.85|2014-09-15 14:07:00|1.41290891556208|4|1380010321|149|0.6104695895098807|0|33|1279|-81.027334|48|34.977331|SINGLE SERVE FLAVOR|0.0|5|STOUF MAC&CHEESE W/BROCC|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00013800447920|FROZEN MEALS|FROZEN|-81.027334|1.4141937624131469|149|1
34.977331|47582d8b04921062c4881597c8e72770f1d1982d|22.79|2015-02-03 18:07:00|1.41290891556208|4|20220200000|149|0.6104695895098807|0|33|299|-81.027334|49|34.977331|ANGUS BEEF|5.7|2|ANGUS BEEF FILET MIGNON CUSTOM|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00202209000007|BEEF|MEAT|-81.027334|1.4141937624131469|149|1
34.977331|3c6f92cdb0a1d5e62b6343545e2366bd1e5cab82|0.37|2014-09-23 15:28:00|1.41290891556208|4||149|0.6104695895098807|0|33|526|-81.027334|64|34.977331|FRESH MUSHROOMS|0.0|4|USA WHITE MUSHROOMS, BULK|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00204085000003|FRESH PRODUCE|PRODUCE|-81.027334|1.4141937624131469|149|1
34.977331|ddd70ad3af4423bb9c001acf811e9abaaf1f5e07|1.79|2014-11-03 15:48:00|1.41290891556208|4|5100001047|149|0.6104695895098807|0|33|212|-81.027334|33|34.977331|CONDENSED SOUP|0.79|1|CAMP COND BROCCOLLI CHEESE|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00051000013477|SOUP|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|cef575705184820ec41430bf2ac7205814d07c7a|3.49|2015-03-08 15:53:00|1.41290891556208|4|2840008294|149|0.6104695895098807|0|33|201|-81.027334|31|34.977331|POTATO CHIPS|0.49|1|LAYS KETTLE REGULAR|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00028400082945|SNACKS|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|06c0d6c45dbcc6cb315cc9e326f9dd7e6cfe8042|3.49|2014-12-28 17:24:00|1.41290891556208|4|2840008294|149|0.6104695895098807|0|33|201|-81.027334|31|34.977331|POTATO CHIPS|0.99|1|LAYS KETTLE REGULAR|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00028400082945|SNACKS|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|03436ff69e64713d65b68309a269494484f7270d|3.49|2014-09-29 15:40:00|1.41290891556208|4|2840008294|149|0.6104695895098807|0|33|201|-81.027334|31|34.977331|POTATO CHIPS|0.99|1|LAYS KETTLE REGULAR|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00028400082945|SNACKS|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|8a4c8ddda86b5f963ece1af7f4b8eb6171d6607c|7.79|2014-09-29 15:41:00|1.41290891556208|4|20943400000|149|0.6104695895098807|0|33|883|-81.027334|145|34.977331|SHRIMP FARM RAISED|4.16|12|31/40 CT EZ PEEL WHITE SHRIMP|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00209434000000|SHRIMP|SEAFOOD|-81.027334|1.4141937624131469|149|1
34.977331|e6e4c2a546253a692bb18a8465460d850b2580f6|3.99|2014-10-18 23:45:00|1.41290891556208|4|4157005982|149|0.6104695895098807|0|33|1148|-81.027334|21|34.977331|ALMONDS|0.99|1|B D ALMONDS B JALAPENO SMK HSE|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00041570052327|NUTS|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|8ffc54bbe0c79799f41a6e176bb739e19c984f9b|3.99|2015-02-25 18:49:00|1.41290891556208|4|4157005982|149|0.6104695895098807|0|33|1148|-81.027334|21|34.977331|ALMONDS|0.0|1|B D ALMONDS B JALAPENO SMK HSE|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00041570052327|NUTS|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|e1644909138416d24bb008d01edd7c2eb28a224e|3.69|2014-11-25 14:46:00|1.41290891556208|4|4178000159|149|0.6104695895098807|0|33|201|-81.027334|31|34.977331|POTATO CHIPS|1.19|1|UTZ CLASSICS B B Q CHIPS|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00041780001795|SNACKS|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|3a238a26bd22925e227753c5772f178029123fc2|3.59|2015-02-26 20:29:00|1.41290891556208|4|4116400022|149|0.6104695895098807|0|33|1469|-81.027334|278|34.977331|REGULAR CUT FRIES|0.0|5|MRS.TLOADED BAKD POTA PIEROGIE|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00041164000482|FROZEN POTATO|FROZEN|-81.027334|1.4141937624131469|149|1
34.977331|cc936fb9a1387448eb7e6789c4ea95a31ee69482|1.79|2015-02-04 16:39:00|1.41290891556208|4|7342000006|149|0.6104695895098807|0|33|322|-81.027334|53|34.977331|SOUR CREAM|0.0|3|DAISY LIGHT SOUR CREAM|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00073420000059|CULTURES|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|e9d246d5c7d1f10f415c3566a12ea1697ec0e6b5|1.98|2014-11-11 14:04:00|1.41290891556208|4|2310001004|149|0.6104695895098807|0|33|158|-81.027334|24|34.977331|NFS-DOG FOOD-WET|0.58|1|PEDIGREE CHOICE CUTS - BEEF|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00023100015279|PET FOOD/SUPPLIES|G1 GROCERY|-81.027334|1.4141937624131469|149|2
34.977331|9c9d085c55f4ff713fb6767759a62e06e4038f56|1.98|2015-01-13 14:15:00|1.41290891556208|4|2310001004|149|0.6104695895098807|0|33|158|-81.027334|24|34.977331|NFS-DOG FOOD-WET|0.38|1|PEDIGREE CHOICE CUTS - BEEF|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00023100015279|PET FOOD/SUPPLIES|G1 GROCERY|-81.027334|1.4141937624131469|149|2
34.977331|e55c40cd69f007bd863c55f7eeab75cf59569368|6.99|2015-01-20 15:53:00|1.41290891556208|4|2301200114|149|0.6104695895098807|0|33|1475|-81.027334|485|34.977331|SUSHI CLASSIC|0.0|6|FULL MOON COMBO|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00023012001148|SUSHI|DELI|-81.027334|1.4141937624131469|149|1
34.977331|9e0465b37ab6ec712ccefb450595b8e980d64543|3.97|2015-02-15 18:55:00|1.41290891556208|4|7203658034|149|0.6104695895098807|0|33|358|-81.027334|100|34.977331|REGULAR BACON|0.0|19|HT REGULAR SLICED BACON|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00072036580344|BACON|CASE READY MEATS|-81.027334|1.4141937624131469|149|1
34.977331|3347259e3231781b855f5a9efaa481425a0656f5|1.98|2015-01-28 16:05:00|1.41290891556208|4|2310001004|149|0.6104695895098807|0|33|158|-81.027334|24|34.977331|NFS-DOG FOOD-WET|0.38|1|PEDIGREE CHOICE CUT BEEF/LIVER|5c4b409524e319a4b23e1d3e4fdd9c11af2e358f|1.8650323203231711|0.61055446569467375|00023100015330|PET FOOD/SUPPLIES|G1 GROCERY|-81.027334|1.4141937624131469|149|2
35.17739|a2d56771598f186e0ac51166dde5b0810f5a4d59|6.79|2015-01-02 13:12:00|1.4094857484078087|3|1200080994|208|0.613961277758128|0|26|54|-80.80146|8|35.17739|DIET|6.79|23|DT PEPSI FRIDGEMATE|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00012000809958|CARBONATED BEVERAGES|BEVERAGE|-80.80146|1.4102515174184975|208|1
35.17739|e84bf3387f132e360b0322306bc22410268dffeb|19.21|2014-09-18 22:37:00|1.4094857484078087|3|20895300000|208|0.613961277758128|0|26|977|-80.80146|201|35.17739|FRESH HT CHICKEN|4.52|2|HT FRESH BNLS CHICKEN BREAST|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00208953000003|POULTRY|MEAT|-80.80146|1.4102515174184975|208|2
35.17739|8c03090a4aa317128a12a1244b19d1bc2159d778|2.49|2015-02-19 19:53:00|1.4094857484078087|3|7203688048|208|0.613961277758128|0|26|526|-80.80146|64|35.17739|FRESH MUSHROOMS|0.2|4|HT SLICED BABY BELLAS|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00072036880482|FRESH PRODUCE|PRODUCE|-80.80146|1.4102515174184975|208|1
35.17739|30f82b947b4fefc360aac5428005790d36f6b32a|1.69|2015-02-25 18:32:00|1.4094857484078087|3|7203688003|208|0.613961277758128|0|26|527|-80.80146|64|35.17739|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00072036880031|FRESH PRODUCE|PRODUCE|-80.80146|1.4102515174184975|208|1
35.17739|80ada84c1e4618b080da1d1ec9e57d15135e9d0e|2.78|2015-01-02 13:07:00|1.4094857484078087|3|7203624015|208|0.613961277758128|0|26|149|-80.80146|23|35.17739|WHSE PASTA CORE|0.7|1|HT PASTA ELBOW MAC 16|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00072036240149|PASTA|G1 GROCERY|-80.80146|1.4102515174184975|208|2
35.17739|b9e2cebbab8e95c2cefdc06c17a0c00a23243a40|1.49|2014-12-04 19:43:00|1.4094857484078087|3|7203611080|208|0.613961277758128|0|26|977|-80.80146|201|35.17739|FRESH HT CHICKEN|0.0|2|HT CHICKEN LIVERS|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00072036110800|POULTRY|MEAT|-80.80146|1.4102515174184975|208|1
35.17739|2a86a723816c220cf2429a94fc51fdbe770dd4c4|2.67|2014-10-19 15:26:00|1.4094857484078087|3|7203653120|208|0.613961277758128|0|26|1273|-80.80146|50|35.17739|BAG VEG NON STEAM|0.0|5|HT CHOPPED ONIONS|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00072036531209|VEGETABLES-FROZEN|FROZEN|-80.80146|1.4102515174184975|208|2
35.17739|54dbcb1913beee7e42642c5ed819038b522df3a1|6.9|2014-12-14 17:28:00|1.4094857484078087|3|7203663995|208|0.613961277758128|0|26|342|-80.80146|57|35.17739|FRESH MILK|0.0|3|HARRIS TEETER 1% MILK|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00072036631275|MILK|DAIRY|-80.80146|1.4102515174184975|208|2
35.17739|a01f3e2c5033907eaf5397912daf2e1dc4cd02fb|3.99|2014-10-13 19:31:00|1.4094857484078087|3|7203663995|208|0.613961277758128|0|26|342|-80.80146|57|35.17739|FRESH MILK|0.0|3|HARRIS TEETER 1% MILK|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00072036631275|MILK|DAIRY|-80.80146|1.4102515174184975|208|1
35.17739|1c0904df7719799b4e40afe7ed0fe7c2191ffbcd|3.99|2014-12-28 07:46:00|1.4094857484078087|3|7203663995|208|0.613961277758128|0|26|342|-80.80146|57|35.17739|FRESH MILK|0.0|3|HARRIS TEETER 1% MILK|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00072036631275|MILK|DAIRY|-80.80146|1.4102515174184975|208|1
35.17739|609790489d96fb04664cecaafee1fe87f7901e95|6.98|2014-11-07 15:42:00|1.4094857484078087|3|7203663995|208|0.613961277758128|0|26|342|-80.80146|57|35.17739|FRESH MILK|0.0|3|HARRIS TEETER 1% MILK|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00072036631275|MILK|DAIRY|-80.80146|1.4102515174184975|208|2
35.17739|be26f8c07cc25c07bd130dd185f561dcb842e9df|11.32|2014-11-20 20:46:00|1.4094857484078087|3|1707710232|208|0.613961277758128|0|26|1455|-80.80146|61|35.17739|DRINKABLE YOGURT|1.78|3|LIFEWAY KEFIR PLAIN|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00017077102322|YOGURT|DAIRY|-80.80146|1.4102515174184975|208|4
35.17739|bf1105102adaf8b2ead3c5a86cd7fd3830b98802|7.78|2014-11-14 14:15:00|1.4094857484078087|3|1707710232|208|0.613961277758128|0|26|1455|-80.80146|61|35.17739|DRINKABLE YOGURT|2.12|3|LIFEWAY KEFIR PLAIN|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00017077102322|YOGURT|DAIRY|-80.80146|1.4102515174184975|208|2
35.17739|61f56a5677e2469acc450e6dff97d62136381c1b|15.56|2015-01-24 12:12:00|1.4094857484078087|3|1707710232|208|0.613961277758128|0|26|1455|-80.80146|61|35.17739|DRINKABLE YOGURT|2.12|3|LIFEWAY KEFIR PLAIN|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00017077102322|YOGURT|DAIRY|-80.80146|1.4102515174184975|208|4
35.17739|c4f21a14981b1205514dfa504f58f6470110ae25|11.67|2015-02-23 19:04:00|1.4094857484078087|3|1707710232|208|0.613961277758128|0|26|1455|-80.80146|61|35.17739|DRINKABLE YOGURT|6.36|3|LIFEWAY KEFIR PLAIN|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00017077102322|YOGURT|DAIRY|-80.80146|1.4102515174184975|208|3
35.17739|55eb87dbbcaae753701a9514423cf528d153d5ef|4.9|2014-09-12 13:24:00|1.4094857484078087|3|1450000253|208|0.613961277758128|0|26|1273|-80.80146|50|35.17739|BAG VEG NON STEAM|1.22|5|BE PEPPER STIR FRY|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00014500505637|VEGETABLES-FROZEN|FROZEN|-80.80146|1.4102515174184975|208|2
35.17739|986e117fc18db455beeea633faa9775ae1b4821f|11.67|2014-12-07 18:47:00|1.4094857484078087|3|1707710232|208|0.613961277758128|0|26|1455|-80.80146|61|35.17739|DRINKABLE YOGURT|6.36|3|LIFEWAY KEFIR PLAIN|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00017077102322|YOGURT|DAIRY|-80.80146|1.4102515174184975|208|3
35.17739|f2d1acb0ab430ef10c4c275a1edebe389dae4640|6.98|2014-10-30 17:43:00|1.4094857484078087|3|4812127620|208|0.613961277758128|0|26|1037|-80.80146|164|35.17739|ENGLISH MUFFINS|1.75|7|THOMAS LITE MULTIGRAIN EM PP|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00048121276201|BREAKFAST|COMMERCIAL BAKERY|-80.80146|1.4102515174184975|208|2
35.17739|bd49bc60ee742470039f5d47598846b79e83cb2f|3.85|2015-02-13 15:14:00|1.4094857484078087|3|4812127620|208|0.613961277758128|0|26|1037|-80.80146|164|35.17739|ENGLISH MUFFINS|1.93|7|THOMAS LITE MULTIGRAIN EM PP|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00048121276201|BREAKFAST|COMMERCIAL BAKERY|-80.80146|1.4102515174184975|208|1
35.17739|6ce66ab3ceaa601d39c8b8a92199e7cb3708efc4|0.99|2014-12-22 10:19:00|1.4094857484078087|3||208|0.613961277758128|0|26|540|-80.80146|64|35.17739|FRESH CELERY|0.0|4|COO CELERY (RPC) 24'S|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00204070000001|FRESH PRODUCE|PRODUCE|-80.80146|1.4102515174184975|208|1
35.17739|1390ccf3f6a5ba274bce9700a5649d8625ed50c3|1.29|2014-09-25 20:18:00|1.4094857484078087|3||208|0.613961277758128|0|26|505|-80.80146|64|35.17739|FRESH SOFT FRUIT|0.09|4|WHITE NECTARINES PLU#|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00233035000008|FRESH PRODUCE|PRODUCE|-80.80146|1.4102515174184975|208|1
35.17739|b5458175ed6a21d5f79d42636495c8b96ebbd75a|3.99|2015-03-09 15:51:00|1.4094857484078087|3|3338310366|208|0.613961277758128|0|26|509|-80.80146|64|35.17739|FRESH CITRUS-REMAINING|0.99|4|MINNEOLA TANGELO 3LB|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00605049366812|FRESH PRODUCE|PRODUCE|-80.80146|1.4102515174184975|208|1
35.17739|21b22510619924a4cb3e57d9d7ffb765023e0cad|3.98|2014-09-23 14:19:00|1.4094857484078087|3|7203678045|208|0.613961277758128|0|26|151|-80.80146|23|35.17739|DSD PASTA CORE|1.48|1|HT TRADER WW PASTA CAPELLINI|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00072036780485|PASTA|G1 GROCERY|-80.80146|1.4102515174184975|208|2
35.17739|9dca79c16d6b166ed3ac415a3f55af8d9e89697e|0.45|2015-01-30 09:03:00|1.4094857484078087|3||208|0.613961277758128|0|26|522|-80.80146|64|35.17739|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00204664000004|FRESH PRODUCE|PRODUCE|-80.80146|1.4102515174184975|208|1
35.17739|0ccba79126235991c32ee65bb6c6b60f020ff2de|1.25|2015-01-17 16:57:00|1.4094857484078087|3||208|0.613961277758128|0|26|522|-80.80146|64|35.17739|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00204664000004|FRESH PRODUCE|PRODUCE|-80.80146|1.4102515174184975|208|1
35.17739|cda5144e875864775f237c2c10433a55f9df4561|3.99|2015-02-06 14:20:00|1.4094857484078087|3|7127923100|208|0.613961277758128|0|26|555|-80.80146|64|35.17739|PACKAGED SALADS|0.99|4|F.E. BABY SPRING SALAD MIX|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00071279231006|FRESH PRODUCE|PRODUCE|-80.80146|1.4102515174184975|208|1
35.17739|305834ae731f6870d97061b341fce05159779696|2.19|2015-01-01 16:17:00|1.4094857484078087|3|4900005010|208|0.613961277758128|0|26|54|-80.80146|8|35.17739|DIET|0.2|23|COKE ZERO 2 LITER|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00049000050141|CARBONATED BEVERAGES|BEVERAGE|-80.80146|1.4102515174184975|208|1
35.17739|04f0a62d1f29292da3ecb77d48c2762e6b3ff87f|2.97|2014-10-25 14:35:00|1.4094857484078087|3||208|0.613961277758128|0|26|507|-80.80146|64|35.17739|FRESH ORANGES|0.19|4|NAVEL ORANGE, FL XL|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00204385000000|FRESH PRODUCE|PRODUCE|-80.80146|1.4102515174184975|208|3
35.17739|bca27e851593e66d99c35f1ab730d3838fe29e7c|8.0|2015-03-07 14:11:00|1.4094857484078087|3||208|0.613961277758128|0|26|500|-80.80146|64|35.17739|FRESH APPLES|4.02|4|FUJI APPLES|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00204131000001|FRESH PRODUCE|PRODUCE|-80.80146|1.4102515174184975|208|1
35.17739|1e92ad34ab507d64dde8559d1d6d220f333b4041|5.0|2014-11-23 09:01:00|1.4094857484078087|3|7203696869|208|0.613961277758128|0|26|1165|-80.80146|87|35.17739|NFS-FRESH CONSUMER BUNCH|0.0|9|CHRISTMS MIX TULIP BUNCHES  ED|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00072036968692|FLORAL|FLORAL|-80.80146|1.4102515174184975|208|1
35.17739|0d665d53c151ed7c3bfa8c77a5130eb6f4fdc18c|1.99|2015-01-03 16:40:00|1.4094857484078087|3|7203663220|208|0.613961277758128|0|26|330|-80.80146|55|35.17739|EGGS|0.0|3|HT GRADE A    LARGE EGGS|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00072036632203|EGGS FRESH|DAIRY|-80.80146|1.4102515174184975|208|1
35.17739|5b1a81b236db7a69c0e0901d2afd605c57c5faa7|1.99|2015-01-10 17:11:00|1.4094857484078087|3|7203663220|208|0.613961277758128|0|26|330|-80.80146|55|35.17739|EGGS|0.74|3|HT GRADE A    LARGE EGGS|5c7c6959fe97458a36f0655cb5a53f9572a8df06|0.7005874551768377|0.61471665291522548|00072036632203|EGGS FRESH|DAIRY|-80.80146|1.4102515174184975|208|1
34.977331|114b52198ed031e36b1b20743549e79d16f28669|2.0|2014-12-19 22:22:00|1.41290891556208|4|4300095562|149|0.6104695895098807|0|33|209|-81.027334|20|34.977331|POWDERED SOFT DRINKS|0.0|1|K-AID UNSWT LEMON LIME 2 QT|5e1924cce633078c9398c2f04c9148cc1e0d8c38|1.1336624329907317|0.61055446569467375|00043000955444|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-81.027334|1.4141937624131469|149|8
34.977331|c9793235bedb02af909c1f18ae42a5099d777144|1.0|2014-10-30 19:00:00|1.41290891556208|4|4300095562|149|0.6104695895098807|0|33|209|-81.027334|20|34.977331|POWDERED SOFT DRINKS|0.0|1|K-AID UNSWT LEMON LIME 2 QT|5e1924cce633078c9398c2f04c9148cc1e0d8c38|1.1336624329907317|0.61055446569467375|00043000955444|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-81.027334|1.4141937624131469|149|4
34.977331|06483e6a48e6fae25143ffa03f6a1d7b7bcf2c74|13.54|2015-02-05 19:11:00|1.41290891556208|4|20140400000|149|0.6104695895098807|0|33|296|-81.027334|49|34.977331|RANCHER BEEF|0.0|2|BEEF LOIN NY STRIP STEAK BNLS|5e1924cce633078c9398c2f04c9148cc1e0d8c38|1.1336624329907317|0.61055446569467375|00201404000003|BEEF|MEAT|-81.027334|1.4141937624131469|149|2
34.977331|c0ac91abda8bb73c7ea3026acfd1f2cb9c4a43be|4.29|2014-09-24 19:02:00|1.41290891556208|4|2840016014|149|0.6104695895098807|0|33|201|-81.027334|31|34.977331|POTATO CHIPS|0.29|1|LAYS CLASSIC|5e1924cce633078c9398c2f04c9148cc1e0d8c38|1.1336624329907317|0.61055446569467375|00028400160148|SNACKS|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|82ea72b86127102d0863091efd8c5a60277b64a9|4.29|2014-12-16 18:59:00|1.41290891556208|4|2840016014|149|0.6104695895098807|0|33|201|-81.027334|31|34.977331|POTATO CHIPS|0.29|1|LAYS CLASSIC|5e1924cce633078c9398c2f04c9148cc1e0d8c38|1.1336624329907317|0.61055446569467375|00028400160148|SNACKS|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|05cba697faf7e74be009f69e6caf66ea78faf4b6|8.97|2014-12-08 19:17:00|1.41290891556208|4|4610001992|149|0.6104695895098807|0|33|317|-81.027334|52|34.977331|CHUNK AND BAR CHEESE|1.5|3|SARGENTO FIESTA PEPPER JACK|5e1924cce633078c9398c2f04c9148cc1e0d8c38|1.1336624329907317|0.61055446569467375|00046100019931|CHEESE|DAIRY|-81.027334|1.4141937624131469|149|3
34.977331|720491adc6264829433340782ab374f53fc959d5|3.0|2014-10-08 08:14:00|1.41290891556208|4|7203698316|149|0.6104695895098807|0|33|1134|-81.027334|57|34.977331|CARTON MILK|0.0|3|HT CHOCOLATE LOWFAT MILK|5e1924cce633078c9398c2f04c9148cc1e0d8c38|1.1336624329907317|0.61055446569467375|00072036983169|MILK|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|2d7cf7ce1435ea254409e9c94d77bd7303d81b47|3.0|2014-09-19 07:54:00|1.41290891556208|4|7203698316|149|0.6104695895098807|0|33|1134|-81.027334|57|34.977331|CARTON MILK|0.0|3|HT CHOCOLATE LOWFAT MILK|5e1924cce633078c9398c2f04c9148cc1e0d8c38|1.1336624329907317|0.61055446569467375|00072036983169|MILK|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|b7a59752e934d2e4913d8694935d4d80601b79e4|5.37|2015-01-12 19:08:00|1.41290891556208|4|5100002457|149|0.6104695895098807|0|33|212|-81.027334|33|34.977331|CONDENSED SOUP|0.12|1|CAMP COND HMSTL CHICKEN NOODLE|5e1924cce633078c9398c2f04c9148cc1e0d8c38|1.1336624329907317|0.61055446569467375|00051000024572|SOUP|G1 GROCERY|-81.027334|1.4141937624131469|149|3
34.977331|5413bc0d35266fc61de73bd350d87d835a7af3d5|3.49|2014-12-07 15:41:00|1.41290891556208|4|2500004786|149|0.6104695895098807|0|33|335|-81.027334|56|34.977331|ORANGE JUICE-REGRIGERATED|0.5|3|MINUTE MAID PREMIUM OJ|5e1924cce633078c9398c2f04c9148cc1e0d8c38|1.1336624329907317|0.61055446569467375|00025000047862|JUICES & DRINKS-REFRIGERATED|DAIRY|-81.027334|1.4141937624131469|149|1
34.977331|3664c01a40fdb8029c3f8935854082f7c13b709f|1.79|2015-02-07 14:40:00|1.41290891556208|4|4300097940|149|0.6104695895098807|0|33|183|-81.027334|28|34.977331|SALAD DRESSINGS-DRY|0.0|1|GOOD SNS DRY DRS ZESTY ITALIAN|5e1924cce633078c9398c2f04c9148cc1e0d8c38|1.1336624329907317|0.61055446569467375|00043000979037|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-81.027334|1.4141937624131469|149|1
35.116638|fc2117fdfb6840b86873c40e28477188527b40be|6.49|2015-02-28 17:51:00|80.856688219393845|1|5210003038|204|35.132181951641783|0|15|220|-80.85013|34|35.175855|PEPPER|0.0|1|MC WHOLE BLACK PEPPER FAM SIZE|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00052100071282|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.85753|80.85754234393255|218|1
35.116638|a4631820686df531cd569a009dc9e0e81fcd10a1|4.69|2014-10-19 14:31:00|80.856688219393845|1|5210000212|204|35.132181951641783|0|15|1245|-80.85013|34|35.175855|SINGLE SPICES|0.0|1|MC GROUND ALLSPICE|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00052100002125|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.85753|80.85754234393255|218|1
35.116638|65940de17044f487c40d162e18572697d09bf334|0.6|2014-12-24 13:30:00|80.856688219393845|1|7047000100|204|35.132181951641783|0|15|687|-80.85013|61|35.175855|BLENDED|0.0|3|YOPLAIT RASPBERRY YOGURT|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00070470003016|YOGURT|DAIRY|-80.85753|80.85754234393255|218|1
35.116638|b7dceb06ab8fb6b2856a6ee62e986f6686e9dff0|1.2|2015-02-21 12:07:00|80.856688219393845|1|7047000100|204|35.132181951641783|0|15|687|-80.85013|61|35.175855|BLENDED|0.1|3|YOPLAIT RASPBERRY YOGURT|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00070470003016|YOGURT|DAIRY|-80.85753|80.85754234393255|218|2
35.116638|6485688af187e3ba887dc159d70fdad9e1d27a12|1.2|2014-10-25 13:30:00|80.856688219393845|1|7047000100|204|35.132181951641783|0|15|687|-80.85013|61|35.175855|BLENDED|0.0|3|YOPLAIT RASPBERRY YOGURT|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00070470003016|YOGURT|DAIRY|-80.85753|80.85754234393255|218|2
35.116638|f35d9ac5e0e127bfc465681d98cb3cfa248de381|1.89|2014-12-04 12:34:00|80.856688219393845|1|7069002210|204|35.132181951641783|0|15|757|-80.85013|3|35.175855|BAKING NUTS|0.2|1|FISHER ALMONDS SLIVERED|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00070690022101|BAKING SUPPLIES|G1 GROCERY|-80.85753|80.85754234393255|218|1
35.116638|60e9216b3eed7d328358ff25ef0f288eb0914df5|1.2|2015-02-01 16:58:00|80.856688219393845|1|7047000100|204|35.132181951641783|0|15|687|-80.85013|61|35.175855|BLENDED|0.0|3|YOPLAIT RASPBERRY YOGURT|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00070470003016|YOGURT|DAIRY|-80.85753|80.85754234393255|218|2
35.116638|db31b94f11532797c49898d314eac61a0da00cfc|1.6|2014-09-23 20:05:00|80.856688219393845|1|7047000100|204|35.132181951641783|0|15|687|-80.85013|61|35.175855|BLENDED|0.6|3|YOPLAIT RASPBERRY YOGURT|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00070470003016|YOGURT|DAIRY|-80.85753|80.85754234393255|218|2
35.116638|e223983681154ae2a5706ab6fe087c154664585f|1.69|2015-01-29 19:05:00|80.856688219393845|1|4900000044|204|35.132181951641783|0|15|54|-80.85013|8|35.175855|DIET|0.0|23|CB DIET DR PEPPER 20OZ NR|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00078000083408|CARBONATED BEVERAGES|BEVERAGE|-80.85753|80.85754234393255|218|1
35.116638|a8297906d396ec06b09d03ab4401fbb297bb3d66|1.69|2015-01-01 18:29:00|80.856688219393845|1|4900000044|204|35.132181951641783|0|15|54|-80.85013|8|35.175855|DIET|0.0|23|CB DIET DR PEPPER 20OZ NR|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00078000083408|CARBONATED BEVERAGES|BEVERAGE|-80.85753|80.85754234393255|218|1
35.116638|5b9d06aa10d2e037824ffa028331399dd230a5ff|7.78|2014-09-14 17:22:00|80.856688219393845|1|7247000222|204|35.132181951641783|0|15|1641|-80.85013|377|35.175855|PACKAGED DONUTS|0.0|14|K K 6 ORIG GLAZED DONUT  PP|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00072470002228|DONUTS|BAKERY|-80.85753|80.85754234393255|218|2
35.116638|4ea4b49bec55e10ff32ab2ddcdca834ba5d92a2a|1.23|2014-11-11 19:18:00|80.856688219393845|1||204|35.132181951641783|0|15|522|-80.85013|64|35.175855|FRESH TOMATOES|0.0|4|HT VINE RIPE TOMATOES|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00204064000000|FRESH PRODUCE|PRODUCE|-80.85753|80.85754234393255|218|1
35.116638|63d9078504e05a158589331412fe7186d1d0a334|2.37|2014-12-22 19:24:00|80.856688219393845|1||204|35.132181951641783|0|15|501|-80.85013|64|35.175855|FRESH PEARS|0.0|4|BARTLETT PEARS|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00204409000009|FRESH PRODUCE|PRODUCE|-80.85753|80.85754234393255|218|1
35.116638|989dcf538f3880486d0ae2a57722ed1a2c029edb|2.69|2014-11-29 17:45:00|80.856688219393845|1||204|35.132181951641783|0|15|501|-80.85013|64|35.175855|FRESH PEARS|0.0|4|BARTLETT PEARS|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00204409000009|FRESH PRODUCE|PRODUCE|-80.85753|80.85754234393255|218|1
35.116638|f8afba44451674f914ee7da2a6a7a3b121a13c90|4.7|2014-12-13 17:50:00|80.856688219393845|1||204|35.132181951641783|0|15|501|-80.85013|64|35.175855|FRESH PEARS|0.94|4|BARTLETT PEARS|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00204409000009|FRESH PRODUCE|PRODUCE|-80.85753|80.85754234393255|218|2
35.116638|1fed19de7e0ca875f055ac626d3745521b021636|4.16|2014-11-17 19:28:00|80.856688219393845|1||204|35.132181951641783|0|15|501|-80.85013|64|35.175855|FRESH PEARS|0.63|4|BARTLETT PEARS|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00204409000009|FRESH PRODUCE|PRODUCE|-80.85753|80.85754234393255|218|1
35.116638|5ccad832d8775aad2784145653d7b02bd364b43f|2.85|2014-12-05 20:09:00|80.856688219393845|1||204|35.132181951641783|0|15|501|-80.85013|64|35.175855|FRESH PEARS|0.0|4|BARTLETT PEARS|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00204409000009|FRESH PRODUCE|PRODUCE|-80.85753|80.85754234393255|218|1
35.116638|d2d1fde4141c278de5f0e9ddab73d8f1d612118b|4.02|2014-11-05 19:56:00|80.856688219393845|1||204|35.132181951641783|0|15|501|-80.85013|64|35.175855|FRESH PEARS|0.0|4|BARTLETT PEARS|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00204409000009|FRESH PRODUCE|PRODUCE|-80.85753|80.85754234393255|218|1
35.116638|02af4e4682340b842ac6763c6d8fe153ed5903c3|2.49|2015-01-10 17:16:00|80.856688219393845|1||204|35.132181947731389|0|15|561|-80.826724|64|35.195689|FR PROD ORGANIC PRODUCE|0.0|4|ORG HASS AVOCADOS|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00294225000000|FRESH PRODUCE|PRODUCE|-80.85753|80.857548278251102|412|1
35.116638|12acb3ad21cfc9e0ca0b5fc4ce7241d922805710|3.89|2014-11-16 21:41:00|80.856688219393845|1|7684010015|204|35.132181951641783|0|15|275|-80.85013|45|35.175855|SUPER PREMIUM ICE CREAM|0.0|5|BEN & JERRY HALF BAKED|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00076840101320|ICE CREAM|FROZEN|-80.85753|80.85754234393255|218|1
35.116638|c40777229ed4c583e67b7ce954ba3d304e0e2d24|3.89|2014-11-14 23:21:00|80.856688219393845|1|7684010015|204|35.132181951641783|0|15|275|-80.85013|45|35.175855|SUPER PREMIUM ICE CREAM|0.0|5|BEN & JERRY HALF BAKED|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00076840101320|ICE CREAM|FROZEN|-80.85753|80.85754234393255|218|1
35.116638|0376e7a81f15d6483eeb0ae4aa083165dd903f3b|3.89|2014-12-20 16:18:00|80.856688219393845|1|7684010015|204|35.132181951641783|0|15|275|-80.85013|45|35.175855|SUPER PREMIUM ICE CREAM|0.0|5|BEN & JERRY HALF BAKED|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00076840101320|ICE CREAM|FROZEN|-80.85753|80.85754234393255|218|1
35.116638|452a242885a37fe62e1f4647f1608e61ba984cae|3.79|2015-02-07 18:39:00|80.856688219393845|1|7684010015|204|35.132181951641783|0|15|275|-80.85013|45|35.175855|SUPER PREMIUM ICE CREAM|0.29|5|BEN & JERRY HALF BAKED|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00076840101320|ICE CREAM|FROZEN|-80.85753|80.85754234393255|218|1
35.116638|fe6631271c7d20179fb873313bf6acbffe695490|3.89|2014-11-21 19:47:00|80.856688219393845|1|7684010015|204|35.132181951641783|0|15|275|-80.85013|45|35.175855|SUPER PREMIUM ICE CREAM|0.0|5|BEN & JERRY HALF BAKED|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00076840101320|ICE CREAM|FROZEN|-80.85753|80.85754234393255|218|1
35.116638|8340cab1b7e4fd813509c0a305231784b22682ab|3.89|2014-11-24 18:51:00|80.856688219393845|1|7684010015|204|35.132181951641783|0|15|275|-80.85013|45|35.175855|SUPER PREMIUM ICE CREAM|0.0|5|BEN & JERRY HALF BAKED|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00076840101320|ICE CREAM|FROZEN|-80.85753|80.85754234393255|218|1
35.116638|13fdfad26a39cd14031eec6a37c15bb84440fbea|3.89|2015-01-03 19:02:00|80.856688219393845|1|7684010015|204|35.132181947731389|0|15|275|-80.826724|45|35.195689|SUPER PREMIUM ICE CREAM|0.0|5|BEN & JERRY HALF BAKED|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00076840101320|ICE CREAM|FROZEN|-80.85753|80.857548278251102|412|1
35.116638|0ce463e78e1ba4a71a51c26a67f32116b2a97fbf|11.98|2014-11-20 20:12:00|80.856688219393845|1|7403008182|204|35.132181951641783|0|15|2017|-80.85013|505|35.175855|STRETCHED CURD CHEESE|2.99|6|SORRENTO FRESH MOZZARELLA|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00074030081827|SPECIALTY CHEESE|DELI|-80.85753|80.85754234393255|218|2
35.116638|fc236355262f49d119691526cd1ec37a4793844c|5.49|2015-02-08 18:23:00|80.856688219393845|1|7203688095|204|35.132181951641783|0|15|526|-80.85013|64|35.175855|FRESH MUSHROOMS|0.0|4|HT PORTOBELLO CAPS,TRAY|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00072036880956|FRESH PRODUCE|PRODUCE|-80.85753|80.85754234393255|218|1
35.116638|95ed0568cd5eef95a048f4367b343d6c56e48ea2|8.29|2014-09-20 09:46:00|80.856688219393845|1|4116710081|204|35.132181947731389|0|15|4388|-80.826724|1210|35.195689|ACID NEUTRALIZER-LIQUID|0.0|17|ROLAIDS ULTRA LIQUID CHERRY|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00041167100813|STOMACH REMEDIES|HBC|-80.85753|80.857548278251102|412|1
35.116638|8ed016536c1774415423ad595471eb7403e02c1c|8.29|2014-10-27 19:11:00|80.856688219393845|1|4116710081|204|35.13218194757431|0|15|4388|-80.844274|1210|35.204336|ACID NEUTRALIZER-LIQUID|0.0|17|ROLAIDS ULTRA LIQUID CHERRY|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00041167100813|STOMACH REMEDIES|HBC|-80.85753|80.857548476848805|61|1
35.116638|aa11645e2bcd54c45fee80b44fd5e30d033fd5fa|1.99|2014-11-22 15:43:00|80.856688219393845|1|3900004504|204|35.132181951641783|0|15|114|-80.85013|14|35.175855|PUMPKIN|0.2|1|LIBBY SOLID PACK PUMPKIN|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00039000045049|DESSERTS/GELS/SYRUPS|G1 GROCERY|-80.85753|80.85754234393255|218|1
35.116638|ed669551a8caa93440f8bb8a48a844604640b397|2.19|2015-02-24 17:24:00|80.856688219393845|1|76857300210|204|35.132181951641783|0|15|544|-80.85013|64|35.175855|FRESH PRODUCE FRSH HERBS|0.0|4|PKG FRESH SAGE|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00768573002202|FRESH PRODUCE|PRODUCE|-80.85753|80.85754234393255|218|1
35.116638|1c7c5c94e38881fe96b49f27cbdffedc00b3dede|2.19|2015-01-13 18:07:00|80.856688219393845|1|76857300210|204|35.132181951641783|0|15|544|-80.85013|64|35.175855|FRESH PRODUCE FRSH HERBS|0.0|4|PKG FRESH ITALIAN PARSLEY|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00768573002301|FRESH PRODUCE|PRODUCE|-80.85753|80.85754234393255|218|1
35.116638|282efc8ae73291bcf35535684fcfcc7e07c2bdd6|2.19|2014-11-03 18:01:00|80.856688219393845|1|76857300210|204|35.132181951641783|0|15|544|-80.85013|64|35.175855|FRESH PRODUCE FRSH HERBS|0.0|4|PKG FRESH ITALIAN PARSLEY|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00768573002301|FRESH PRODUCE|PRODUCE|-80.85753|80.85754234393255|218|1
35.116638|1e7fabc596a6fa6d0b1b82f21a1045bd8fda84c6|4.0|2014-10-15 21:21:00|80.856688219393845|1|65780295163|204|35.132181951641783|0|15|1165|-80.85013|87|35.175855|NFS-FRESH CONSUMER BUNCH|0.66|9|BUNCH- ALSTROEMERIA   RIVERD|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00657802951636|FLORAL|FLORAL|-80.85753|80.85754234393255|218|1
35.116638|2d804be64bfd3725f7949ddfb4caabc3c9de02aa|2.49|2014-09-18 17:31:00|80.856688219393845|1|60504939530|204|35.132181951641783|0|15|509|-80.85013|64|35.175855|FRESH CITRUS-REMAINING|0.0|4|LEMONS, SMALL 1LB BAG|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00605049395300|FRESH PRODUCE|PRODUCE|-80.85753|80.85754234393255|218|1
35.116638|cb20f58604ef11f4255cb0efd3f2aef26d6d72d0|12.0|2014-09-27 17:23:00|80.856688219393845|1|65780295163|204|35.132181951641783|0|15|1165|-80.85013|87|35.175855|NFS-FRESH CONSUMER BUNCH|0.0|9|BUNCH- ALSTROEMERIA   RIVERD|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00657802951636|FLORAL|FLORAL|-80.85753|80.85754234393255|218|3
35.116638|13d4802eeedcf6916b1756fd01dc8ccd7ebf7dfe|9.02|2015-03-05 17:38:00|80.856688219393845|1||204|35.132181951641783|0|15|500|-80.85013|64|35.175855|FRESH APPLES|0.0|4|HONEY CRISP APPLE|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00233283000003|FRESH PRODUCE|PRODUCE|-80.85753|80.85754234393255|218|1
35.116638|3b900bad1ecfd7486a29f250f5cbbd496d4851a6|4.82|2015-02-11 17:28:00|80.856688219393845|1||204|35.132181951641783|0|15|500|-80.85013|64|35.175855|FRESH APPLES|0.0|4|HONEY CRISP APPLE|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00233283000003|FRESH PRODUCE|PRODUCE|-80.85753|80.85754234393255|218|1
35.116638|3d1cd0fef2c6b4a83528c6ae749986844c9512e0|5.98|2014-09-17 20:32:00|80.856688219393845|1|5010017170|204|35.132181951641783|0|15|1499|-80.85013|33|35.175855|RTS MICROWAVE|0.0|1|HC MW SP CHS TORTELLINI|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00050100171926|SOUP|G1 GROCERY|-80.85753|80.85754234393255|218|2
35.116638|e8bd077fa319e196494f12a1c0a0efda3e1b0678|2.49|2014-11-09 19:14:00|80.856688219393845|1|7156766109|204|35.132181951641783|0|15|52|-80.85013|7|35.175855|PKG NON CHOC|0.0|1|JBELLY 20 FLAVORS|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00071567661096|CANDY|G1 GROCERY|-80.85753|80.85754234393255|218|1
35.116638|e8e3849c51f49900c92934e1622775d1f9c66066|1.2|2015-03-08 17:52:00|80.856688219393845|1|7047000641|204|35.132181951641783|0|15|688|-80.85013|61|35.175855|LIGHT|0.0|3|YOPLAIT LIGHT STRAWBERRY|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00070470006505|YOGURT|DAIRY|-80.85753|80.85754234393255|218|2
35.116638|9816d0ec735954cb72520d8cbda3c2862f2b8920|4.98|2014-09-10 15:33:00|80.856688219393845|1|7156766109|204|35.132181951641783|0|15|52|-80.85013|7|35.175855|PKG NON CHOC|0.0|1|JBELLY 20 FLAVORS|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00071567661096|CANDY|G1 GROCERY|-80.85753|80.85754234393255|218|2
35.116638|62cda5b8180145d48455502f42852f1f5f594e8f|3.59|2014-11-19 19:51:00|80.856688219393845|1|4850002013|204|35.132181951641783|0|15|335|-80.85013|56|35.175855|ORANGE JUICE-REGRIGERATED|0.59|3|TROPICANA PP HOMESTYLE|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00048500301395|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.85753|80.85754234393255|218|1
35.116638|e6fd06dd5a52577aa2640020b068bab24395fff6|10.98|2014-12-14 17:11:00|80.856688219393845|1|20895300000|204|35.132181951641783|0|15|977|-80.85013|201|35.175855|FRESH HT CHICKEN|5.49|2|HT FRESH BNLS CHICKEN BREAST|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00208953000003|POULTRY|MEAT|-80.85753|80.85754234393255|218|1
35.116638|47367fd57e8ec715e5ff33843a2f6cf26ad489f3|15.99|2015-02-15 14:49:00|80.856688219393845|1|3980000605|204|35.132181951641783|0|15|8445|-80.85013|1769|35.175855|ALKALINE C|0.0|18|(FE) ENERGIZER C FAMILY PK E|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00039800006059|BATTERY & FLASHLIGHT|GM|-80.85753|80.85754234393255|218|1
35.116638|1165bed6adc704faa44cc472a0fbb10f0e80420e|0.99|2014-11-13 18:46:00|80.856688219393845|1|7203676207|204|35.132181951641783|0|15|1218|-80.85013|273|35.175855|ASIAN OTHER|0.2|1|HT TRADER WATER CHESTNUTS SLIC|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00072036762078|ASIAN PREP. FOODS|G1 GROCERY|-80.85753|80.85754234393255|218|1
35.116638|5052384367cae590fc2d5e30692e3ccce1a8e9bb|0.99|2014-12-09 18:57:00|80.856688219393845|1|7203676207|204|35.132181951641783|0|15|1218|-80.85013|273|35.175855|ASIAN OTHER|0.0|1|HT TRADER WATER CHESTNUTS SLIC|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00072036762078|ASIAN PREP. FOODS|G1 GROCERY|-80.85753|80.85754234393255|218|1
35.116638|1befbe5d4475dae4221cb475bb728bfe17a469d5|2.69|2014-09-13 17:48:00|80.856688219393845|1|7203663996|204|35.132181951641783|0|15|342|-80.85013|57|35.175855|FRESH MILK|0.0|3|HARRIS TEETER WHOLE MILK|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00072036639967|MILK|DAIRY|-80.85753|80.85754234393255|218|1
35.116638|eb89d8876caa142502d4355c966dbcbbe0d6bdf8|16.72|2015-02-22 14:38:00|80.856688219393845|1|20249700000|204|35.132181951641783|0|15|297|-80.85013|49|35.175855|GROUND BEEF|0.84|2|NY STRIP STEAKBURGER 80% LEAN|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00202497000000|BEEF|MEAT|-80.85753|80.85754234393255|218|2
35.116638|0efdc1e64846adf66fabf38163be5355b2123c46|3.2|2015-01-23 17:56:00|80.856688219393845|1||204|35.132181951641783|0|15|531|-80.85013|64|35.175855|FRESH CORN|0.0|4|COO YELLOW CORN|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00204078000003|FRESH PRODUCE|PRODUCE|-80.85753|80.85754234393255|218|4
35.116638|67bfb17f1560076b7d777843c82e8a159450305b|6.98|2014-09-29 19:06:00|80.856688219393845|1||204|35.132181951641783|0|15|542|-80.85013|64|35.175855|FRESH VEGETABLES REMAIN|0.49|4|COO ARTICHOKES, JBO (RPC)|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00204084000004|FRESH PRODUCE|PRODUCE|-80.85753|80.85754234393255|218|2
35.116638|5cb5aee45d320bdca269b2acf4903ad7fedc6c21|2.29|2014-10-05 19:13:00|80.856688219393845|1||204|35.132181951641783|0|15|501|-80.85013|64|35.175855|FRESH PEARS|0.23|4|BOSC PEARS|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00204413000002|FRESH PRODUCE|PRODUCE|-80.85753|80.85754234393255|218|1
35.116638|5d7f2f589d99c35bcd7441e9c253d04c59e444ea|0.61|2015-02-14 18:28:00|80.856688219393845|1||204|35.132181951641783|0|15|524|-80.85013|64|35.175855|FRESH PROD FRESH ONIONS|0.0|4|COO YELLOW ONIONS, LRG|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00204665000003|FRESH PRODUCE|PRODUCE|-80.85753|80.85754234393255|218|1
35.116638|8b998c256b2ae176df14b9fefca7b25911bc37ee|4.19|2014-10-14 18:31:00|80.856688219393845|1|2100000201|204|35.132181951641783|0|15|317|-80.85013|52|35.175855|CHUNK AND BAR CHEESE|1.69|3|KRAFT SHARP CHEDDAR CHUNK|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00021000002016|CHEESE|DAIRY|-80.85753|80.85754234393255|218|1
35.116638|72ed4e992b572285f1a49006ca01518c2236ab39|5.39|2014-12-28 16:34:00|80.856688219393845|1|3000006720|204|35.132181951641783|0|15|1433|-80.85013|9|35.175855|GRANOLA|0.4|1|QKR NAT GRANOLA OAT HONEY RAIS|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00030000067208|CEREAL|G1 GROCERY|-80.85753|80.85754234393255|218|1
35.116638|b96262068989a072ad0f4e33edca9b60bbb2fe20|5.39|2015-01-17 19:13:00|80.856688219393845|1|3000006720|204|35.132181951641783|0|15|1433|-80.85013|9|35.175855|GRANOLA|0.6|1|QKR NAT GRANOLA OAT HONEY RAIS|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00030000067208|CEREAL|G1 GROCERY|-80.85753|80.85754234393255|218|1
35.116638|9acc7ead512ae3d7335408d3e265459bd3e9aa68|1.39|2014-10-12 16:04:00|80.856688219393845|1|4150005807|204|35.132181951641783|0|15|80|-80.85013|34|35.175855|SEASONING PACKETS|0.0|1|FRENCH'S ORIGINAL CHILI-O|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00041500058078|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.85753|80.85754234393255|218|1
35.116638|6502a88c9d3340f3bda3f312f38500c4cf5a0e60|2.85|2014-12-07 17:17:00|80.856688219393845|1|4400000055|204|35.132181951641783|0|15|88|-80.85013|13|35.175855|FLAKED SODA CRACKERS|0.35|1|NABISCO PREMIUMS|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00044000000578|CRACKERS|G1 GROCERY|-80.85753|80.85754234393255|218|1
35.116638|895aa4a6355a0b0cfe27c3c7bab79d1f13ddd860|1.79|2014-11-26 19:21:00|80.856688219393845|1|7203663157|204|35.132181951641783|0|15|1134|-80.85013|57|35.175855|CARTON MILK|0.0|3|HARRIS TEETER WHOLE MILK|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00072036631572|MILK|DAIRY|-80.85753|80.85754234393255|218|1
35.116638|352aa3382991b26cb5f9269efa1cebd3e17f8981|3.67|2014-10-21 19:20:00|80.856688219393845|1|7203655019|204|35.132181951641783|0|15|332|-80.85013|52|35.175855|STRING/SNACK|0.0|3|HT STRING CHEESE|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00072036550194|CHEESE|DAIRY|-80.85753|80.85754234393255|218|1
35.116638|4f932fc0eb10f4a04218330ad4a6c43f3a6e5aea|8.69|2014-10-16 19:31:00|80.856688219393845|1|7203653118|204|35.132181951641783|0|15|1243|-80.85013|21|35.175855|MIXED NUTS CASHEWS|2.7|1|HT CASHEWS HALVES|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00072036531186|NUTS|G1 GROCERY|-80.85753|80.85754234393255|218|1
35.116638|8ef0df2cbee92850624e4a865c8cd2d90b681b27|3.69|2015-02-19 17:33:00|80.856688219393845|1|7127925101|204|35.132181951641783|0|15|555|-80.85013|64|35.175855|PACKAGED SALADS|0.0|4|F.E. AMERICAN SALAD|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00071279241005|FRESH PRODUCE|PRODUCE|-80.85753|80.85754234393255|218|1
35.116638|4e3b7137f6c67c27a789da2bb9d3a07133d2057f|4.49|2014-10-01 20:13:00|80.856688219393845|1|87989000001|204|35.132181947731389|0|15|1982|-80.826724|480|35.195689|DRY GOODS CRACKERS|0.0|6|ORIGINAL MULTI-SEED CRACKERS|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00879890000014|DRY GOODS|DELI|-80.85753|80.857548278251102|412|1
35.116638|43ce105b480db6d687317c06d3f1d0fcd625ad82|1.49|2014-12-16 20:17:00|80.856688219393845|1|1530044051|204|35.132181951641783|0|15|1439|-80.85013|274|35.175855|DRY DINNERS|0.0|1|PASTA RONI ANGEL HAIR HERB|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00015300440517|PREP FOODS DINNERS|G1 GROCERY|-80.85753|80.85754234393255|218|1
35.116638|4d81a4927a8788cc4d0f8c952356b175eb6a89c7|9.99|2014-10-25 19:22:00|80.856688219393845|1|83074600117|204|35.132181942070169|0|15|458|-80.810056|82|35.219587|CRAFT BEER|0.0|16|GREEN FLASH WEST COAST IPA 4PK|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00830746001173|DOMESTIC BEER|BEER|-80.85753|80.857554437239529|401|1
35.116638|d6761b7ddb92e38a194f69da300ca9e729cee877|1.38|2014-09-25 18:15:00|80.856688219393845|1||204|35.132181951641783|0|15|505|-80.85013|64|35.175855|FRESH SOFT FRUIT|0.1|4|WHITE NECTARINES PLU#|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00233035000008|FRESH PRODUCE|PRODUCE|-80.85753|80.85754234393255|218|1
35.116638|99f94a58a004acd65b78d5e766711000dfe8519a|4.39|2015-01-15 19:30:00|80.856688219393845|1|4400003037|204|35.132181951641783|0|15|90|-80.85013|13|35.175855|SNACK CRACKERS|1.39|1|WHEAT THINS ORIGINAL|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00044000030377|CRACKERS|G1 GROCERY|-80.85753|80.85754234393255|218|1
35.116638|000ff081f3887d28de44057310f0114c7716b1c0|9.98|2014-12-17 20:33:00|80.856688219393845|1|7146426060|204|35.132181951641783|0|15|577|-80.85013|136|35.175855|OTHER MERCH FR MSC JUICE|0.0|4|BOLTHOUSE CARROT JUICE|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00071464200602|OTHER MERCHANDISE|PRODUCE|-80.85753|80.85754234393255|218|2
35.116638|8baa2a741a7df92df5693745cd94e9cd4199310c|8.89|2014-11-06 18:09:00|80.856688219393845|1|1410009655|204|35.132181951641783|0|15|87|-80.85013|13|35.175855|CHEESE CRACKERS|0.9|1|PF BULK GOLDFISH CHEDDAR|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00014100096559|CRACKERS|G1 GROCERY|-80.85753|80.85754234393255|218|1
35.116638|f873f86c058e67115f8e4ccea5454d881afe34a2|2.89|2014-10-26 19:27:00|80.856688219393845|1|3120000293|204|35.132181951641783|0|15|116|-80.85013|17|35.175855|DRIED CRANBERRIES|0.39|1|OS CRAISIN CHERRY FLAVOR|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00031200002921|FRUIT-DRIED|G1 GROCERY|-80.85753|80.85754234393255|218|1
35.116638|420a3f529339860bf008734f8e03f74d6bd2f408|3.79|2015-02-11 20:16:00|80.856688219393845|1|7684010015|204|35.132181951641783|0|15|275|-80.85013|45|35.175855|SUPER PREMIUM ICE CREAM|0.0|5|BEN&JERRY COFFEE TOFFEE CRUNCH|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00076840100118|ICE CREAM|FROZEN|-80.85753|80.85754234393255|218|1
35.116638|c152057db4afa0ef83af9d5056f7b6c04b9acde3|3.79|2015-01-18 17:58:00|80.856688219393845|1|7684010015|204|35.132181951641783|0|15|275|-80.85013|45|35.175855|SUPER PREMIUM ICE CREAM|0.0|5|BEN&JERRY COFFEE TOFFEE CRUNCH|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00076840100118|ICE CREAM|FROZEN|-80.85753|80.85754234393255|218|1
35.116638|5e84e972ac7e0b06638d1439dc1ecd8831494ba5|12.89|2014-11-30 17:26:00|80.856688219393845|1|30005475756|204|35.132181951641783|0|15|4615|-80.85013|1215|35.175855|VITAMIN-MULTIPLE-ADULT|0.0|17|CENTRUM MEN|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00300054757562|VITAMINS & SUPPLEMENTS|HBC|-80.85753|80.85754234393255|218|1
35.116638|d0ebfc5b02f92f5040062db21180614d38d8b7c6|0.63|2014-10-09 19:34:00|80.856688219393845|1||204|35.132181951641783|0|15|522|-80.85013|64|35.175855|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00204664000004|FRESH PRODUCE|PRODUCE|-80.85753|80.85754234393255|218|1
35.116638|29d7153aefc48f90c12d633b90035f2ba9512f70|1.15|2014-10-06 17:59:00|80.856688219393845|1|7203614992|204|35.132181951641783|0|15|115|-80.85013|16|35.175855|REMAINING FRUIT|0.15|1|HT MANDARIN ORANGE LS|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00072036146687|FRUIT-CAN/JAR|G1 GROCERY|-80.85753|80.85754234393255|218|1
35.116638|e394193a939b4f14db4f4e5ab7bb5e1f51792d5f|1.89|2014-10-07 19:35:00|80.856688219393845|1|2400034616|204|35.132181951641783|0|15|1221|-80.85013|275|35.175855|PASTA SC VALUE|0.0|1|CONTADINA SQZ PIZZA SC|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00024000346166|PASTA SAUCES|G1 GROCERY|-80.85753|80.85754234393255|218|1
35.116638|9364346766b781d06454c468a11de95b9a3d9efc|5.9|2014-12-16 21:02:00|80.856688219393845|1|7203663125|204|35.132181947731389|0|15|1262|-80.826724|57|35.195689|HALF N HALF WHIPPING CREAM|1.9|3|HT WHIPPING CREAM|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00072036631251|MILK|DAIRY|-80.85753|80.857548278251102|412|2
35.116638|524395e46ac52674f2c7a4bf161ecd52d6b5de9a|3.35|2014-12-31 07:58:00|80.856688219393845|1|1600042040|204|35.132181951641783|0|15|13|-80.85013|2|35.175855|ROLLS/BISCUIT MIXES|0.0|1|BC BISQUICK|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00016000420403|BAKING MIXES|G1 GROCERY|-80.85753|80.85754234393255|218|1
35.116638|57e161eb9e8fce23128fa8d889028c620ed7e8cd|2.19|2014-11-04 17:32:00|80.856688219393845|1|31254662542|204|35.132181951641783|0|15|4207|-80.85013|1200|35.175855|COUGH DROP-ADULT|0.0|17|HALLS SF H/LEMON 62213|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00312546622135|COUGH/COLD/SINUS|HBC|-80.85753|80.85754234393255|218|1
35.116638|1b8df3fe313e1cb97bd6f383a413c152be555111|3.69|2014-09-28 17:41:00|80.856688219393845|1|5000012734|204|35.132181951641783|0|15|341|-80.85013|57|35.175855|CREAMERS|1.19|3|COFFEEMATE FRENCH VANILLA|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00050000322756|MILK|DAIRY|-80.85753|80.85754234393255|218|1
35.116638|a7eae2458e152075a2cb04620703805af80cedea|3.39|2014-11-02 19:51:00|80.856688219393845|1|5000012734|204|35.132181951641783|0|15|341|-80.85013|57|35.175855|CREAMERS|0.0|3|COFFEEMATE FRENCH VANILLA|5f1c0f580d2899c6f85f020d8a43ef86b7cedb84|1.0740497477077775|35.134355925261694|00050000322756|MILK|DAIRY|-80.85753|80.85754234393255|218|1
34.937113|c31ed6e517775b565a663e7224760cd8f35ed55c|2.39|2014-09-11 18:14:00|80.828402574597021|4|5100002549|372|35.201287466225793|0|8|1221|-81.027334|275|34.977331|PASTA SC VALUE|0.39|1|PREGO SC TRADITIONAL|5f44b7d54e2bd5cbfd35363afb882fabb5cb9472|18.253819376591427|35.209978091326001|00051000025494|PASTA SAUCES|G1 GROCERY|-80.837892|80.838032073693185|149|1
34.937113|316cf96743109e543b56653b65337dbabb9d1c87|11.98|2015-01-27 18:03:00|80.828402574597021|4|20526100000|372|35.201287466225793|0|8|1935|-81.027334|465|34.977331|CHEF CASE|0.0|6|LUMP CRABCAKES|5f44b7d54e2bd5cbfd35363afb882fabb5cb9472|18.253819376591427|35.209978091326001|00205261000008|COLD PREPARED FOODS|DELI|-80.837892|80.838032073693185|149|1
34.937113|924e43de66b024df15ad3e4a56533f778a7922a6|2.59|2014-11-11 18:21:00|80.828402574597021|4|7203663996|372|35.201287466225793|0|8|342|-81.027334|57|34.977331|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|5f44b7d54e2bd5cbfd35363afb882fabb5cb9472|18.253819376591427|35.209978091326001|00072036631299|MILK|DAIRY|-80.837892|80.838032073693185|149|1
34.937113|d36d10ca5c97fc179a7d863e9fe162660832a63e|17.26|2014-10-07 18:32:00|80.828402574597021|4|5000|372|35.201287466225793|0|8|49|-81.027334|7|34.977331|BULK CANDY|9.27|1|JBELLY PLU#|5f44b7d54e2bd5cbfd35363afb882fabb5cb9472|18.253819376591427|35.209978091326001|00000000050000|CANDY|G1 GROCERY|-80.837892|80.838032073693185|149|1
35.43259|e2ac01ef599322558347d76c664afcf5c8846600|7.99|2014-12-19 12:45:00|1.4057311447477159|3|31284353637|202|0.6184153580092175|0|52|4308|-80.605588|1205|35.43259|ASPIRIN|0.0|17|EBAYER 81MG REGIMEN|5f55d4cf2d4b946f6749d8c117f2527c71f3c3d5|9.70732144626205|0.6209993146566879|00312843536371|PAIN RELIEF|HBC|-80.605588|1.406832906106031|202|1
35.43259|86a0ede51844ccbdc80f5fec3ee9f6c165648141|10.71|2014-09-12 11:34:00|1.4057311447477159|3|20891800000|202|0.6184153580092175|0|52|657|-80.605588|201|35.43259|STR MDE VALUE ADD POLTRY|1.34|2|SKEWERED CHICKEN KABOB|5f55d4cf2d4b946f6749d8c117f2527c71f3c3d5|9.70732144626205|0.6209993146566879|00208919000009|POULTRY|MEAT|-80.605588|1.406832906106031|202|1
35.43259|09bf09e081077a09551b1594df82989855168364|2.65|2015-01-09 11:53:00|1.4057311447477159|3|4119691401|202|0.6184153580092175|0|52|1201|-80.605588|33|35.43259|RTS CANNED|0.0|1|PROG RICH HRT STEAK BURGER VEG|5f55d4cf2d4b946f6749d8c117f2527c71f3c3d5|9.70732144626205|0.6209993146566879|00041196421699|SOUP|G1 GROCERY|-80.605588|1.406832906106031|202|1
35.43259|4de7706258d30e722ddb4a6dfd713df783bc2e74|4.59|2014-10-17 12:39:00|1.4057311447477159|3|7033041756|202|0.6184153580092175|0|52|6680|-80.605588|1564|35.43259|MECHANICAL PENCIL|0.0|18|BIC MECH PENCIL METALLIC .5MM|5f55d4cf2d4b946f6749d8c117f2527c71f3c3d5|9.70732144626205|0.6209993146566879|00070330417564|SCHOOL & OFFICE SUPPLY|GM|-80.605588|1.406832906106031|202|1
35.43259|bfe303ae690a8556f8efc76adcf0230103aa21a3|14.19|2014-10-24 11:22:00|1.4057311447477159|3|7023015366|202|0.6184153580092175|0|52|730|-80.605588|24|35.43259|NFS-CAT LITTER|0.0|1|TIDY CATS LGHTWEIGHT LITTR 8.5|5f55d4cf2d4b946f6749d8c117f2527c71f3c3d5|9.70732144626205|0.6209993146566879|00070230153661|PET FOOD/SUPPLIES|G1 GROCERY|-80.605588|1.406832906106031|202|1
35.43259|7ec787b5499d97aff087de1333965c5a71b44c7d|1.79|2015-01-30 11:53:00|1.4057311447477159|3|5100001047|202|0.6184153580092175|0|52|212|-80.605588|33|35.43259|CONDENSED SOUP|0.54|1|CAMP COND NEW ENG CLAM CHOWDER|5f55d4cf2d4b946f6749d8c117f2527c71f3c3d5|9.70732144626205|0.6209993146566879|00051000013675|SOUP|G1 GROCERY|-80.605588|1.406832906106031|202|1
35.43259|25cf011c10461bbea5eccc60197384bac298d019|2.69|2014-12-05 13:27:00|1.4057311447477159|3|4114312010|202|0.6184153580092175|0|52|119|-80.605588|17|35.43259|RAISINS|0.0|1|SUN MAID 6PK RAISINS|5f55d4cf2d4b946f6749d8c117f2527c71f3c3d5|9.70732144626205|0.6209993146566879|00041143120101|FRUIT-DRIED|G1 GROCERY|-80.605588|1.406832906106031|202|1
35.43259|23fb7d1907d306485075afaed3a4d35d490d3712|3.99|2014-11-01 17:24:00|80.606823361882718|3|7005700120|202|35.573077086425243|0|57|677|-80.746334|150|35.41832|SEASONINGS|0.0|12|PHILLIPS BLACKENING SEASONING|5f55d4cf2d4b946f6749d8c117f2527c71f3c3d5|9.70732144626205|35.500309569604553|00070057001206|CONDIMENTS|SEAFOOD|-80.605588|80.605724539114249|190|1
35.024332|8718dd3de04e25231e07ea9cc99646a00d44df88|1.89|2014-10-24 14:55:00|1.4091206135396188|2|4150000025|343|0.6112899117116106|0|47|78|-80.760919|11|35.024332|MUSTARD|0.04|1|FRENCHS MUSTARD YELLOW 14|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00041500000251|CONDIMENTS|G1 GROCERY|-80.760919|1.4095439434864463|343|1
35.024332|5659192d2810bc6dba76ca10a7fda18097a55c4f|3.49|2015-01-02 15:53:00|1.4091206135396188|2|3800001611|343|0.6112899117116106|0|47|61|-80.760919|9|35.024332|RTE CEREAL ADULT|0.99|1|KELLOGG SPECIAL K 12 OZ BOX|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00038000016110|CEREAL|G1 GROCERY|-80.760919|1.4095439434864463|343|1
35.024332|0621f4c0bb2dc2a1753b24bf3bd9a498780ae297|3.69|2014-09-23 15:04:00|1.4091206135396188|2|3700025574|343|0.6112899117116106|0|47|725|-80.760919|66|35.024332|NFS-DISHWASHING LIQUID|0.69|1|IVORY LIQ DISH GENTLE CLASSIC|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00037000255741|DETERGENTS|G1 GROCERY|-80.760919|1.4095439434864463|343|1
35.024332|5585d59317895648f5a309f85fd6dcd89c345858|3.49|2015-01-29 14:39:00|1.4091206135396188|2|3800001611|343|0.6112899117116106|0|47|61|-80.760919|9|35.024332|RTE CEREAL ADULT|0.0|1|KELLOGG SPECIAL K 12 OZ BOX|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00038000016110|CEREAL|G1 GROCERY|-80.760919|1.4095439434864463|343|1
35.024332|83d289356fa3a2967aff8a027e2e35934b877b8f|3.49|2015-02-05 14:07:00|1.4091206135396188|2|3800001611|343|0.6112899117116106|0|47|61|-80.760919|9|35.024332|RTE CEREAL ADULT|0.0|1|KELLOGG SPECIAL K 12 OZ BOX|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00038000016110|CEREAL|G1 GROCERY|-80.760919|1.4095439434864463|343|1
35.024332|dd2776a69515f06405d36a6e1f0099f92165eaaa|3.69|2015-01-10 17:28:00|1.4091206135396188|2|7203698007|343|0.6112899117116106|0|47|423|-80.760919|72|35.024332|NFS-DISPOSE PLATES/BOWLS|1.19|1|"YH 9"" HEAVY DUTY PAPER PLATES"|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00072036980076|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.760919|1.4095439434864463|343|1
35.024332|0e1a2c54ae29822bb877e183ba697296d1d60d7a|2.99|2015-03-02 16:56:00|1.4091206135396188|2|81204900640|343|0.6112899117116106|0|47|504|-80.760919|64|35.024332|FRESH BERRIES|0.0|4|BLUEBERRIES 6 OZ|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00891700002124|FRESH PRODUCE|PRODUCE|-80.760919|1.4095439434864463|343|1
35.024332|bcb7602cee437ec457ee81125bc2effbba8b264e|3.79|2015-03-06 15:04:00|1.4091206135396188|2|4470000063|343|0.6112899117116106|0|47|359|-80.760919|101|35.024332|MEAT WIENERS|0.0|19|OSCAR MAYER WIENER|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00044700000632|WIENERS|CASE READY MEATS|-80.760919|1.4095439434864463|343|1
35.024332|b448017ec6fc0e1a164e86c4e39023ab10e8d5a9|3.49|2014-10-06 12:29:00|1.4091206135396188|2|4470000063|343|0.6112899117116106|0|47|359|-80.760919|101|35.024332|MEAT WIENERS|0.0|19|OSCAR MAYER WIENER|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00044700000632|WIENERS|CASE READY MEATS|-80.760919|1.4095439434864463|343|1
35.024332|1a98f1f6e7b70dc8d80b51fe404aa402858c627f|1.99|2015-01-21 12:59:00|1.4091206135396188|2|5100002549|343|0.6112899117116106|0|47|1221|-80.760919|275|35.024332|PASTA SC VALUE|0.32|1|PREGO SC TRADITIONAL|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00051000025494|PASTA SAUCES|G1 GROCERY|-80.760919|1.4095439434864463|343|1
35.024332|8e9fc72e718fabb9c9f4e4660ca2934fe9f2914d|11.85|2015-01-24 10:23:00|1.4091206135396188|2|74816261452|343|0.6112899117116106|0|47|1460|-80.760919|40|35.024332|FROZEN BREAD AND ROLLS|0.0|5|SCHUBERTS DINNER YEAST ROLLS|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00748162621021|FROZEN DOUGH|FROZEN|-80.760919|1.4095439434864463|343|3
35.024332|811a881783d236717e988694522a076abc10179e|3.95|2015-02-16 13:31:00|1.4091206135396188|2|74816261452|343|0.6112899117116106|0|47|1460|-80.760919|40|35.024332|FROZEN BREAD AND ROLLS|0.0|5|SCHUBERTS DINNER YEAST ROLLS|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00748162621021|FROZEN DOUGH|FROZEN|-80.760919|1.4095439434864463|343|1
35.024332|ff1a73252055ca2fcc4d5bd45143dec71ce95052|3.95|2014-12-16 15:20:00|1.4091206135396188|2|74816261452|343|0.6112899117116106|0|47|1460|-80.760919|40|35.024332|FROZEN BREAD AND ROLLS|1.45|5|SCHUBERTS DINNER YEAST ROLLS|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00748162621021|FROZEN DOUGH|FROZEN|-80.760919|1.4095439434864463|343|1
35.024332|1a7c4f1a9463c0240c37ccb5253e8251abebc9a3|11.75|2014-09-18 14:52:00|1.4091206135396188|2|20140400000|343|0.6112899117116106|0|47|296|-80.760919|49|35.024332|RANCHER BEEF|0.0|2|BEEF LOIN NY STRIP STEAK BNLS|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00201404000003|BEEF|MEAT|-80.760919|1.4095439434864463|343|1
35.024332|a74aa49e11c0ca08f43f4243f199e053457b1a95|3.58|2014-12-01 17:46:00|80.805842308733688|2|5100005977|343|35.058763625319919|0|49|212|-80.758228|33|34.95459|CONDENSED SOUP|0.24|1|CAMP HLTHY REQ CREAM MUSHROOM|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|35.053350220983141|00051000060075|SOUP|G1 GROCERY|-80.760919|80.760949072798837|182|2
35.024332|cd095ce5d3db95c0719c1845e4cb620bdbf4086f|3.49|2014-10-30 13:04:00|80.805842308733688|2|20455000000|343|35.058763625319919|0|49|542|-80.758228|64|34.95459|FRESH VEGETABLES REMAIN|0.0|4|BRUSSEL SPROUTS 1LB (RPC)|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|35.053350220983141|00094922577160|FRESH PRODUCE|PRODUCE|-80.760919|80.760949072798837|182|1
35.024332|83e8f876c5979855504bd8c950a4f93524326478|2.49|2014-12-23 16:13:00|1.4091206135396188|2|60504939530|343|0.6112899117116106|0|47|509|-80.760919|64|35.024332|FRESH CITRUS-REMAINING|0.0|4|LEMONS, SMALL 1LB BAG|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00605049395300|FRESH PRODUCE|PRODUCE|-80.760919|1.4095439434864463|343|1
35.024332|4126c0d6696c13ddf4e0da584b2bcfeb7ad00a50|1.29|2014-10-07 17:56:00|1.4091206135396188|2|2700041916|343|0.6112899117116106|0|47|95|-80.760919|14|35.024332|SINGLE/SERVE R-T-S DESSERTS|0.29|1|SNACK PACK VANILLA|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00027000419014|DESSERTS/GELS/SYRUPS|G1 GROCERY|-80.760919|1.4095439434864463|343|1
35.024332|868de563de4ac8d2a0953d5b205d0236887fec86|4.79|2015-02-23 16:23:00|1.4091206135396188|2|37513770335|343|0.6112899117116106|0|47|4820|-80.760919|1235|35.024332|ADHESIVE BANDAGE LIQ PWD PST|0.0|17|NEW SKIN LIQUID BANDAGE|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00375137703354|FIRST AID|HBC|-80.760919|1.4095439434864463|343|1
35.024332|acb1a8c8f1231784e26a97d70500e8fa49af294d|4.99|2014-11-18 15:17:00|1.4091206135396188|2|7203688079|343|0.6112899117116106|0|47|523|-80.760919|64|35.024332|FRESH POTATOES|0.0|4|HT WHITE POTATO 5LB BAG|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00072036880796|FRESH PRODUCE|PRODUCE|-80.760919|1.4095439434864463|343|1
35.024332|cc92adff812dc5820c6e3e3c09a87b3811c1756c|4.29|2014-12-27 15:59:00|1.4091206135396188|2|74816261502|343|0.6112899117116106|0|47|1460|-80.760919|40|35.024332|FROZEN BREAD AND ROLLS|1.29|5|SCHUBERTS SWT HAWAIIAN ROLLS|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00748162615020|FROZEN DOUGH|FROZEN|-80.760919|1.4095439434864463|343|1
35.024332|228e538179a3ec0910413be1fc86cc86ee9de77a|3.69|2014-10-14 13:03:00|1.4091206135396188|2|2059300015|343|0.6112899117116106|0|47|1459|-80.760919|40|35.024332|FROZEN BISCUITS|0.0|5|MARY B'S THIN BISCUITS|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00020593000287|FROZEN DOUGH|FROZEN|-80.760919|1.4095439434864463|343|1
35.024332|6cc49c921efa6b543e4b7ca0e64704be982ed06e|5.89|2015-01-12 15:41:00|1.4091206135396188|2|5210000396|343|0.6112899117116106|0|47|1245|-80.760919|34|35.024332|SINGLE SPICES|0.0|1|E  MC CILANTRO LEAVES|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00052100003962|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.760919|1.4095439434864463|343|1
35.024332|32f51608a3b9bdd9ed2199312e69659109850378|7.99|2015-01-12 15:21:00|1.4091206135396188|2|31284353637|343|0.6112899117116106|0|47|4308|-80.760919|1205|35.024332|ASPIRIN|0.0|17|EBAYER 81MG REGIMEN|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00312843536371|PAIN RELIEF|HBC|-80.760919|1.4095439434864463|343|1
35.024332|8dec72a0521f0b677ece330c51010e4cb9597b08|5.39|2015-02-27 12:19:00|1.4091206135396188|2|4116710041|343|0.6112899117116106|0|47|4394|-80.760919|1210|35.024332|ACID NEUTRALIZER-SWALLOW|1.4|17|ROLAIDS ULTRA FRUIT TABLETS|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00041167100417|STOMACH REMEDIES|HBC|-80.760919|1.4095439434864463|343|1
35.024332|d5641469c59678dfadd399696cb776b2c86458be|3.99|2014-12-12 14:44:00|1.4091206135396188|2|5783602064|343|0.6112899117116106|0|47|522|-80.760919|64|35.024332|FRESH TOMATOES|0.0|4|CAMPARI TOMATO 16 OZ|6126a902933e6e25f25bada1cf10bd6cba737c98|2.379142768498045|0.61242566243833529|00057836020641|FRESH PRODUCE|PRODUCE|-80.760919|1.4095439434864463|343|1
35.318911|e2481e7613c11fd8e3a6ecb916b3f90e20ca04ac|1.16|2014-11-16 18:45:00|80.780380710856576|2||167|35.350705649277756|0|48|524|-80.737839|64|35.297134|FRESH PROD FRESH ONIONS|0.0|4|COO YELLOW ONIONS, LRG|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00204665000003|FRESH PRODUCE|PRODUCE|-80.780702|80.78070323080172|258|1
35.318911|76b8ea496edc715cc0a5fca5f238d2583d81dcb7|13.99|2014-11-26 23:50:00|80.780380710856576|2|8200072908|167|35.350705649277756|0|48|461|-80.737839|84|35.297134|FLAVORED MALT BEVERAGE|0.0|16|SMIRNOFF TWISTED VARIETY 12PK|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00082000729082|SPECIALTY|BEER|-80.780702|80.78070323080172|258|1
35.318911|8ac2e457ec2109815608cf3f5a02821faf5d2ab5|1.25|2015-02-26 20:36:00|80.780380710856576|2|5100002421|167|35.350705649277756|0|48|214|-80.737839|33|35.297134|BROTH|0.0|1|SWANSON BROTH CHICKEN|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00051000024312|SOUP|G1 GROCERY|-80.780702|80.78070323080172|258|1
35.318911|546be9193b99a529a0cecc136edd499a70f4ac5a|11.99|2014-09-12 13:36:00|80.780380710856576|2|2301286481|167|35.350705610304743|0|48|1477|-80.80146|485|35.17739|SUSHI HYBRID|0.0|6|"CHEF SAMPLER ""A"""|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00023012864811|SUSHI|DELI|-80.780702|80.780763035958614|208|1
35.318911|a63740bef608a96bea6a69dce323e7ac0aaf3390|2.38|2015-02-08 22:01:00|80.780380710856576|2|2970000146|167|35.350705649277756|0|48|165|-80.737839|26|35.297134|DEHYDRATED POTATOES|0.0|1|IDAHOAN MASHD APPLWD SMK BACON|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00029700021504|PREPARED FOODS-DRY MIXES|G1 GROCERY|-80.780702|80.78070323080172|258|2
35.318911|c65b4db54674214024b82715858ac2a00889d85d|2.38|2014-11-23 23:29:00|80.780380710856576|2|2970000146|167|35.350705649277756|0|48|165|-80.737839|26|35.297134|DEHYDRATED POTATOES|0.0|1|IDAHOAN MASHD APPLWD SMK BACON|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00029700021504|PREPARED FOODS-DRY MIXES|G1 GROCERY|-80.780702|80.78070323080172|258|2
35.318911|99e0ab2f97ff013f28263d84ed9e8cfe9bde47b0|3.57|2014-11-30 16:44:00|80.780380710856576|2|2970000146|167|35.350705649277756|0|48|165|-80.737839|26|35.297134|DEHYDRATED POTATOES|0.0|1|IDAHOAN MASHD LOADED|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00029700001483|PREPARED FOODS-DRY MIXES|G1 GROCERY|-80.780702|80.78070323080172|258|3
35.318911|ad76d3b2fe4924aae88ed95e28e5e14a88a7b978|1.19|2014-11-19 22:19:00|80.780380710856576|2|2970000146|167|35.350705649277756|0|48|165|-80.737839|26|35.297134|DEHYDRATED POTATOES|0.0|1|IDAHOAN MASHD LOADED|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00029700001483|PREPARED FOODS-DRY MIXES|G1 GROCERY|-80.780702|80.78070323080172|258|1
35.318911|b2b3d363ccc5c769641575626fb98d87de768e63|4.0|2014-12-20 22:57:00|80.780380710856576|2|66440177739|167|35.350705649277756|0|48|1165|-80.737839|87|35.297134|NFS-FRESH CONSUMER BUNCH|0.0|9|BUNCH- JUMBO SUNFLOWER 3 ST|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00664401777390|FLORAL|FLORAL|-80.780702|80.78070323080172|258|1
35.318911|3727e54d80c1b200b2194a84eda20ab58e1f1c6b|4.0|2015-02-21 18:37:00|80.780380710856576|2|66440177739|167|35.350705649277756|0|48|1165|-80.737839|87|35.297134|NFS-FRESH CONSUMER BUNCH|0.0|9|BUNCH- JUMBO SUNFLOWER 3 ST|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00664401777390|FLORAL|FLORAL|-80.780702|80.78070323080172|258|1
35.318911|7a60ad92ca4519b08db034993f9e0866a43b63d3|2.19|2014-11-12 19:10:00|80.780380710856576|2|76857300210|167|35.350705649277756|0|48|544|-80.737839|64|35.297134|FRESH PRODUCE FRSH HERBS|0.0|4|PKG FRESH DILL|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00768573002103|FRESH PRODUCE|PRODUCE|-80.780702|80.78070323080172|258|1
35.318911|bd6f39318e8732bb6bbb218d80c0dadae07a5cb5|0.89|2015-01-12 23:25:00|80.780380710856576|2||167|35.350705649277756|0|48|507|-80.737839|64|35.297134|FRESH ORANGES|0.1|4|NAVEL ORANGE, LRG|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00233107000004|FRESH PRODUCE|PRODUCE|-80.780702|80.78070323080172|258|1
35.318911|e6ced2338cdf58b49125d657c86fb879a66e065b|0.89|2014-09-18 21:24:00|80.780380710856576|2||167|35.350705649277756|0|48|507|-80.737839|64|35.297134|FRESH ORANGES|0.0|4|NAVEL ORANGE, LRG|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00233107000004|FRESH PRODUCE|PRODUCE|-80.780702|80.78070323080172|258|1
35.318911|1eb11381c8cd83ca3fb57db568eb1d462ef9d1f8|5.98|2014-12-23 18:04:00|80.780380710856576|2|4144900210|167|35.350705649277756|0|48|231|-80.737839|37|35.297134|INSTANT TEA|0.98|1|ALPINE SPICED CIDER REGULAR|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00041449002101|TEA|G1 GROCERY|-80.780702|80.78070323080172|258|2
35.318911|7d4fa67c3b01461faa24241fc04574eb920ca5ab|2.99|2014-11-05 18:59:00|80.780380710856576|2|4144900210|167|35.350705649277756|0|48|231|-80.737839|37|35.297134|INSTANT TEA|0.49|1|ALPINE SPICED CIDER REGULAR|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00041449002101|TEA|G1 GROCERY|-80.780702|80.78070323080172|258|1
35.318911|c8088e174a799ff90444b5f7d1d9dfabc8139af8|3.49|2015-01-29 23:25:00|80.780380710856576|2|2389649770|167|35.350705649277756|0|48|200|-80.737839|31|35.297134|MICROWAVE POPCORN|0.0|1|POPSECRET HOME STYLE 3 CT|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00023896246802|SNACKS|G1 GROCERY|-80.780702|80.78070323080172|258|1
35.318911|23b578a82672510da39de73a9a43d118459c0c20|3.85|2015-01-05 21:49:00|80.780380710856576|2|2100060464|167|35.350705649277756|0|48|315|-80.737839|52|35.297134|CHEESE-PROCESSED-SLICED|0.0|3|KRAFT SHARP CHEDDAR SINGLES|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00021000616480|CHEESE|DAIRY|-80.780702|80.78070323080172|258|1
35.318911|de0e5fc7fd43f7784b39504b990ca8755a3f959f|3.85|2014-12-15 01:03:00|80.780380710856576|2|2100060464|167|35.350705649277756|0|48|315|-80.737839|52|35.297134|CHEESE-PROCESSED-SLICED|0.85|3|KRAFT SHARP CHEDDAR SINGLES|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00021000616480|CHEESE|DAIRY|-80.780702|80.78070323080172|258|1
35.318911|54ed4f2981ec838adc7fa062cc27c102454df6fa|7.99|2014-11-02 17:03:00|80.780380710856576|2|1497490009|167|35.350705649277756|0|48|463|-80.737839|84|35.297134|HARD CIDER|0.0|16|WOODCHUCK SEASONAL 6PK|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00014974900099|SPECIALTY|BEER|-80.780702|80.78070323080172|258|1
35.318911|9f06ac162ac2dd169abb27b10b878b6441948ed3|2.59|2014-12-27 00:37:00|80.780380710856576|2|2073509418|167|35.350705649277756|0|48|365|-80.737839|56|35.297134|REFRIGERATED TEAS|0.09|3|TURKEY HILL P&C LEMONADE|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00020735094280|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.780702|80.78070323080172|258|1
35.318911|8cbc9057a881386c70db5fd0a7ee75906537e558|6.99|2015-02-16 20:31:00|80.780380710856576|2|3125903235|167|35.350705649277756|0|48|9937|-80.737839|885|35.297134|NFS POP SAUV/FUME BLANC|0.0|13|YELLOW TAIL SAUV BLANC|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00031259032351|POPULAR (4-$7.99)|WINE|-80.780702|80.78070323080172|258|1
35.318911|d2d8f4cee432cac89993195e27b221ce488475a8|3.99|2014-11-14 22:42:00|80.780380710856576|2|2685106106|167|35.350705649277756|0|48|6871|-80.737839|1582|35.297134|CAT FOOD & CAT NIP|0.0|18|KOOKAMUNGA CATNIP 06106|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00026851061069|PET NEEDS|GM|-80.780702|80.78070323080172|258|1
35.318911|14561cff6b884922ef98c7b44957bc2844076149|3.99|2014-11-08 19:50:00|80.780380710856576|2|7203698196|167|35.350705649277756|0|48|275|-80.737839|45|35.297134|SUPER PREMIUM ICE CREAM|0.0|5|HTT ESPRESSO CHIP GELATO|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00072036042088|ICE CREAM|FROZEN|-80.780702|80.78070323080172|258|1
35.318911|9f10a6db5cfd687ba6ee49b835911cc538817fdd|0.79|2014-11-09 21:15:00|80.780380710856576|2|7203641055|167|35.350705649277756|0|48|257|-80.737839|39|35.297134|TOMATOES|0.12|1|HT TOMATOES DICED CHILIES|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00072036410566|VEGETABLES-CAN/JAR|G1 GROCERY|-80.780702|80.78070323080172|258|1
35.318911|a857b9fd7709d34fa88aa9113e616b1ace67c2f2|2.0|2015-03-04 13:56:00|80.780380710856576|2|5100002549|167|35.350705649277756|0|48|1221|-80.737839|275|35.297134|PASTA SC VALUE|0.0|1|PREGO SC ALFREDO|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00051000197597|PASTA SAUCES|G1 GROCERY|-80.780702|80.78070323080172|258|1
35.318911|8a59813cc705ecf23bdf82026808304e6a28a2c5|1.89|2014-12-21 22:23:00|80.780380710856576|2|5100900934|167|35.350705649277756|0|48|3939|-80.737839|1075|35.297134|SHAVING CREAM MEN-CREAM|0.4|17|BARBASOL ALOE SHAVE CREAM|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00051009002731|SHAVING NEEDS/MEN HAIR|HBC|-80.780702|80.78070323080172|258|1
35.318911|25f14a9fb1ddd36a6d0e8a653e1787d63db61a70|5.58|2015-01-07 14:16:00|80.780380710856576|2|5200032669|167|35.350705649277756|0|48|171|-80.737839|20|35.297134|ISOTONIC DRINKS|0.41|1|GATORADE LEMON-LIME|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00052000338324|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.780702|80.78070323080172|258|2
35.318911|55b20e771ba3e096fb9959b3c41c1fe1ebe2810e|3.35|2015-01-23 23:07:00|80.780380710856576|2|5000012734|167|35.350705649277756|0|48|341|-80.737839|57|35.297134|CREAMERS|0.0|3|COFFEEMATE PEPPERMINT MOCHA|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00050000886104|MILK|DAIRY|-80.780702|80.78070323080172|258|1
35.318911|f1894244fb509e1fbcda9754982bf26920c6ea65|3.39|2015-01-11 17:44:00|80.780380710856576|2|5000012734|167|35.350705649277756|0|48|341|-80.737839|57|35.297134|CREAMERS|0.89|3|COFFEEMATE PEPPERMINT MOCHA|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00050000886104|MILK|DAIRY|-80.780702|80.78070323080172|258|1
35.318911|f6a93f525c2cc9699e1b60052e7e06349e3c4b39|3.19|2015-03-04 13:58:00|80.780380710856576|2|5000062231|167|35.350705649277756|0|48|326|-80.737839|54|35.297134|COOKIES/BROWNIES-REFRIGERATED|0.0|3|NESTLE CHOC. CHIP BAR COOKIES|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00050000622313|DOUGH PRODUCTS|DAIRY|-80.780702|80.78070323080172|258|1
35.318911|de766b70d37f337b6b0d2d160db36483ae18fac0|3.19|2015-03-01 22:39:00|80.780380710856576|2|5000062231|167|35.350705649277756|0|48|326|-80.737839|54|35.297134|COOKIES/BROWNIES-REFRIGERATED|0.0|3|NESTLE CHOC. CHIP BAR COOKIES|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00050000622313|DOUGH PRODUCTS|DAIRY|-80.780702|80.78070323080172|258|1
35.318911|8270343207e6797defba0b072b40269ccfe49a29|3.19|2015-01-19 21:53:00|80.780380710856576|2|5000062231|167|35.350705649277756|0|48|326|-80.737839|54|35.297134|COOKIES/BROWNIES-REFRIGERATED|0.0|3|NESTLE CHOC. CHIP BAR COOKIES|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00050000622313|DOUGH PRODUCTS|DAIRY|-80.780702|80.78070323080172|258|1
35.318911|7fad852bf776683eb3ebdff0bb2a6d68c1a59975|3.39|2014-10-22 01:15:00|80.780380710856576|2|5000012734|167|35.350705649277756|0|48|341|-80.737839|57|35.297134|CREAMERS|0.89|3|COFFEEMATE PEPPERMINT MOCHA|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00050000886104|MILK|DAIRY|-80.780702|80.78070323080172|258|1
35.318911|874e6d3de822082cb2666e9e85f69f0afe557209|4.49|2014-12-08 00:40:00|80.780380710856576|2||167|35.350705649277756|0|48|529|-80.737839|64|35.297134|FRESH ASPARAGUS|0.7|4|GREEN  ASPARAGUS|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00204080000008|FRESH PRODUCE|PRODUCE|-80.780702|80.78070323080172|258|1
35.318911|dc93e958764f89b73fc0c0d0dbb94e2389b93931|4.03|2015-02-10 19:25:00|80.780380710856576|2||167|35.350705649277756|0|48|529|-80.737839|64|35.297134|FRESH ASPARAGUS|1.01|4|GREEN  ASPARAGUS|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00204080000008|FRESH PRODUCE|PRODUCE|-80.780702|80.78070323080172|258|1
35.318911|ff34b4f62689d5f7611f83a367e1803cd16bd87f|8.62|2014-11-26 02:59:00|80.780380710856576|2||167|35.350705649277756|0|48|529|-80.737839|64|35.297134|FRESH ASPARAGUS|1.92|4|GREEN  ASPARAGUS|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00204080000008|FRESH PRODUCE|PRODUCE|-80.780702|80.78070323080172|258|1
35.318911|0c8e05da651e85a1095527336424a06145d9d8d7|7.99|2014-10-05 10:37:00|80.780380710856576|2|7203620028|167|35.350705486783326|0|48|1435|-80.992182|19|35.103409|SHELF STABLE SPREADS|0.0|1|HT ALMOND BUTTER|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00072036200280|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.780702|80.780826610732717|88|1
35.318911|e0f870d44d86bf6ccb22721340ac9ef6277434e4|8.99|2014-10-16 19:10:00|80.780380710856576|2|8992427896|167|35.350705649277756|0|48|455|-80.737839|82|35.297134|DOMESTIC PREMIUM 12PK&>|0.0|16|YUENGLING LAGER 12PK 12OZ BTL|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00089924278962|DOMESTIC BEER|BEER|-80.780702|80.78070323080172|258|1
35.318911|a2bff884de74cbf37d6994ab3de7f1cc0c798aee|2.87|2014-12-31 21:23:00|80.780380710856576|2|8130831863|167|35.350705303080211|0|48|9935|-81.027334|885|34.977331|NFS POP CAB SAUV|0.0|13|OAK CREEK CABERNET|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00081308318639|POPULAR (4-$7.99)|WINE|-80.780702|80.78088388057958|149|1
35.318911|ed1dc0fe7064247320ddd4e77296d17dd8715d3a|9.99|2015-02-12 22:25:00|80.780380710856576|2|8992427896|167|35.350705649277756|0|48|455|-80.737839|82|35.297134|DOMESTIC PREMIUM 12PK&>|0.0|16|YUENGLING LAGER 12PK 12OZ BTL|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00089924278962|DOMESTIC BEER|BEER|-80.780702|80.78070323080172|258|1
35.318911|962335707d0d57a379d5f8eac244306fbd2e02bd|3.89|2014-10-24 00:12:00|80.780380710856576|2|7684010015|167|35.350705649277756|0|48|275|-80.737839|45|35.297134|SUPER PREMIUM ICE CREAM|0.0|5|BEN & JERRY S'MORES|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00076840101771|ICE CREAM|FROZEN|-80.780702|80.78070323080172|258|1
35.318911|6ac4fca28a0bc2fdcf1fde6cf3c078d46e94aebb|3.89|2014-12-17 23:14:00|80.780380710856576|2|7684010015|167|35.350705649277756|0|48|275|-80.737839|45|35.297134|SUPER PREMIUM ICE CREAM|0.0|5|BEN & JERRY S'MORES|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00076840101771|ICE CREAM|FROZEN|-80.780702|80.78070323080172|258|1
35.318911|1ced05e3255d78b0d837a3d085620f378b94bc98|3.79|2015-03-07 23:57:00|80.780380710856576|2|7684010015|167|35.350705649277756|0|48|275|-80.737839|45|35.297134|SUPER PREMIUM ICE CREAM|0.29|5|BEN & JERRY S'MORES|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00076840101771|ICE CREAM|FROZEN|-80.780702|80.78070323080172|258|1
35.318911|e03c7012679cc76a7093c60465af09ad10946186|3.89|2014-12-09 00:22:00|80.780380710856576|2|7684010015|167|35.350705649277756|0|48|275|-80.737839|45|35.297134|SUPER PREMIUM ICE CREAM|0.0|5|BEN & JERRY S'MORES|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00076840101771|ICE CREAM|FROZEN|-80.780702|80.78070323080172|258|1
35.318911|1a72e5afca3e85796d959d8a8b0f0782748dbf08|6.39|2014-11-04 22:51:00|80.780380710856576|2|5150072001|167|35.350705649277756|0|48|125|-80.737839|19|35.297134|PEANUT BUTTER|0.0|1|JIF EXTRA CRUNCHY PEANUT BUTTE|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00051500720028|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.780702|80.78070323080172|258|1
35.318911|bd88090f4c7cb55793f62caf6b0523f3cfd6dbdc|4.49|2014-11-05 18:27:00|80.780380710856576|2|5100012938|167|35.350705649277756|0|48|212|-80.737839|33|35.297134|CONDENSED SOUP|0.0|1|CAMP COND CHICKEN NOODLE 4PK|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00051000129383|SOUP|G1 GROCERY|-80.780702|80.78070323080172|258|1
35.318911|2a56dbaa8ed09146d33c72ee69f7ffde41b616ce|7.49|2014-10-18 00:29:00|80.780380710856576|2|76108880053|167|35.350705649277756|0|48|1941|-80.737839|465|35.297134|COLD PREP FOODS MEALS|0.0|6|CHICKEN TIKKA W/JASMINE RICE|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00761088800530|COLD PREPARED FOODS|DELI|-80.780702|80.78070323080172|258|1
35.318911|ce128d4115faca5171e5313b2353548bf6fdcabe|7.49|2014-09-30 00:06:00|80.780380710856576|2|76108880053|167|35.350705649277756|0|48|1941|-80.737839|465|35.297134|COLD PREP FOODS MEALS|0.0|6|CHICKEN TIKKA W/JASMINE RICE|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00761088800530|COLD PREPARED FOODS|DELI|-80.780702|80.78070323080172|258|1
35.318911|d441d2e3b21e4015f36f69f722fe92436dcee9c7|7.49|2014-10-30 23:44:00|80.780380710856576|2|76108880053|167|35.350705649277756|0|48|1941|-80.737839|465|35.297134|COLD PREP FOODS MEALS|0.0|6|CHICKEN TIKKA W/JASMINE RICE|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00761088800530|COLD PREPARED FOODS|DELI|-80.780702|80.78070323080172|258|1
35.318911|1f85476b58be729c3d3b320896b64b5ae8217fd6|7.49|2014-10-13 00:30:00|80.780380710856576|2|76108880053|167|35.350705649277756|0|48|1941|-80.737839|465|35.297134|COLD PREP FOODS MEALS|0.0|6|CHICKEN TIKKA W/JASMINE RICE|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00761088800530|COLD PREPARED FOODS|DELI|-80.780702|80.78070323080172|258|1
35.318911|adf10ebf2c6bf3012c13a1df2f4026f11bd58deb|7.49|2014-09-25 23:55:00|80.780380710856576|2|76108880053|167|35.350705649277756|0|48|1941|-80.737839|465|35.297134|COLD PREP FOODS MEALS|0.0|6|CHICKEN TIKKA W/JASMINE RICE|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00761088800530|COLD PREPARED FOODS|DELI|-80.780702|80.78070323080172|258|1
35.318911|01a82c3efe9dcb9748451290b4b8ead6b1457871|10.99|2015-03-04 22:03:00|80.780380710856576|2|85283210625|167|35.350705649277756|0|48|9969|-80.737839|887|35.297134|NFS-S/PREM-OTHER RED|0.0|13|CAMPO VIEJO TEMPRANILLO|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00852832106258|SUPER PREMIUM ($11-$14.99)|WINE|-80.780702|80.78070323080172|258|1
35.318911|3ab3325b2c980bad82828fe8c5ece6d3dcecc933|11.99|2015-01-04 22:28:00|80.780380710856576|2|8224228043|167|35.350705649277756|0|48|9960|-80.737839|887|35.297134|NFS-S/PREM-CAB SAUVIGNON|0.0|13|NOBLE VINES 337 CABERNET SAUV|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00082242280433|SUPER PREMIUM ($11-$14.99)|WINE|-80.780702|80.78070323080172|258|1
35.318911|b75ad049add42ce2a9a94c43fb24c550bdd348cb|11.99|2014-12-11 23:28:00|80.780380710856576|2|8224228043|167|35.350705649277756|0|48|9960|-80.737839|887|35.297134|NFS-S/PREM-CAB SAUVIGNON|0.0|13|NOBLE VINES 337 CABERNET SAUV|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00082242280433|SUPER PREMIUM ($11-$14.99)|WINE|-80.780702|80.78070323080172|258|1
35.318911|a4a016445d7221aff357fad923217ef185824693|12.99|2015-01-18 01:09:00|80.780380710856576|2|8224228043|167|35.350705649277756|0|48|9960|-80.737839|887|35.297134|NFS-S/PREM-CAB SAUVIGNON|0.0|13|NOBLE VINES 337 CABERNET SAUV|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00082242280433|SUPER PREMIUM ($11-$14.99)|WINE|-80.780702|80.78070323080172|258|1
35.318911|882c9040c745c4aaf7802cc582c7a697f90f4532|11.99|2014-12-16 21:17:00|80.780380710856576|2|8224228043|167|35.350705649277756|0|48|9960|-80.737839|887|35.297134|NFS-S/PREM-CAB SAUVIGNON|0.0|13|NOBLE VINES 337 CABERNET SAUV|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00082242280433|SUPER PREMIUM ($11-$14.99)|WINE|-80.780702|80.78070323080172|258|1
35.318911|74e1f55c5f5a598c081b99b7ff8278884800ff9c|2.87|2014-10-16 19:46:00|80.780380710856576|2|7203602031|167|35.350705649277756|0|48|387|-80.737839|65|35.297134|NFS-REMAIN CHAR/LOGS/ACC|0.0|1|HT LIGHTER FLUID CAN|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00072036020314|CHARCOAL/LOGS/ACCESSORIES|G1 GROCERY|-80.780702|80.78070323080172|258|1
35.318911|8ed85783a5ef8fb5474c67d3c1b05ae85e644794|3.49|2014-12-19 23:29:00|80.780380710856576|2|20455000000|167|35.350705649277756|0|48|542|-80.737839|64|35.297134|FRESH VEGETABLES REMAIN|0.49|4|BRUSSEL SPROUTS 1LB (RPC)|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00094922577160|FRESH PRODUCE|PRODUCE|-80.780702|80.78070323080172|258|1
35.318911|06de9326872690e008713951c8e52f81669a02c4|5.99|2014-10-12 02:12:00|80.780380710856576|2|7203695041|167|35.350705649277756|0|48|1654|-80.737839|381|35.297134|DESSERT CAKES|0.0|14|2 CT. CHOC OVERLOAD TORTE|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00072036950413|CAKES|BAKERY|-80.780702|80.78070323080172|258|1
35.318911|bc5dc56fbf1a30f4ac441af0453e2385f27a18c7|9.99|2014-10-06 18:55:00|80.780380710856576|2|3100067010|167|35.350705649277756|0|48|1280|-80.737839|48|35.297134|MULTI SERVE MEALS|4.0|5|PF CHANG ORANGE CHICKEN|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00031000670023|FROZEN MEALS|FROZEN|-80.780702|80.78070323080172|258|1
35.318911|fa63e00aa07d7a2f6319a666901527b1578b3817|9.99|2014-09-25 01:12:00|80.780380710856576|2|3100067010|167|35.350705649277756|0|48|1280|-80.737839|48|35.297134|MULTI SERVE MEALS|4.0|5|PF CHANG ORANGE CHICKEN|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00031000670023|FROZEN MEALS|FROZEN|-80.780702|80.78070323080172|258|1
35.318911|d26dc8866886becd34bfe0e379f146c8498d675d|3.99|2014-12-04 23:40:00|80.780380710856576|2|7203663995|167|35.350705649277756|0|48|342|-80.737839|57|35.297134|FRESH MILK|0.0|3|HARRIS TEETER 2% MILK|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00072036639981|MILK|DAIRY|-80.780702|80.78070323080172|258|1
35.318911|aa04431ad8673b2621d89d861080297ef8a3c330|3.99|2014-09-29 01:50:00|80.780380710856576|2|7203663995|167|35.350705649277756|0|48|342|-80.737839|57|35.297134|FRESH MILK|1.02|3|HARRIS TEETER 2% MILK|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00072036639981|MILK|DAIRY|-80.780702|80.78070323080172|258|1
35.318911|b6039867d19e3cf9bb9c135d698b9d291b8c04eb|2.79|2014-11-11 13:35:00|80.780380710856576|2|3450015179|167|35.350705649277756|0|48|312|-80.737839|51|35.297134|BUTTER|0.0|3|LOL CINNAMON SUGAR BUTTER|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00034500151184|BUTTER & MARGARINE|DAIRY|-80.780702|80.78070323080172|258|1
35.318911|8933adfe7773ef025bac1bfe7c1a411b6a56b497|7.99|2014-09-15 22:07:00|80.780380710856576|2|64786510001|167|35.350705649277756|0|48|4195|-80.737839|1200|35.297134|COUGH & COLD REMEDY-ADULT|2.0|17|(FE)(JHK)AIRBORNE REG  ORANGE|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00647865100010|COUGH/COLD/SINUS|HBC|-80.780702|80.78070323080172|258|1
35.318911|d7b020dd9916348eb359d5091ae9d03023982f3e|7.99|2014-12-28 23:05:00|80.780380710856576|2|64786510001|167|35.350705649277756|0|48|4195|-80.737839|1200|35.297134|COUGH & COLD REMEDY-ADULT|0.0|17|(FE)(JHK)AIRBORNE REG  ORANGE|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00647865100010|COUGH/COLD/SINUS|HBC|-80.780702|80.78070323080172|258|1
35.318911|7683b162d43b75cd2f9879350f1ae3fe3e383a2b|6.49|2014-11-12 17:03:00|80.780380710856576|2|7203670500|167|35.350705649277756|0|48|4186|-80.737839|1200|35.297134|ALLERGY REMEDY-ADULT|0.0|17|HT ALLERGY RELIEF CAPSULES|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00072036705006|COUGH/COLD/SINUS|HBC|-80.780702|80.78070323080172|258|1
35.318911|02df96601e56bff7552fa6cf7a092cab073179ed|1.39|2014-09-20 01:45:00|80.780380710856576|2|1254667609|167|35.350705649277756|0|48|48|-80.737839|7|35.297134|REGISTER GUM|0.0|1|TRIDENT WHITE PEPPERMINT|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00012546676090|CANDY|G1 GROCERY|-80.780702|80.78070323080172|258|1
35.318911|3febfd047adf26a5bbf7e96ff7b2e66b4ef5a67b|1.39|2015-01-04 13:45:00|80.780380710856576|2|1254667609|167|35.350705649277756|0|48|48|-80.737839|7|35.297134|REGISTER GUM|0.0|1|TRIDENT WHITE PEPPERMINT|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00012546676090|CANDY|G1 GROCERY|-80.780702|80.78070323080172|258|1
35.318911|25f755e2498d6baa3bbf015ad31a874917005cf4|2.0|2015-01-29 23:23:00|80.780380710856576|2||167|35.350705649277756|0|48|511|-80.737839|64|35.297134|FRESH AVOCADOS|0.75|4|AVOCADOS, HASS XL 36CT|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00204770000004|FRESH PRODUCE|PRODUCE|-80.780702|80.78070323080172|258|1
35.318911|440aa1af1057df52d6e362e38285f085776dc34d|21.98|2014-12-13 00:27:00|80.780380710856576|2|1820000769|167|35.350705649277756|0|48|455|-80.737839|82|35.297134|DOMESTIC PREMIUM 12PK&>|0.0|16|BUD LIGHT 12PK 12OZ BTL|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00018200007699|DOMESTIC BEER|BEER|-80.780702|80.78070323080172|258|2
35.318911|2499e175f3f3553b03b3700d4106a33dadd607d8|1.99|2014-10-25 22:50:00|80.780380710856576|2|7203676016|167|35.350705649277756|0|48|151|-80.737839|23|35.297134|DSD PASTA CORE|0.0|1|HT TRADER PASTA FETTUCCINI|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00072036760227|PASTA|G1 GROCERY|-80.780702|80.78070323080172|258|1
35.318911|0b6dada07aa1486854eeb83973bbe30310e9fbaf|14.99|2014-11-20 21:58:00|80.780380710856576|2|1820053308|167|35.350705649277756|0|48|455|-80.737839|82|35.297134|DOMESTIC PREMIUM 12PK&>|0.0|16|BUD LIGHT 18PK BOTTLES|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00018200533082|DOMESTIC BEER|BEER|-80.780702|80.78070323080172|258|1
35.318911|70634c2eee5f720c2211078f6fe86fab0b2bd8a0|14.99|2014-10-22 18:07:00|80.780380710856576|2|1820053308|167|35.350705649277756|0|48|455|-80.737839|82|35.297134|DOMESTIC PREMIUM 12PK&>|0.0|16|BUD LIGHT 18PK BOTTLES|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00018200533082|DOMESTIC BEER|BEER|-80.780702|80.78070323080172|258|1
35.318911|e1dc6f048e2a5144694222c10bc395c3e68df716|3.99|2014-09-16 22:39:00|80.780380710856576|2|7203663995|167|35.350705649277756|0|48|342|-80.737839|57|35.297134|FRESH MILK|0.0|3|HARRIS TEETER WHOLE MILK|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00072036639950|MILK|DAIRY|-80.780702|80.78070323080172|258|1
35.318911|5263c3ff3db587c9c736b268249b51bada6d2802|8.99|2014-09-16 00:09:00|80.780380710856576|2|70436120024|167|35.350705649277756|0|48|458|-80.737839|82|35.297134|CRAFT BEER|0.0|16|GREAT LAKES EDM FITZGERALD 6PK|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00704361200245|DOMESTIC BEER|BEER|-80.780702|80.78070323080172|258|1
35.318911|7275bfe7c5941b0772a509f4782bd3a6b952953b|4.19|2014-10-30 09:33:00|80.780380710856576|2|7778200276|167|35.350705649277756|0|48|361|-80.737839|105|35.297134|BREAKFAST SAUSAGE|0.85|19|JOHNSONVILLE BROWN SUGAR HONEY|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00077782013573|BREAKFAST SAUSAGE|CASE READY MEATS|-80.780702|80.78070323080172|258|1
35.318911|29ffa14de34f965aa9dfea9c02f284b74da8f613|8.99|2014-10-20 23:22:00|80.780380710856576|2|8382012393|167|35.350705649277756|0|48|459|-80.737839|83|35.297134|IMPORT BEER|0.0|16|GUINNESS STOUT 6PK 12OZ BTL|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00083820123937|IMPORT BEER|BEER|-80.780702|80.78070323080172|258|1
35.318911|b6cb30908f0e3b8ef62d4b8e706a483c472c686f|6.99|2015-01-16 23:52:00|80.780380710856576|2|8992427891|167|35.350705649277756|0|48|457|-80.737839|82|35.297134|DOMESTIC SINGLES/SIX PACKS|0.0|16|YUENGLING AMBER LG 6PK12OZ BTL|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00089924278917|DOMESTIC BEER|BEER|-80.780702|80.78070323080172|258|1
35.318911|22f42338ecc6bf7b12654be1e68b583a45f039f2|8.99|2014-11-24 22:07:00|80.780380710856576|2|8382012393|167|35.350705649277756|0|48|459|-80.737839|83|35.297134|IMPORT BEER|0.0|16|GUINNESS STOUT 6PK 12OZ BTL|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00083820123937|IMPORT BEER|BEER|-80.780702|80.78070323080172|258|1
35.318911|8c4049337b2e24b9c9e8d8ec9e623d46719b4e9d|7.99|2014-09-21 22:25:00|80.780380710856576|2|2000045764|167|35.350705649277756|0|48|1280|-80.737839|48|35.297134|MULTI SERVE MEALS|0.0|5|OEP ENCHILADAS CHICKEN 6CT|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00020000457642|FROZEN MEALS|FROZEN|-80.780702|80.78070323080172|258|1
35.318911|4393c32f5b8fd67231517fc997e2b379934190b8|5.59|2014-11-27 13:16:00|80.780380710856576|2|3309200400|167|35.350705649277756|0|48|1250|-80.737839|12|35.297134|SPECIALTY COOKIES|0.6|1|HANS FREITAG DESIREE COOKIES|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00033092004007|COOKIES|G1 GROCERY|-80.780702|80.78070323080172|258|1
35.318911|3aadf8404da3889cea5d08afe3415b19cac9e620|7.99|2014-10-28 22:51:00|80.780380710856576|2|2210000288|167|35.350705649277756|0|48|454|-80.737839|82|35.297134|DOMESTIC ECONOMY 12PK&>|0.0|16|PABST 12PK 12OZ BTL|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00022100002883|DOMESTIC BEER|BEER|-80.780702|80.78070323080172|258|1
35.318911|ac314dfe2bcab269027d43efc9f4eb60376f1523|8.29|2014-10-15 23:56:00|80.780380710856576|2|2066200512|167|35.350705649277756|0|48|1280|-80.737839|48|35.297134|MULTI SERVE MEALS|1.3|5|NEWMANS ORANGE CHICKEN|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00020662005168|FROZEN MEALS|FROZEN|-80.780702|80.78070323080172|258|1
35.318911|eac382abcd36fc452f4f95a0814bd67924a11e95|0.77|2014-09-20 23:33:00|80.780380710856576|2||167|35.350705649277756|0|48|502|-80.737839|64|35.297134|FRESH BANANAS|0.0|4|BANANAS, YELLOW|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00204011000008|FRESH PRODUCE|PRODUCE|-80.780702|80.78070323080172|258|1
35.318911|8e74e729e09bee63cd038dc0a0e0a7950b9345cd|3.25|2014-11-27 13:23:00|80.780380710856576|2|7203656080|167|35.350705649277756|0|48|333|-80.737839|52|35.297134|PARMESAN CHEESE|0.0|3|HT SHREDDED PARMESAN CHEESE|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00072036550187|CHEESE|DAIRY|-80.780702|80.78070323080172|258|1
35.318911|c86bd31eab71a96a99c02cd133807e7f7f1e98a6|1.65|2014-11-29 21:52:00|80.780380710856576|2|7203663215|167|35.350705649277756|0|48|330|-80.737839|55|35.297134|EGGS|0.0|3|HT GRADE A    JUMBO WHITE EGGS|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00072036632159|EGGS FRESH|DAIRY|-80.780702|80.78070323080172|258|1
35.318911|22b8f45b6bd50d8f52b5fa4ea067e6855f8e4de9|2.49|2014-10-20 14:36:00|80.780380710856576|2|1410008550|167|35.350705303080211|0|48|87|-81.027334|13|34.977331|CHEESE CRACKERS|1.24|1|PP PF GF FLAV BLST QUESO FIEST|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00014100040200|CRACKERS|G1 GROCERY|-80.780702|80.78088388057958|149|1
35.318911|ac0940e675dd190eab43188a67de74f09e028cc1|3.58|2015-01-03 23:45:00|80.780380710856576|2|5100002457|167|35.350705649277756|0|48|212|-80.737839|33|35.297134|CONDENSED SOUP|0.54|1|CAMP COND KIDS DOUBLE NOODLE|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00051000028280|SOUP|G1 GROCERY|-80.780702|80.78070323080172|258|2
35.318911|d5f4780ae51b3289885f442f1c2aa7b53c67c84e|3.99|2014-12-10 00:05:00|80.780380710856576|2|81829001364|167|35.350705649277756|0|48|685|-80.737839|61|35.297134|GREEK|0.49|3|CHOBANI INDULGENT 4% MINT&CHOC|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00818290013637|YOGURT|DAIRY|-80.780702|80.78070323080172|258|1
35.318911|88e0be717a187f77cb84a2cfed80225ff4949d8f|1.49|2015-01-01 14:01:00|80.780380710856576|2|3000004150|167|35.350705649277756|0|48|60|-80.737839|9|35.297134|HOT CEREAL|0.0|1|QUAKER 18 QUICK GRITS|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00030000041505|CEREAL|G1 GROCERY|-80.780702|80.78070323080172|258|1
35.318911|a253d8fa52655d158d93d50311f9c980538de9a9|23.98|2014-09-10 21:22:00|80.780380710856576|2|82471033315|167|35.350705649277756|0|48|663|-80.737839|154|35.297134|FISH FILLETS/STEAKS PKGD|6.04|12|PIER 33 VP SALMON PORTION|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00824710333155|FISH FILLETS/STEAKS|SEAFOOD|-80.780702|80.78070323080172|258|2
35.318911|4f6a5965cd5a5ea178e87bcda1bab3eff15389ae|4.99|2014-09-30 14:58:00|1.4094857484078087|2|7146426060|167|0.616431285168843|0|26|577|-80.780702|136|35.318911|OTHER MERCH FR MSC JUICE|0.0|4|BOLTHOUSE PROTEIN PLUS COFFEE|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|0.61471665291522548|00071464016289|OTHER MERCHANDISE|PRODUCE|-80.780702|1.4098892219723687|167|1
35.318911|a7f499a3476209086a0dcd988fa87fa7f39f7d01|1.0|2014-12-30 16:18:00|80.780380710856576|2|3400000031|167|35.350705649277756|0|48|47|-80.737839|7|35.297134|REGISTER BARS|0.0|1|YORK PEPPERMINT PATTIES|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00034000003303|CANDY|G1 GROCERY|-80.780702|80.78070323080172|258|1
35.318911|30519213857fc190f8759fe205ec25712029d185|12.99|2015-01-02 18:07:00|80.780380710856576|2|7199076400|167|35.350705649277756|0|48|458|-80.737839|82|35.297134|CRAFT BEER|0.0|16|GEORGE KILLIANS 12PK 12OZ BTL|65142bb50acbff925c72c3e982ade6b7cb8da651|2.196933484858633|35.351085445956379|00071990764005|DOMESTIC BEER|BEER|-80.780702|80.78070323080172|258|1
35.585842|b87efdd3928a97fa9ef0ce925c45ae433f3adbeb|1.59|2014-12-26 18:44:00|80.895431304315082|4|7800023046|99|35.766165373191292|0|10|54|-80.497332|8|35.667941|DIET|0.59|23|DIET CF  CHEERWINE 2 LTR NR|676165f2b3e1f45687bf8b5d915556e47fb38135|12.459951315393052|35.810118468028598|00070925000409|CARBONATED BEVERAGES|BEVERAGE|-80.875654|80.876228264307514|178|1
35.585842|bb0823c530d4297f1a509784c87751c864a72882|11.07|2014-12-10 19:12:00|80.895431304315082|4|7729806718|99|35.766165373191292|0|10|1277|-80.497332|279|35.667941|FROZEN SNACKS|0.0|5|NANCY'S QUICHE FLORENTINE|676165f2b3e1f45687bf8b5d915556e47fb38135|12.459951315393052|35.810118468028598|00077298067282|FROZEN SANDWICH AND SNACKS|FROZEN|-80.875654|80.876228264307514|178|3
35.323246|6e04d6e8a79627c6059ac298dcac3b6d9ca5757a|3.49|2014-10-19 21:13:00|80.945255278477163|4|88491212971|166|35.387151815317949|0|13|81|-80.764523|9|35.341927|RTE CEREAL KIDS|1.74|1|POST PEBBLES COCOA|67fb0a7556932dff7124297da6c91f530c8b4ade|4.415739782503714|35.37387923947206|00884912129512|CEREAL|G1 GROCERY|-80.945176|80.94525546950922|220|1
35.323246|754f85cdd05e0144d580c81ab6f58d7867374c16|10.709999999999999|2015-01-22 20:30:00|80.945255278477163|4|7203603100|166|35.387151825807301|0|13|757|-80.66939|3|35.28326|BAKING NUTS|0.0|1|HT WALNUT PIECES|67fb0a7556932dff7124297da6c91f530c8b4ade|4.415739782503714|35.37387923947206|00072036031006|BAKING SUPPLIES|G1 GROCERY|-80.945176|80.945241573569547|46|3
35.323246|f2fbf2376b741b755e2b3ae055b4692aa3f75a61|12.99|2014-09-27 15:38:00|80.945255278477163|4|20496000000|166|35.387151345522867|0|13|755|-81.027334|87|34.977331|NFS-BALLOONS|0.0|9|*BALLOONS|67fb0a7556932dff7124297da6c91f530c8b4ade|4.415739782503714|35.37387923947206|00204960000005|FLORAL|FLORAL|-80.945176|80.945486782007492|149|1
35.323246|de7d13dc9000a4439faeae002dc87fe66b4dbd54|2.27|2014-10-11 12:05:00|80.945255278477163|4|7203611029|166|35.387151825807301|0|13|55|-80.66939|8|35.28326|REGULAR|0.0|23|HT GRAPE 12PK|67fb0a7556932dff7124297da6c91f530c8b4ade|4.415739782503714|35.37387923947206|00072036110497|CARBONATED BEVERAGES|BEVERAGE|-80.945176|80.945241573569547|46|1
35.43259|3504df7fb96c15fb77c1c6fc3ff2dc7e9f108cb0|2.99|2014-09-15 13:31:00|1.4057311447477159|4|76026391110|202|0.6184153580092175|0|52|1439|-80.605588|274|35.43259|DRY DINNERS|0.99|1|BEAR CREEK PASTA GARLIC HERB|68bd396075d990144925865b9999699071d78777|2.868847793342135|0.6209993146566879|00760263911603|PREP FOODS DINNERS|G1 GROCERY|-80.605588|1.406832906106031|202|1
35.444064|15023c5250c72355db475d8955f0ebdaa10d3a12|7.78|2014-12-04 16:32:00|1.4102725052409182|4|5450019352|121|0.6186156170875914|0|1|359|-80.995484|101|35.444064|MEAT WIENERS|1.95|19|BALL PARK BUN SIZE MEAT FRANK|6efec0bde4fa18bda44ce99c775ce6837be83e33|2.245710274202341|0.61833652052202714|00054500193274|WIENERS|CASE READY MEATS|-80.995484|1.413637875046387|121|2
35.28326|9c284685a08c455f196ac505f8ae3fd840213f12|12.99|2014-12-21 17:35:00|1.4094857484078087|4|4179021426|46|0.6158090578372145|0|26|194|-80.66939|30|35.28326|OLIVE OIL|5.0|1|BERTOLLI EX VIRGIN OLIVE OIL|738217b8e86a4f67281233587df1e84544b62832|3.4231797194294327|0.61471665291522548|00041790214260|SHORTENING/OIL|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.17739|32a8a71c88c57e40eff71b10c138bff86d6af258|4.99|2014-10-28 11:18:00|80.801203185414451|4|7203688080|208|35.193171645283492|0|24|523|-80.78468|64|35.096737|FRESH POTATOES|2.5|4|HT YUKON GOLD 5 LB BAG|745069b5266b7b8cca50102741e4692b27a35b7e|1.0904738957015905|35.194272495053255|00072036880802|FRESH PRODUCE|PRODUCE|-80.80146|80.801474744890854|30|1
35.17739|04241f1b4ec616b91129a5cd88b825f7ffc50839|5.29|2014-09-16 11:36:00|80.801203185414451|4|5100007874|208|35.193171645283492|0|24|264|-80.78468|307|35.096737|DESSERT CAKES FROZEN|0.0|5|PEP FARM PUFF PASTRY SHEETS|745069b5266b7b8cca50102741e4692b27a35b7e|1.0904738957015905|35.194272495053255|00051000078742|DESSERTS FROZEN|FROZEN|-80.80146|80.801474744890854|30|1
35.17739|5276e9b8e04bbd6b3ec0fddba457b0e551dda3b3|3.99|2014-12-02 12:31:00|80.801203185414451|4|7203663995|208|35.193171645283492|0|24|342|-80.78468|57|35.096737|FRESH MILK|1.52|3|HARRIS TEETER 2% MILK|745069b5266b7b8cca50102741e4692b27a35b7e|1.0904738957015905|35.194272495053255|00072036639981|MILK|DAIRY|-80.80146|80.801474744890854|30|1
35.17739|942a8ee9741ea6905bae1784e58e813542e68b50|1.79|2014-09-13 19:20:00|80.801203185414451|4|7800020345|208|35.193171645283492|0|24|55|-80.78468|8|35.096737|REGULAR|0.0|23|SCHWEPPES CLUB SODA 1 LTR|745069b5266b7b8cca50102741e4692b27a35b7e|1.0904738957015905|35.194272495053255|00078000203455|CARBONATED BEVERAGES|BEVERAGE|-80.80146|80.801474744890854|30|1
35.219587|795588562536e83ec7e1394269e04521046ad279|2.85|2015-02-06 20:26:00|80.810069425230125|4|7203604237|401|35.23738395181487|0|23|41|-80.80146|6|35.17739|BREAKFAST BARS|0.88|1|HT BAR CEREAL APPLE LF|74a9a0011d6c31d99ea4a4709f678a0d9d590c35|1.2297264906938778|35.240679762029046|00072036042385|BREAKFAST FOODS|G1 GROCERY|-80.810056|80.810064715205272|208|1
35.219587|a8f23766e52850e47bd55f13037077f53e67454b|2.85|2015-03-02 20:07:00|80.810069425230125|4|7203604237|401|35.23738395181487|0|23|41|-80.80146|6|35.17739|BREAKFAST BARS|0.88|1|HT BAR CEREAL APPLE LF|74a9a0011d6c31d99ea4a4709f678a0d9d590c35|1.2297264906938778|35.240679762029046|00072036042385|BREAKFAST FOODS|G1 GROCERY|-80.810056|80.810064715205272|208|1
35.219587|cd02e5e48143655b1b17a08d08fcea2a8b7bf8f3|2.85|2015-01-30 20:10:00|80.810069425230125|4|7203604237|401|35.23738395181487|0|23|41|-80.80146|6|35.17739|BREAKFAST BARS|0.88|1|HT BAR CEREAL APPLE LF|74a9a0011d6c31d99ea4a4709f678a0d9d590c35|1.2297264906938778|35.240679762029046|00072036042385|BREAKFAST FOODS|G1 GROCERY|-80.810056|80.810064715205272|208|1
35.219587|f0dadbc9d0062d58a7a060ce386d08f96df7b43d|1.79|2014-09-18 18:20:00|80.810069425230125|4|4850001775|401|35.237383948043764|0|23|335|-80.825175|56|35.152722|ORANGE JUICE-REGRIGERATED|0.79|3|TROPICANA PP CALCIUM 12 OZ|74a9a0011d6c31d99ea4a4709f678a0d9d590c35|1.2297264906938778|35.240679762029046|00048500017760|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.810056|80.810072646901688|160|1
35.219587|60a196f73b696b41065a3243b412ca82ec5e2930|2.79|2014-12-20 23:05:00|80.810069425230125|4|3800031120|401|35.237383949635444|0|23|44|-80.85013|6|35.175855|TOASTER PASTRIES-SHELF STABLE|0.0|1|KELL POPTART 12CT STRAWBERY|74a9a0011d6c31d99ea4a4709f678a0d9d590c35|1.2297264906938778|35.240679762029046|00038000317200|BREAKFAST FOODS|G1 GROCERY|-80.810056|80.810069864096988|218|1
35.219587|b5aa159b401307d8d94c8c9e87e0e6efd80384be|2.79|2014-12-04 19:32:00|80.810069425230125|4|3800031120|401|35.23738395181487|0|23|44|-80.80146|6|35.17739|TOASTER PASTRIES-SHELF STABLE|0.0|1|KELL POPTART 12CT STRAWBERY|74a9a0011d6c31d99ea4a4709f678a0d9d590c35|1.2297264906938778|35.240679762029046|00038000317200|BREAKFAST FOODS|G1 GROCERY|-80.810056|80.810064715205272|208|1
35.219587|119ae95fbceaa3788d7cb23727f6a657cbcfcdfe|2.19|2014-12-04 20:11:00|80.810069425230125|4|82348214040|401|35.23738395181487|0|23|1615|-80.80146|371|35.17739|LOCAL BREAD|0.0|14|NOVA BAGUETTE|74a9a0011d6c31d99ea4a4709f678a0d9d590c35|1.2297264906938778|35.240679762029046|00823482140404|BREAD|BAKERY|-80.810056|80.810064715205272|208|1
35.219587|f48efc10bc0195ae70ec2980ca2b2321106e32bd|2.99|2014-09-21 18:35:00|80.810069425230125|4|1600081341|401|35.237383949635444|0|23|8|-80.85013|2|35.175855|BROWNIE MIXES|0.99|1|BC SUP/HERSHEY ULTIMATE FUDGE|74a9a0011d6c31d99ea4a4709f678a0d9d590c35|1.2297264906938778|35.240679762029046|00016000813397|BAKING MIXES|G1 GROCERY|-80.810056|80.810069864096988|218|1
35.219587|7811da66320094baa500fc78924529f05c830a59|7.98|2014-12-24 15:40:00|80.810069425230125|4|7203618980|401|35.237383949635444|0|23|8436|-80.85013|1769|35.175855|ALKALINE AAA|5.98|18|HT AAA BATTERIES|74a9a0011d6c31d99ea4a4709f678a0d9d590c35|1.2297264906938778|35.240679762029046|00072036189813|BATTERY & FLASHLIGHT|GM|-80.810056|80.810069864096988|218|2
35.219587|ee9cd09db6e874b94039ce246a956cf23c635793|1.27|2014-12-07 18:22:00|80.810069425230125|4|7203603112|401|35.237383949635444|0|23|209|-80.85013|20|35.175855|POWDERED SOFT DRINKS|0.0|1|HT DRINK MIX PINK LEMONADE OTG|74a9a0011d6c31d99ea4a4709f678a0d9d590c35|1.2297264906938778|35.240679762029046|00072036031105|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.810056|80.810069864096988|218|1
35.219587|2ec9dd5f4600f097914f92e89327be41fa67ec1e|0.94|2014-10-12 18:25:00|80.810069425230125|4|7248600220|401|35.237383949635444|0|23|11|-80.85013|2|35.175855|MUFFIN MIXES|0.0|1|JIFFY CORN MUFFIN MIX|74a9a0011d6c31d99ea4a4709f678a0d9d590c35|1.2297264906938778|35.240679762029046|00072486002205|BAKING MIXES|G1 GROCERY|-80.810056|80.810069864096988|218|2
35.219587|80c3d6f578256a474b3183c9461c71793c7d628c|20.39|2014-09-10 10:04:00|80.810069425230125|4|3700085934|401|35.23738395181487|0|23|1206|-80.80146|67|35.17739|NFS-BOX DIAPERS|2.4|1|LUVS BIG BOX SIZE 4|74a9a0011d6c31d99ea4a4709f678a0d9d590c35|1.2297264906938778|35.240679762029046|00037000859352|DISPOSABLE DIAPERS|G1 GROCERY|-80.810056|80.810064715205272|208|1
35.219587|008ea99271044cd9274948be8aebca73121ea57f|9.99|2015-03-02 21:08:00|80.810069425230125|4|7203661033|401|35.23738395181487|0|23|666|-80.80146|145|35.17739|PACKAGED COOKED|0.0|12|HT COOKED SHRIMP RING 10OZ|74a9a0011d6c31d99ea4a4709f678a0d9d590c35|1.2297264906938778|35.240679762029046|00072036610331|SHRIMP|SEAFOOD|-80.810056|80.810064715205272|208|1
35.219587|af1abfb0893a405122553de737f206c83a0303bc|10.7|2015-01-23 18:24:00|80.810069425230125|4|5450019322|401|35.237383948043764|0|23|359|-80.825175|101|35.152722|MEAT WIENERS|2.67|19|BALL PARK WHITE TURKEY FRANKS|74a9a0011d6c31d99ea4a4709f678a0d9d590c35|1.2297264906938778|35.240679762029046|00054500100869|WIENERS|CASE READY MEATS|-80.810056|80.810072646901688|160|2
35.219587|4106b6f838a3c746ce654f0cec9308e79b9baa5b|2.65|2015-01-05 15:05:00|80.810069425230125|4|4119640471|401|35.237383947815992|0|23|1201|-80.849471|33|35.161696|RTS CANNED|0.65|1|PROG LIGHT CHICKEN NOODLE|74a9a0011d6c31d99ea4a4709f678a0d9d590c35|1.2297264906938778|35.240679762029046|00041196404821|SOUP|G1 GROCERY|-80.810056|80.81007300791066|35|1
35.219587|1b12e04d753a0cf75803d38adb47086260cdac69|2.59|2014-09-26 19:30:00|80.810069425230125|4|3620000250|401|35.23738395181487|0|23|1221|-80.80146|275|35.17739|PASTA SC VALUE|1.3|1|RAGU SC OWS TRADITIONAL|74a9a0011d6c31d99ea4a4709f678a0d9d590c35|1.2297264906938778|35.240679762029046|00036200002506|PASTA SAUCES|G1 GROCERY|-80.810056|80.810064715205272|208|1
35.219587|19425638269b30b3a9cb79fbc37e5678d2e97121|1.59|2014-09-26 17:53:00|80.810069425230125|4|7800015240|401|35.237383948043764|0|23|55|-80.825175|8|35.152722|REGULAR|0.2|23|C DRY GINGER ALE NR 20 OZ|74a9a0011d6c31d99ea4a4709f678a0d9d590c35|1.2297264906938778|35.240679762029046|00078000152401|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.810072646901688|160|1
35.219587|e125fc13780ff9f83336e0c9c657ebcb6ef5d17a|1.19|2014-09-28 18:29:00|80.810069425230125|4|4000000051|401|35.237383949635444|0|23|47|-80.85013|7|35.175855|REGISTER BARS|0.0|1|STARBURST ORIG FRUIT CHEWS|74a9a0011d6c31d99ea4a4709f678a0d9d590c35|1.2297264906938778|35.240679762029046|00040000000518|CANDY|G1 GROCERY|-80.810056|80.810069864096988|218|1
35.219587|2a56959c89136dcb17e93cb136bdb9859d33c6ff|3.5|2014-10-20 13:56:00|1.4094857484078087|4|7203698425|401|0.6146977543425921|0|26|254|-80.810056|892|35.219587|PREMIUM PIZZA|0.5|5|HT THIN CRUST SUPREME PIZZA|74a9a0011d6c31d99ea4a4709f678a0d9d590c35|1.2297264906938778|0.61471665291522548|00072036984272|FROZEN PIZZA|FROZEN|-80.810056|1.4104015459209989|401|1
35.500972|015e1d7eadb018293a71b96d363743854985bb8c|2.78|2015-02-15 20:05:00|80.8939826282094|4|2200000488|268|35.528154857117684|0|2|48|-80.861571|7|35.444615|REGISTER GUM|0.69|1|(FE)ORBIT SPEARMINT GUM 14 PC|74fa232f8842d37badbcf394aef76e80a07b2621|1.8782701108672621|35.490689277687849|00022000004840|CANDY|G1 GROCERY|-80.860108|80.860127744643364|340|2
35.103409|ed1553e3e1314528320d6f5772fed3ed21f970e7|6.98|2015-02-24 19:02:00|1.4132775322775095|4|88491212971|88|0.6126700657242101|0|58|81|-80.992182|9|35.103409|RTE CEREAL KIDS|1.75|1|POST PEBBLES FRUITY|79142e600cc43ddffb2448c84e274dade95cfa0d|0.8414931495528609|0.61177642288969325|00884912129710|CEREAL|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|a97b533f978332a2027afc9403b7adb95315a0db|5.69|2015-03-05 18:32:00|1.4132775322775095|4|5190001602|88|0.6126700657242101|0|58|839|-80.992182|102|35.103409|STACK PACKS|0.7|19|LOF PREMIUM HONEY TURKEY|79142e600cc43ddffb2448c84e274dade95cfa0d|0.8414931495528609|0.61177642288969325|00051900016059|LUNCHMEATS|CASE READY MEATS|-80.992182|1.413580244274486|88|1
35.103409|df6bb9d2cdb647533da1cb686cf2e0e591947c2d|2.5|2014-12-28 09:06:00|1.4132775322775095|4|7203697755|88|0.6126700657242101|0|58|81|-80.992182|9|35.103409|RTE CEREAL KIDS|0.53|1|HT CER FROSTED FLAKES|79142e600cc43ddffb2448c84e274dade95cfa0d|0.8414931495528609|0.61177642288969325|00072036977557|CEREAL|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|205207d83057f541e845152010971bf31a610f93|2.89|2014-12-06 06:51:00|1.4132775322775095|4|7203697887|88|0.6126700657242101|0|58|61|-80.992182|9|35.103409|RTE CEREAL ADULT|0.92|1|HT CER CRUNCH GRAN RAISIN BRAN|79142e600cc43ddffb2448c84e274dade95cfa0d|0.8414931495528609|0.61177642288969325|00072036978899|CEREAL|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|c22530e959b6200ae49af1eb877fa8f1c55a26c7|5.29|2014-12-16 15:18:00|1.4132775322775095|4|5150024177|88|0.6126700657242101|0|58|125|-80.992182|19|35.103409|PEANUT BUTTER|1.3|1|JIF CREAMY PEANUT BUTTER|79142e600cc43ddffb2448c84e274dade95cfa0d|0.8414931495528609|0.61177642288969325|00051500241776|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|d9cf655f5516fc0a7be6a74f3c8f51a0a4d71d16|8.7|2014-10-24 11:37:00|1.4132775322775095|4|4400002747|88|0.6126700657242101|0|58|91|-80.992182|13|35.103409|SPRAYED BUTTER CRACKERS|2.17|1|RITZ HONEY WHEAT|79142e600cc43ddffb2448c84e274dade95cfa0d|0.8414931495528609|0.61177642288969325|00044000031169|CRACKERS|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|cb1a6905355cd9f3288acd5de0e58e437bad52c7|10.99|2015-02-14 09:01:00|1.4132775322775095|4|20499400000|88|0.6126700657242101|0|58|755|-80.992182|87|35.103409|NFS-BALLOONS|2.0|9|"*AD - 36"" Jumbo Balloon"|79142e600cc43ddffb2448c84e274dade95cfa0d|0.8414931495528609|0.61177642288969325|00204994000002|FLORAL|FLORAL|-80.992182|1.413580244274486|88|1
35.103409|dfd43b6681c83c745d756119676ea183217f3a0b|6.78|2015-01-30 15:35:00|1.4132775322775095|4|4330130577|88|0.6126700657242101|0|58|1469|-80.992182|278|35.103409|REGULAR CUT FRIES|1.7|5|CHECKER'S FAMOUS FRIES|79142e600cc43ddffb2448c84e274dade95cfa0d|0.8414931495528609|0.61177642288969325|00043301305818|FROZEN POTATO|FROZEN|-80.992182|1.413580244274486|88|2
35.103409|a215056d212706d605d95ef6a837214c08395352|3.75|2014-09-27 08:26:00|1.4132775322775095|4|7433610102|88|0.6126700657242101|0|58|342|-80.992182|57|35.103409|FRESH MILK|0.0|3|HIGHLAND CREST WHOLE MILK|79142e600cc43ddffb2448c84e274dade95cfa0d|0.8414931495528609|0.61177642288969325|00074336879203|MILK|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|9f32dbaabeac155fd0bfc091503178d229ebc831|3.18|2014-10-18 13:27:00|1.4132775322775095|4|78533176189|88|0.6126700657242101|0|58|359|-80.992182|101|35.103409|MEAT WIENERS|0.62|19|GWALTNEY GREAT DOGS|79142e600cc43ddffb2448c84e274dade95cfa0d|0.8414931495528609|0.61177642288969325|00785331761898|WIENERS|CASE READY MEATS|-80.992182|1.413580244274486|88|2
35.103409|af2270404a90aae6d690230b6db53045db0cb4ed|6.98|2015-01-20 15:43:00|1.4132775322775095|4|7203660027|88|0.6126700657242101|0|58|361|-80.992182|105|35.103409|BREAKFAST SAUSAGE|0.49|19|HT BREAKFAST LINKS MAPLE|79142e600cc43ddffb2448c84e274dade95cfa0d|0.8414931495528609|0.61177642288969325|00072036600301|BREAKFAST SAUSAGE|CASE READY MEATS|-80.992182|1.413580244274486|88|2
35.103409|bdbcd52663f9162f1be6322fb4d049d2dd3ceb92|6.49|2015-02-14 09:06:00|1.4132775322775095|4|81483201002|88|0.6126700657242101|0|58|4010|-80.992182|1080|35.103409|DENTURE CLEANER PRODUCT|0.0|17|EFFERDENT DENTURE TAB NB|79142e600cc43ddffb2448c84e274dade95cfa0d|0.8414931495528609|0.61177642288969325|00814832010027|ORAL HYGIENE|HBC|-80.992182|1.413580244274486|88|1
35.103409|1a90608c542475fd73eeb634aca8efba84d60013|5.69|2014-12-31 20:54:00|1.4132775322775095|4|7203663043|88|0.6126700657242101|0|58|974|-80.992182|201|35.103409|FRESH TURKEY|0.0|2|HT 85% LEAN GROUND TURKEY|79142e600cc43ddffb2448c84e274dade95cfa0d|0.8414931495528609|0.61177642288969325|00072036630438|POULTRY|MEAT|-80.992182|1.413580244274486|88|1
35.053394|fd08011bb99abcde7de1a1164dc5bdb55510d0c3|6.99|2014-12-31 21:03:00|80.848351720559364|4|7203695205|11|35.096368251988459|0|25|1673|-80.850065|383|35.030252|PASTRY CASE CAKES|4.0|14|FFM PUMPKIN CAKE ROLL|7f4d0cec8b70fda386e7fef54e4ca8ddb6bcfdb1|2.9694171245934355|35.082633588753836|00072036952059|PASTRY CASE|BAKERY|-80.848528|80.848541020953135|470|1
35.053394|78325658f89417ca782f09530a84331cadc1c78c|2.99|2014-12-07 16:57:00|80.848351720559364|4|3338365583|11|35.096368251988459|0|25|522|-80.850065|64|35.030252|FRESH TOMATOES|0.2|4|SWEET GRAPE TOMATO (PINT)|7f4d0cec8b70fda386e7fef54e4ca8ddb6bcfdb1|2.9694171245934355|35.082633588753836|00072036880284|FRESH PRODUCE|PRODUCE|-80.848528|80.848541020953135|470|1
35.053394|09c1fd98f3ae90bb6b431031021302cd1dd43673|1.85|2014-09-17 18:35:00|80.848351720559364|4|7203663157|11|35.096368251988459|0|25|1134|-80.850065|57|35.030252|CARTON MILK|0.0|3|HARRIS TEETER WHOLE MILK|7f4d0cec8b70fda386e7fef54e4ca8ddb6bcfdb1|2.9694171245934355|35.082633588753836|00072036631572|MILK|DAIRY|-80.848528|80.848541020953135|470|1
35.053394|c7efb3287d7f1ae19f9b7c6cc4c825f3cf158254|1.85|2014-10-01 21:04:00|80.848351720559364|4|7203663157|11|35.096368251988459|0|25|1134|-80.850065|57|35.030252|CARTON MILK|0.0|3|HARRIS TEETER WHOLE MILK|7f4d0cec8b70fda386e7fef54e4ca8ddb6bcfdb1|2.9694171245934355|35.082633588753836|00072036631572|MILK|DAIRY|-80.848528|80.848541020953135|470|1
35.053394|f22078336324aad26f56b9f817888d2212eabc25|2.89|2014-12-02 21:00:00|80.848351720559364|4|7203663102|11|35.096368251988459|0|25|339|-80.850065|57|35.030252|EGGNOGS/DRINKS|0.39|3|I/O HARRIS TEETER EGG NOG|7f4d0cec8b70fda386e7fef54e4ca8ddb6bcfdb1|2.9694171245934355|35.082633588753836|00072036631022|MILK|DAIRY|-80.848528|80.848541020953135|470|1
35.053394|a2d18fe4beb5702a725e6287af181bdc0bea7d68|2.46|2014-11-07 18:12:00|80.848351720559364|4|20895100000|11|35.096368251988459|0|25|977|-80.850065|201|35.030252|FRESH HT CHICKEN|0.0|2|HT FRESH CHICKEN THIGHS|7f4d0cec8b70fda386e7fef54e4ca8ddb6bcfdb1|2.9694171245934355|35.082633588753836|00208951000005|POULTRY|MEAT|-80.848528|80.848541020953135|470|1
35.053394|b3f1ec08fc7e131c5d5773c20369d6f87687a3eb|3.19|2015-01-23 17:36:00|80.848351720559364|4|76352830603|11|35.096368252333768|0|25|1134|-80.816172|57|35.059823|CARTON MILK|0.0|3|PROMISED LAND CHOCOLATE MILK|7f4d0cec8b70fda386e7fef54e4ca8ddb6bcfdb1|2.9694171245934355|35.082633588753836|00763528306039|MILK|DAIRY|-80.848528|80.848539190811451|66|1
35.053394|a4e4bb0a81e67d60b0b6cd0ae9a4809c773578f5|3.49|2014-11-19 19:22:00|80.848351720559364|4|85225100001|11|35.096368251988459|0|25|339|-80.850065|57|35.030252|EGGNOGS/DRINKS|0.5|3|I/O SUTHRN COMF EGG NOG|7f4d0cec8b70fda386e7fef54e4ca8ddb6bcfdb1|2.9694171245934355|35.082633588753836|00852251000014|MILK|DAIRY|-80.848528|80.848541020953135|470|1
35.053394|64bc2e280a824b7b5298eee9a5a9331e009d7614|3.69|2014-10-18 17:03:00|80.848351720559364|4|7332103401|11|35.096368251425048|0|25|1277|-80.847383|279|35.024464|FROZEN SNACKS|0.79|5|SP PRETZEL SOFTSTIX BUFFALO|7f4d0cec8b70fda386e7fef54e4ca8ddb6bcfdb1|2.9694171245934355|35.082633588753836|00073321073282|FROZEN SANDWICH AND SNACKS|FROZEN|-80.848528|80.848543551325875|317|1
35.053394|2980c1f9a12c42d1558366fb854f3c6ed386749b|4.99|2015-01-17 20:10:00|1.4091206135396188|4|7336070341|11|0.6117971392988252|0|47|30|-80.848528|4|35.053394|CARBONATED WATER|1.49|1|LACROIX WTR BERRY 12PK|7f4d0cec8b70fda386e7fef54e4ca8ddb6bcfdb1|2.9694171245934355|0.61242566243833529|00073360743412|BOTTLED WATER|G1 GROCERY|-80.848528|1.411073008990826|11|1
35.053394|9be7f4c7fe9f635e29f61a8971e2137640d6c6c9|0.87|2015-02-21 18:46:00|80.848351720559364|4|7203610114|11|35.096368251425048|0|25|55|-80.847383|8|35.024464|REGULAR|0.0|23|HT GRAPE 2 LITER|7f4d0cec8b70fda386e7fef54e4ca8ddb6bcfdb1|2.9694171245934355|35.082633588753836|00072036110244|CARBONATED BEVERAGES|BEVERAGE|-80.848528|80.848543551325875|317|1
35.053394|e75f95e7c3266c2b6b029f44add7416878c0a3d8|1.49|2015-01-07 17:32:00|80.848351720559364|4|4900005537|11|35.096368251425048|0|25|54|-80.847383|8|35.024464|DIET|0.49|23|COKE ZERO 1.25 LITER BOTTLE|7f4d0cec8b70fda386e7fef54e4ca8ddb6bcfdb1|2.9694171245934355|35.082633588753836|00049000055412|CARBONATED BEVERAGES|BEVERAGE|-80.848528|80.848543551325875|317|1
35.053394|aebfad6f518a98ecd7556674aeed9a4abc457a67|2.0|2015-03-02 16:41:00|80.848351720559364|4|2840000210|11|35.096368251988459|0|25|204|-80.850065|31|35.030252|TORTILLA CHIPS|0.0|1|SANTITAS BLENDED CORN|7f4d0cec8b70fda386e7fef54e4ca8ddb6bcfdb1|2.9694171245934355|35.082633588753836|00028400002110|SNACKS|G1 GROCERY|-80.848528|80.848541020953135|470|1
35.053394|6ffe86583ac15b62d97a22c4e26ef5b586f965dc|0.87|2015-03-06 17:15:00|80.848351720559364|4|7203610114|11|35.096368251988459|0|25|55|-80.850065|8|35.030252|REGULAR|0.0|23|HT CRANBERRY GINGER AL 2 LITER|7f4d0cec8b70fda386e7fef54e4ca8ddb6bcfdb1|2.9694171245934355|35.082633588753836|00072036983916|CARBONATED BEVERAGES|BEVERAGE|-80.848528|80.848541020953135|470|1
35.053394|714149baa54cb2a958ca9aa59ea0f5ac0b4dcce7|1.99|2014-11-26 15:00:00|80.848351720559364|4|78616233800|11|35.096368251988459|0|25|31|-80.850065|4|35.030252|NON CARBONATED WATER|0.99|1|CB SMARTWATER 1 LTR PET SINGLE|7f4d0cec8b70fda386e7fef54e4ca8ddb6bcfdb1|2.9694171245934355|35.082633588753836|00786162338006|BOTTLED WATER|G1 GROCERY|-80.848528|80.848541020953135|470|1
35.053394|53f84c316ee8ce9e07d3b7257c861bc5189a5862|3.98|2014-10-03 17:46:00|80.848351720559364|4|78616233800|11|35.096368251988459|0|25|31|-80.850065|4|35.030252|NON CARBONATED WATER|1.48|1|CB SMARTWATER 1 LTR PET SINGLE|7f4d0cec8b70fda386e7fef54e4ca8ddb6bcfdb1|2.9694171245934355|35.082633588753836|00786162338006|BOTTLED WATER|G1 GROCERY|-80.848528|80.848541020953135|470|2
35.053394|fd99551ec134eef300c46f71fef77aa818a8c701|2.29|2014-10-25 17:16:00|80.848351720559364|4|63256500002|11|35.096368251425048|0|25|31|-80.847383|4|35.024464|NON CARBONATED WATER|0.62|1|CB FIJI WATER 1 LITER SINGLE|7f4d0cec8b70fda386e7fef54e4ca8ddb6bcfdb1|2.9694171245934355|35.082633588753836|00632565000029|BOTTLED WATER|G1 GROCERY|-80.848528|80.848543551325875|317|1
35.053394|1fc76e565f40b2cd0acf12d4eb449078fe9b8828|3.49|2014-10-17 18:13:00|80.848351720559364|4|7203695269|11|35.096368251425048|0|25|1895|-80.847383|450|35.024464|TEA|2.52|6|FFM GALLON LEMONADE|7f4d0cec8b70fda386e7fef54e4ca8ddb6bcfdb1|2.9694171245934355|35.082633588753836|00072036953032|BEVERAGES|DELI|-80.848528|80.848543551325875|317|1
35.053394|378c32e8e2d493ab0070391ac3c996bb80fe042f|0.99|2014-12-23 17:36:00|80.848351720559364|4|7203695306|11|35.096368177289072|0|25|1895|-80.70901|450|35.17335|TEA|0.0|6|FFM ORANGE JUICE|7f4d0cec8b70fda386e7fef54e4ca8ddb6bcfdb1|2.9694171245934355|35.082633588753836|00072036018953|BEVERAGES|DELI|-80.848528|80.848626768430819|174|1
35.318911|e69f2601a6a84d83c34b2b0344db45296ade2753|4.49|2015-03-09 20:05:00|80.779636304526477|4|1895914003|167|35.379166076554554|0|17|580|-80.737839|136|35.297134|OTHER MERCH DRESSINGS|0.0|4|PANERA CAESAR DRESSING|8252c6529f4a0189773b5a295bb4e4d7f50f1558|4.16348028119543|35.392509581117899|00018959140005|OTHER MERCHANDISE|PRODUCE|-80.780702|80.78070433335462|258|1
35.318911|fcaa85e32d68b1845e5015512280e51062a16dba|7.99|2014-11-07 18:40:00|80.779636304526477|4|85360200400|167|35.37916607363595|0|17|678|-80.764523|152|35.341927|SEAFOOD SALADS/DIPS DIPS|0.0|12|BIG T CRAB DIP|8252c6529f4a0189773b5a295bb4e4d7f50f1558|4.16348028119543|35.392509581117899|00853602004002|SALADS/DIPS|SEAFOOD|-80.780702|80.780725111286841|220|1
35.318911|8799e98b4f421e28f720d74fab1e2e7237111071|7.99|2014-11-21 17:56:00|80.779636304526477|4|85360200400|167|35.379166076554554|0|17|678|-80.737839|152|35.297134|SEAFOOD SALADS/DIPS DIPS|0.0|12|BIG T CRAB DIP|8252c6529f4a0189773b5a295bb4e4d7f50f1558|4.16348028119543|35.392509581117899|00853602004002|SALADS/DIPS|SEAFOOD|-80.780702|80.78070433335462|258|1
35.318911|c287c6f4ebdb3aac552089c7f60a63a7dbe97787|1.77|2014-10-03 18:10:00|80.779636304526477|4|4497921004|167|35.379166076584454|0|17|1469|-80.814133|278|35.333742|REGULAR CUT FRIES|0.0|5|BUYERS BEST CRINKLE CUT FRIES|8252c6529f4a0189773b5a295bb4e4d7f50f1558|4.16348028119543|35.392509581117899|00044979210046|FROZEN POTATO|FROZEN|-80.780702|80.780702164527725|472|1
35.318911|436b13681bf5d2a7586832135b3391986c9018eb|2.69|2014-10-03 18:16:00|80.779636304526477|4|5250005112|167|35.379166076584454|0|17|181|-80.814133|28|35.333742|SEAFOOD SAUCES|0.0|1|DUKES TARTAR SC SQZ|8252c6529f4a0189773b5a295bb4e4d7f50f1558|4.16348028119543|35.392509581117899|00052500051129|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.780702|80.780702164527725|472|1
35.318911|195592ae12383878b4ebdde1e047e8b58bf5a44e|5.49|2014-11-13 06:46:00|80.779636304526477|4|5100018866|167|35.379166076031403|0|17|137|-80.66939|20|35.28326|TOMATO & VEGETABLE JUICE|0.5|1|V8 FUSION+ENERGY PEACH MANGO|8252c6529f4a0189773b5a295bb4e4d7f50f1558|4.16348028119543|35.392509581117899|00051000196255|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.780702|80.780712010476662|46|1
35.318911|d3e95303cf2e89bdbce54db28ad704748bef94ab|10.19|2014-09-26 16:33:00|80.779636304526477|4|20829200000|167|35.379166076584454|0|17|660|-80.814133|154|35.333742|FISH FILLETS WILD CGHT|1.02|12|WC FRESH HADDOCK FILLETS (NO)|8252c6529f4a0189773b5a295bb4e4d7f50f1558|4.16348028119543|35.392509581117899|00208292000009|FISH FILLETS/STEAKS|SEAFOOD|-80.780702|80.780702164527725|472|1
35.318911|52eef01e259c97ea08336b64e42256ca55af9f6e|1.66|2014-10-13 21:20:00|80.779636304526477|4|4280011400|167|35.379166076584454|0|17|255|-80.814133|892|35.333742|VALUE PIZZA|0.41|5|TOTINO'S CHEESE PIZZA|8252c6529f4a0189773b5a295bb4e4d7f50f1558|4.16348028119543|35.392509581117899|00042800113009|FROZEN PIZZA|FROZEN|-80.780702|80.780702164527725|472|1
35.318911|b304814d5e4a9de637d0d13eb7ca733773f00e15|2.99|2015-03-09 20:06:00|80.779636304526477|4|5250006714|167|35.379166076554554|0|17|182|-80.737839|28|35.297134|MAYO|0.0|1|DUKES MAYO 11.5 SQZ|8252c6529f4a0189773b5a295bb4e4d7f50f1558|4.16348028119543|35.392509581117899|00052500067144|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.780702|80.78070433335462|258|1
35.318911|8c96173d0bc7e6d980d7e15b3a702bc778f2733e|1.65|2014-09-21 17:59:00|80.779636304526477|4|7203663215|167|35.379166076584454|0|17|330|-80.814133|55|35.333742|EGGS|0.0|3|HT GRADE A    JUMBO WHITE EGGS|8252c6529f4a0189773b5a295bb4e4d7f50f1558|4.16348028119543|35.392509581117899|00072036632159|EGGS FRESH|DAIRY|-80.780702|80.780702164527725|472|1
35.318911|a6e2c840ffbc947584b290b88467e701a4fb51bd|2.85|2014-11-12 18:40:00|80.779636304526477|4|4133500053|167|35.379166076031403|0|17|184|-80.66939|28|35.28326|SALAD DRESSINGS-LIQUID|0.0|1|KENS DRS CAESAR CREAMY|8252c6529f4a0189773b5a295bb4e4d7f50f1558|4.16348028119543|35.392509581117899|00041335001768|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.780702|80.780712010476662|46|1
35.318911|e48bcfbd08c962d369d647bc03941a910d321c33|7.99|2014-11-21 18:52:00|80.779636304526477|4|85360200400|167|35.379166076554554|0|17|678|-80.737839|152|35.297134|SEAFOOD SALADS/DIPS DIPS|0.0|12|BIG T SHRIMP DIP|8252c6529f4a0189773b5a295bb4e4d7f50f1558|4.16348028119543|35.392509581117899|00853602004040|SALADS/DIPS|SEAFOOD|-80.780702|80.78070433335462|258|1
35.318911|47fd87a155f652fe2d5b536e7df28a2a81ccb174|1.97|2015-03-09 20:11:00|80.779636304526477|4|2410010523|167|35.379166076554554|0|17|1252|-80.737839|12|35.297134|LUNCH BOX COOKIES|0.0|1|SUNSHINE CHEEZT IT RED FAT CDY|8252c6529f4a0189773b5a295bb4e4d7f50f1558|4.16348028119543|35.392509581117899|00024100940196|COOKIES|G1 GROCERY|-80.780702|80.78070433335462|258|1
35.318911|daff6984961a07cd0180c9f45e04c0ec01bb35af|4.29|2014-11-13 19:48:00|80.779636304526477|4|2840016014|167|35.379166076031403|0|17|201|-80.66939|31|35.28326|POTATO CHIPS|0.29|1|LAYS WAVY LIGHTLY SALTED|8252c6529f4a0189773b5a295bb4e4d7f50f1558|4.16348028119543|35.392509581117899|00028400160124|SNACKS|G1 GROCERY|-80.780702|80.780712010476662|46|1
35.318911|b8062aa096e5f594ddcafd330bfa5dcca865babb|5.99|2014-11-08 20:07:00|80.779636304526477|4|7203663044|167|35.379166076031403|0|17|974|-80.66939|201|35.28326|FRESH TURKEY|0.0|2|HT 93% LEAN GROUND TURKEY|8252c6529f4a0189773b5a295bb4e4d7f50f1558|4.16348028119543|35.392509581117899|00072036630445|POULTRY|MEAT|-80.780702|80.780712010476662|46|1
35.318911|b2ef5cf2c4cdb28eea0b68e1519e502ae4e0511b|7.99|2014-09-20 19:51:00|80.779636304526477|4|3040021526|167|35.379166076584454|0|17|426|-80.814133|72|35.333742|NFS-PAPER TOWELS|2.0|1|SPARKLE 8 RL REGULAR PRINT|8252c6529f4a0189773b5a295bb4e4d7f50f1558|4.16348028119543|35.392509581117899|00030400216503|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.780702|80.780702164527725|472|1
35.585842|6b9a53dc5722333b0c98ee2f444ea33ea83989a2|14.38|2014-11-01 11:56:00|1.4102725052409182|4|7080004118|99|0.6210901099944839|0|1|358|-80.875654|100|35.585842|REGULAR BACON|3.6|19|SMITHFIELD THICK SLC BACON|8554faa7d156520dbcd84ac0b232c92a3545f7e4|2.701560123183571|0.61833652052202714|00070800041251|BACON|CASE READY MEATS|-80.875654|1.411546447003722|99|2
35.585842|116d7fd88148a22d474346219c0453e2341522fc|1.87|2014-12-20 14:52:00|1.4102725052409182|4|7203688081|99|0.6210901099944839|0|1|524|-80.875654|64|35.585842|FRESH PROD FRESH ONIONS|0.0|4|YELLOW ONIONS 3LB BAG|8554faa7d156520dbcd84ac0b232c92a3545f7e4|2.701560123183571|0.61833652052202714|00033383600024|FRESH PRODUCE|PRODUCE|-80.875654|1.411546447003722|99|1
35.006282|14265cfdc758c1245055389ffa5a0496a92fb35b|5.99|2015-01-09 10:41:00|80.562862110758871|2|7261345844|60|35.062278583226735|0|21|1513|-80.7007|66|35.06858|NFS-LAUNDRY DETERGENT PODS|3.0|1|ALL PACS FREE&CLR 24CT|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|35.054042368968126|00072613458448|DETERGENTS|G1 GROCERY|-80.562829|80.562830704304375|273|1
35.006282|18d3e5d23bbf259a247690e17f2b52b1a9af5ed3|4.69|2015-01-10 12:32:00|80.562862110758871|2|7261345111|60|35.062278583226735|0|21|417|-80.7007|71|35.06858|NFS-FABRIC SOFTENERS|1.69|1|SNUGGLE SPARKLE SHEETS 80CT|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|35.054042368968126|00072613451111|LAUNDRY SUPPLIES|G1 GROCERY|-80.562829|80.562830704304375|273|1
35.006282|d4fdc3e3499c083fa17425307512210fdb593463|3.09|2015-01-17 17:55:00|1.4091206135396188|2|20328700000|60|0.6109748797816256|0|47|641|-80.562829|137|35.006282|PREMIUM PORK|0.0|2|PORK LOIN RIB END CHOPS BNLS|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|0.61242566243833529|00203287000002|PORK|MEAT|-80.562829|1.4060866207711706|60|1
35.006282|d4db1eaa7d99442a8c9338e7974b9319afe6708f|2.19|2014-11-08 17:47:00|1.4091206135396188|2|7203698771|60|0.6109748797816256|0|47|176|-80.562829|72|35.006282|NFS-DISPOSE CUPS|0.4|1|YH FOAM CUPS 10 OZ|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|0.61242566243833529|00072036987716|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.562829|1.4060866207711706|60|1
35.006282|3fb451a09cfa4cf2a0b4a9cc2e599358de6f00ec|3.5999999999999996|2014-12-14 18:03:00|80.562862110758871|2|89470001004|60|35.062278547561078|0|21|685|-80.62331|61|35.140781|GREEK|0.6000000000000001|3|CHOBANI SEASONAL GREEN TEA|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|35.054042368968126|00818290013866|YOGURT|DAIRY|-80.562829|80.562906204784099|39|3
35.006282|b761d36a6b6adf6bb22955fa978695ad8c8d1ec0|20.759999999999998|2014-11-16 13:38:00|1.4091206135396188|2|20895300000|60|0.6109748797816256|0|47|977|-80.562829|201|35.006282|FRESH HT CHICKEN|5.26|2|HT FRESH BNLS CHICKEN BREAST|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|0.61242566243833529|00208953000003|POULTRY|MEAT|-80.562829|1.4060866207711706|60|2
35.006282|58d377c922ff6a0008cbeeeba56f3bc166457eac|3.39|2014-09-20 14:49:00|80.562862110758871|2|60502100099|60|35.062278564801773|0|21|1246|-80.654118|34|35.123768|SPICE BLENDS|0.4|1|MRS DASH TABLE BLEND|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|35.054042368968126|00605021000994|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.562829|80.562884503636255|473|1
35.006282|be64486e45a5a8d437a403c7b5d4692fc1b2628e|2.99|2015-02-19 17:21:00|1.4091206135396188|2|70601011292|60|0.6109748797816256|0|47|1219|-80.562829|275|35.006282|PASTA SC CORE|0.99|1|BARILLA SC MARINARA|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|0.61242566243833529|00706010112923|PASTA SAUCES|G1 GROCERY|-80.562829|1.4060866207711706|60|1
35.006282|b57c5322ca8ac9684550bfbc8b22800386827849|8.38|2014-10-17 10:54:00|80.562862110758871|2|31015805306|60|35.062278583226735|0|21|4010|-80.7007|1080|35.06858|DENTURE CLEANER PRODUCT|0.0|17|POLIDENT 3 MINUTE TABS NB|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|35.054042368968126|00310158053064|ORAL HYGIENE|HBC|-80.562829|80.562830704304375|273|2
35.006282|04e948bd4c52b0d59abed46cdd79f2b2adb7e92a|8.38|2015-01-07 12:07:00|80.562862110758871|2|31015805306|60|35.062278583226735|0|21|4010|-80.7007|1080|35.06858|DENTURE CLEANER PRODUCT|0.0|17|POLIDENT 3 MINUTE TABS NB|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|35.054042368968126|00310158053064|ORAL HYGIENE|HBC|-80.562829|80.562830704304375|273|2
35.006282|56ebf78d792eacec0ed97d9b3526740b3f4a3f95|3.5999999999999996|2014-10-05 14:41:00|80.562862110758871|2|68954408130|60|35.062278583201362|0|21|685|-80.64817|61|35.04711|GREEK|0.0|3|FAGE 0% WITH HONEY|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|35.054042368968126|00689544081258|YOGURT|DAIRY|-80.562829|80.562831672536859|129|3
35.006282|8ff5abe9744d4b134346ae2360b342fc0a9cf603|1.49|2014-09-18 17:45:00|80.562862110758871|2||60|35.062278564801773|0|21|561|-80.654118|64|35.123768|FR PROD ORGANIC PRODUCE|0.0|4|COO ORG CUCUMBERS|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|35.054042368968126|00294062000003|FRESH PRODUCE|PRODUCE|-80.562829|80.562884503636255|473|1
35.006282|2872807bf216c047f9a7ccbf9f0a0559f162cf73|3.69|2014-10-28 20:01:00|1.4091206135396188|2|2059300015|60|0.6109748797816256|0|47|1459|-80.562829|40|35.006282|FROZEN BISCUITS|0.0|5|MARY B'S SOUTHERN MADE BISCUIT|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|0.61242566243833529|00020593000188|FROZEN DOUGH|FROZEN|-80.562829|1.4060866207711706|60|1
35.006282|5aa395c0a6d6ccbfedd913dfe61aa4cf26de535b|1.27|2014-12-24 16:22:00|1.4091206135396188|2|5963500189|60|0.6109748797816256|0|47|1461|-80.562829|40|35.006282|FROZEN GARLIC TOAST AND BRD|0.0|5|FURLANI TEXAS TOAST|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|0.61242566243833529|00059635001890|FROZEN DOUGH|FROZEN|-80.562829|1.4060866207711706|60|1
35.006282|d5d22b0ba11ad0d493547d8efa638372e4880510|0.45|2014-11-30 17:34:00|1.4091206135396188|2||60|0.6109748797816256|0|47|522|-80.562829|64|35.006282|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|0.61242566243833529|00204664000004|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|1
35.006282|ce209bdf0769dcdffe8dd7e6d25ef8fcfef775a4|4.49|2014-10-15 11:10:00|80.562862110758871|2|30521309100|60|35.062278564801773|0|21|3200|-80.654118|1015|35.123768|HAND & BODY EXPERIENTIAL|1.0|17|VICL MEN LTN BODY/FACE X-STR|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|35.054042368968126|00305210416390|HAND & BODY LOTION/SUN CARE|HBC|-80.562829|80.562884503636255|473|1
35.006282|55b41ac69044006e167f78b36de77c6a5289dba1|4.19|2015-01-08 11:16:00|80.562862110758871|2|38137003016|60|35.062278583226735|0|21|5189|-80.7007|1305|35.06858|BABY POWDER|1.69|17|J&J BABY POWDER LAVENDER 03017|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|35.054042368968126|00381370030171|BABY HBC|HBC|-80.562829|80.562830704304375|273|1
35.006282|2aeef16a4a93528f9732ad6d0afd2e78820c0216|1.95|2015-01-03 15:40:00|1.4091206135396188|2|1450001098|60|0.6109748797816256|0|47|1272|-80.562829|50|35.006282|BAG VEG STEAM|0.0|5|BE STEAMFRESH WHL GRN BRN RICE|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|0.61242566243833529|00014500012807|VEGETABLES-FROZEN|FROZEN|-80.562829|1.4060866207711706|60|1
35.006282|dc1be8188adb76adaecc9f66fb768bff3149202b|3.59|2015-01-25 17:12:00|1.4091206135396188|2|88491212611|60|0.6109748797816256|0|47|61|-80.562829|9|35.006282|RTE CEREAL ADULT|0.0|1|POST G GRAIN RAISIN DATE PECAN|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|0.61242566243833529|00884912126115|CEREAL|G1 GROCERY|-80.562829|1.4060866207711706|60|1
35.006282|a9bb42d7c238ca33675fd25311f653e054d8b283|3.39|2014-10-20 11:50:00|80.562862110758871|2|7550000011|60|35.062278583226735|0|21|76|-80.7007|11|35.06858|MEAT SAUCES|0.89|1|TEXAS PETE WING BUFFALO|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|35.054042368968126|00075500000119|CONDIMENTS|G1 GROCERY|-80.562829|80.562830704304375|273|1
35.006282|2fc7c71aa9dba56fa6206c536c2e6545aed633fd|2.99|2014-10-01 19:25:00|1.4091206135396188|2|7341013546|60|0.6109748797816256|0|47|1035|-80.562829|163|35.006282|SANDWICH ROLL|0.0|7|ARN HNY WHEAT SANDWICH THIN PP|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|0.61242566243833529|00073410135433|BUNS/ROLLS|COMMERCIAL BAKERY|-80.562829|1.4060866207711706|60|1
35.006282|c1bff3b4256eb970302d2b13bf37ebbeec2b0d2c|3.25|2015-02-14 16:08:00|1.4091206135396188|2|7203656080|60|0.6109748797816256|0|47|318|-80.562829|52|35.006282|SHREDDED/GRATED CHEESE|0.0|3|HT GOURMENT SHARP BLEND|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|0.61242566243833529|00072036600783|CHEESE|DAIRY|-80.562829|1.4060866207711706|60|1
35.006282|6b23d1ee078e921f8e376d86e7b6f7f728db3872|19.77|2015-01-11 13:56:00|80.562862110758871|2|3320097202|60|35.062278583226735|0|21|1513|-80.7007|66|35.06858|NFS-LAUNDRY DETERGENT PODS|3.3000000000000003|1|A&H TOSS N DONE POWR PAK|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|35.054042368968126|00033200972020|DETERGENTS|G1 GROCERY|-80.562829|80.562830704304375|273|3
35.006282|5ca562c425270412a680acea9e3d5c5adc191195|0.47|2014-10-30 16:35:00|80.562862110758871|2|7248600220|60|35.062278564801773|0|21|11|-80.654118|2|35.123768|MUFFIN MIXES|0.0|1|JIFFY CORN MUFFIN MIX|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|35.054042368968126|00072486002205|BAKING MIXES|G1 GROCERY|-80.562829|80.562884503636255|473|1
35.006282|142a6327b24a9bf6eb2bdbe52b5bf46a55cb6a7f|5.98|2015-01-13 11:09:00|80.562862110758871|2|3700012340|60|35.062278583226735|0|21|3874|-80.7007|1070|35.06858|SOLID-FEMALE|0.98|17|SECRET SOLID WS POWDER FRESH|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|35.054042368968126|00037000124511|DEODORANT|HBC|-80.562829|80.562830704304375|273|2
35.006282|d4467417d6a40020c5036ee9e6cd588c3f091eaa|6.36|2014-10-19 18:22:00|80.562862110758871|2|4650073332|60|35.062278583226735|0|21|393|-80.7007|68|35.06858|NFS-AIR FRESHENERS|2.36|1|GLADE AEROSOL LAVENDR VANILLA|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|35.054042368968126|00046500733345|FRESHENERS/DEODORIZERS|G1 GROCERY|-80.562829|80.562830704304375|273|4
35.006282|dcbdc4d82e313a7b8a8ad24706d0b6951369e8f3|4.79|2014-11-22 16:12:00|1.4091206135396188|2|1200010041|60|0.6109748797816256|0|47|54|-80.562829|8|35.006282|DIET|2.4|23|DIET MTN DEW 16 OZ 6 PK|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|0.61242566243833529|00012000107061|CARBONATED BEVERAGES|BEVERAGE|-80.562829|1.4060866207711706|60|1
35.006282|950bde89807a6e397de4277d2c76bbdcb2051dbb|4.39|2015-01-30 16:26:00|80.562862110758871|2|4400002747|60|35.062278547561078|0|21|91|-80.62331|13|35.140781|SPRAYED BUTTER CRACKERS|2.19|1|RITZ FRESH STACKS|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|35.054042368968126|00044000031138|CRACKERS|G1 GROCERY|-80.562829|80.562906204784099|39|1
35.006282|b24fc648e98348231d15b83e3cb8b6b2f961e3e5|4.0|2014-11-23 13:31:00|1.4091206135396188|2|7726006180|60|0.6109748797816256|0|47|727|-80.562829|7|35.006282|SEASONAL CANDY-SINGLE FAC|1.0|1|I/O(C15)RS PPRMNT BRK BLLON BR|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|0.61242566243833529|00077260061805|CANDY|G1 GROCERY|-80.562829|1.4060866207711706|60|4
35.006282|3623a081a1df380bbf4bfddf13065ebf95b81692|2.19|2015-01-19 13:16:00|80.562862110758871|2|1200000496|60|35.062278583201362|0|21|55|-80.64817|8|35.04711|REGULAR|0.52|23|C/F PEPSI 2LTR NR|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|35.054042368968126|00012000004926|CARBONATED BEVERAGES|BEVERAGE|-80.562829|80.562831672536859|129|1
35.006282|b3da761b0aa2df115702132a57fc92baf7962ea9|6.98|2015-01-10 12:33:00|80.562862110758871|2|8087800218|60|35.062278583226735|0|21|3548|-80.7007|1045|35.06858|HAIR CARE SHPOO 2 IN 1'S|0.0|17|PANTENE SH 2N1 VOLUME|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|35.054042368968126|00080878042203|HAIR & SCALP CARE|HBC|-80.562829|80.562830704304375|273|2
35.006282|5b74aebdef4574844ca3ebfc60f1f0c8c0c7fe18|1.0|2015-02-12 16:57:00|80.562862110758871|2||60|35.062278547561078|0|21|1639|-80.62331|377|35.140781|BULK (DONUTS)|0.0|14|OLD KK BULK DONUT CODE|89291454cfc66b675261bba584e1904b0d2eb8f5|3.8692286752613088|35.054042368968126|00072470005298|DONUTS|BAKERY|-80.562829|80.562906204784099|39|1
35.323246|029717dfd39fc8cf885d3c42d0851f298a53a1c1|4.99|2014-11-02 16:56:00|1.4102725052409182|3|1111018700|166|0.6165069451919168|0|1|1647|-80.945176|379|35.323246|PACKAGED MUFFINS|2.5|14|FFM 4 CT DBL CHOC CHIP MUFFIN|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|0.61833652052202714|00011110187024|MUFFINS|BAKERY|-80.945176|1.4127598348062935|166|1
35.323246|cac548796e88c5f8dea7fcd1dd5dd8d0ce3f51e7|6.89|2014-10-14 11:38:00|80.945290274299126|3|7261345083|166|35.414868531832361|0|44|389|-80.995484|66|35.444064|NFS-LAUNDRY DETERGENTS|1.89|1|WISK ULTRA|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00072613450831|DETERGENTS|G1 GROCERY|-80.945176|80.945291222334149|121|1
35.323246|ad036109c5000a7bf924756d78e69acb77a0121f|3.75|2014-09-24 18:01:00|80.945290274299126|3|7433610102|166|35.414868531832361|0|44|342|-80.995484|57|35.444064|FRESH MILK|0.0|3|HIGHLAND CREST WHOLE MILK|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00074336879203|MILK|DAIRY|-80.945176|80.945291222334149|121|1
35.323246|a5e7c8c8d8962d971cf6d8bb5adc6bdacbb59642|0.97|2014-11-22 16:42:00|1.4102725052409182|3|7203688002|166|0.6165069451919168|0|1|527|-80.945176|64|35.323246|FRESH CARROTS|0.0|4|HT WHOLE CARROTS 2LB BAG|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|0.61833652052202714|00072036880024|FRESH PRODUCE|PRODUCE|-80.945176|1.4127598348062935|166|1
35.323246|c3aea333d697a5f9d7d55a458aaedb10693929fe|5.29|2014-09-28 16:30:00|1.4102725052409182|3|7203651143|166|0.6165069451919168|0|1|252|-80.945176|45|35.323246|PREMIUM ICE CREAM|2.29|5|HT ALL NATURAL TRPL CHOCOLATE|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|0.61833652052202714|00072036980113|ICE CREAM|FROZEN|-80.945176|1.4127598348062935|166|1
35.323246|83c471e3d290a5dda74d4dec9b9b0fe4c6bb6973|5.29|2014-10-28 19:14:00|1.4102725052409182|3|7203651143|166|0.6165069451919168|0|1|252|-80.945176|45|35.323246|PREMIUM ICE CREAM|0.0|5|HT ALL NATURAL TRPL CHOCOLATE|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|0.61833652052202714|00072036980113|ICE CREAM|FROZEN|-80.945176|1.4127598348062935|166|1
35.323246|e5c62f7d98bf4232e290bf58acc07a081715a5e1|5.29|2015-01-27 18:53:00|80.945290274299126|3|7203651143|166|35.414868531832361|0|44|252|-80.995484|45|35.444064|PREMIUM ICE CREAM|5.29|5|HT ALL NATURAL TRPL CHOCOLATE|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00072036980113|ICE CREAM|FROZEN|-80.945176|80.945291222334149|121|1
35.323246|2e95e04aa035b6df472fe8864ff5ff990b5ed5f9|5.98|2014-12-13 15:14:00|1.4102725052409182|3|64420933250|166|0.6165069451919168|0|1|8|-80.945176|2|35.323246|BROWNIE MIXES|0.98|1|D HINES MILK CHOC BROWNIE MIX|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|0.61833652052202714|00644209332496|BAKING MIXES|G1 GROCERY|-80.945176|1.4127598348062935|166|2
35.323246|8901d60f527989ba195619c30209037550009d5e|2.99|2015-02-26 18:05:00|1.4102725052409182|3|64420933250|166|0.6165069451919168|0|1|8|-80.945176|2|35.323246|BROWNIE MIXES|0.5|1|D HINES MILK CHOC BROWNIE MIX|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|0.61833652052202714|00644209332496|BAKING MIXES|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|a3e027783fb620915c7c467270b6bc87972c9cbf|3.99|2014-10-26 16:48:00|1.4102725052409182|3|7079660028|166|0.6165069451919168|0|1|161|-80.945176|25|35.323246|PEPPERS|0.4|1|CENTO ROASTED PEPPERS 12|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|0.61833652052202714|00070796600289|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|bda57456f817eab520f31b1b6d3ca053f973aca6|4.39|2014-11-09 16:51:00|1.4102725052409182|3|5150003357|166|0.6165069451919168|0|1|126|-80.945176|19|35.323246|PRESERVES/MARMALADE|1.4|1|DICKINSON SDLS BLACKBERRY|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|0.61833652052202714|00051500033579|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|b102b810e13d9c476cbce4f90a9f8a1478ddb746|1.69|2015-02-20 17:03:00|1.4102725052409182|3|5480005009|166|0.6165069451919168|0|1|238|-80.945176|38|35.323246|RICE FLAVORED|0.69|1|UNCLE BENS C INN CHICKEN R/V|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|0.61833652052202714|00054800050093|RICE GRAINS AND BEANS|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|7d1b8cb8725d0f101df45f33028b14b29f97e5c5|3.79|2014-12-23 17:35:00|1.4102725052409182|3|5565367020|166|0.6165069451919168|0|1|92|-80.945176|13|35.323246|REMAINING CRACKERS|0.79|1|DARE BRETON CRACKERS|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|0.61833652052202714|00055653670209|CRACKERS|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|57f8811cd4302970a740adaf08d759bd1ca325d3|9.49|2014-10-11 18:08:00|1.4102725052409182|3|5400011971|166|0.6165069451919168|0|1|427|-80.945176|72|35.323246|NFS-TOILET TISSUE|2.5|1|SCOTT 1000 WHITE 8 ROLL|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|0.61833652052202714|00054000119712|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|c08f4012bc2d252bbe96178a57852dc6c2f59efe|2.99|2014-11-19 16:28:00|80.945290274299126|3|8201110007|166|35.414868531832361|0|44|1250|-80.995484|12|35.444064|SPECIALTY COOKIES|0.99|1|MURRAY GINGER SNAPS|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00082011100078|COOKIES|G1 GROCERY|-80.945176|80.945291222334149|121|1
35.323246|7d0585477621fb168a2bb6e248764b1db6fbd986|5.98|2014-12-05 15:34:00|80.945290274299126|3|8201110007|166|35.414868531832361|0|44|1250|-80.995484|12|35.444064|SPECIALTY COOKIES|0.99|1|MURRAY GINGER SNAPS|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00082011100078|COOKIES|G1 GROCERY|-80.945176|80.945291222334149|121|2
35.323246|161aa65dea8f72045d23627061e673c72a87e21b|1.99|2014-09-10 13:31:00|80.945290274299126|3|78616233800|166|35.414868531832361|0|44|31|-80.995484|4|35.444064|NON CARBONATED WATER|0.99|1|CB SMARTWATER 1 LTR PET SINGLE|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00786162338006|BOTTLED WATER|G1 GROCERY|-80.945176|80.945291222334149|121|1
35.323246|5d1bd93a5d2ffeaef495c0b8e9a9fdd6b72d8776|5.63|2014-10-17 18:11:00|80.945290274299126|3||166|35.414868545717489|0|44|500|-80.80146|64|35.17739|FRESH APPLES|2.12|4|HONEY CRISP APPLE|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00233283000003|FRESH PRODUCE|PRODUCE|-80.945176|80.945273209668315|208|1
35.323246|4dc52478317d80e876e550652c1443abe3f8dc40|2.39|2015-02-27 17:45:00|1.4102725052409182|3|7203698241|166|0.6165069451919168|0|1|442|-80.945176|76|35.323246|NFS-COOKING-STORAGE BAGS|0.72|1|YH RESEALABLE SANDWICH BAGS|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|0.61833652052202714|00072036982414|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|a87a7e118a965964572e601f241a50d318815554|5.29|2015-01-05 17:59:00|1.4102725052409182|3|7203651143|166|0.6165069451919168|0|1|252|-80.945176|45|35.323246|PREMIUM ICE CREAM|2.65|5|HT ALL NATURAL NATURALLY VAN|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|0.61833652052202714|00072036511430|ICE CREAM|FROZEN|-80.945176|1.4127598348062935|166|1
35.323246|4865e01fce242a738c2a6438cc803c07204245c9|3.34|2014-09-16 17:37:00|1.4102725052409182|3|7203643010|166|0.6165069451919168|0|1|252|-80.945176|45|35.323246|PREMIUM ICE CREAM|0.0|5|HT PREM PEANUT BUTTER CUP IC|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|0.61833652052202714|00072036430250|ICE CREAM|FROZEN|-80.945176|1.4127598348062935|166|1
35.323246|e899ad8087531be4b2825de798f4ccae400bdd47|6.67|2014-11-14 19:09:00|80.945290274299126|3|7203643010|166|35.414868531832361|0|44|252|-80.995484|45|35.444064|PREMIUM ICE CREAM|0.0|5|HT PREM PEANUT BUTTER CUP IC|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00072036430250|ICE CREAM|FROZEN|-80.945176|80.945291222334149|121|2
35.323246|a45fbb2fdad8f5d4907633f545b728ce67054ebe|3.34|2014-10-07 19:01:00|1.4102725052409182|3|7203643010|166|0.6165069451919168|0|1|252|-80.945176|45|35.323246|PREMIUM ICE CREAM|0.84|5|HT PREM PEANUT BUTTER CUP IC|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|0.61833652052202714|00072036430250|ICE CREAM|FROZEN|-80.945176|1.4127598348062935|166|1
35.323246|726dd73f58c43cb1d6660be5aeef05e16098bf1a|3.58|2014-10-31 19:32:00|1.4102725052409182|3|5100001047|166|0.6165069451919168|0|1|212|-80.945176|33|35.323246|CONDENSED SOUP|1.58|1|CAMP COND TOMATO BISQUE|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|0.61833652052202714|00051000015877|SOUP|G1 GROCERY|-80.945176|1.4127598348062935|166|2
35.323246|88b227d51e14d346e59338117cddfde5f8285d41|3.99|2014-09-19 15:09:00|1.4102725052409182|3|4850002013|166|0.6165069451919168|0|1|335|-80.945176|56|35.323246|ORANGE JUICE-REGRIGERATED|0.99|3|TROPICANA PP HOMESTYLE|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|0.61833652052202714|00048500301395|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.945176|1.4127598348062935|166|1
35.323246|73a52117ce7a2a4b9929de495f81ecdf548753fc|1.67|2014-12-16 18:59:00|80.945290274299126|3|7203670851|166|35.414868531832361|0|44|1262|-80.995484|57|35.444064|HALF N HALF WHIPPING CREAM|0.0|3|HIGHLAND CREST HALF&HALF|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00072036708519|MILK|DAIRY|-80.945176|80.945291222334149|121|1
35.323246|78fca90f97f18d51de8b5c8c318058c42fc29f45|1.87|2015-02-11 18:31:00|1.4102725052409182|3|7203670851|166|0.6165069451919168|0|1|1262|-80.945176|57|35.323246|HALF N HALF WHIPPING CREAM|0.0|3|HIGHLAND CREST HALF&HALF|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|0.61833652052202714|00072036708519|MILK|DAIRY|-80.945176|1.4127598348062935|166|1
35.323246|fa528275ae0c1b5ffdd6c340fbab9fde16c6195b|1.67|2014-11-28 19:31:00|80.945290274299126|3|7203670851|166|35.414868531832361|0|44|1262|-80.995484|57|35.444064|HALF N HALF WHIPPING CREAM|0.0|3|HIGHLAND CREST HALF&HALF|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00072036708519|MILK|DAIRY|-80.945176|80.945291222334149|121|1
35.323246|235db8e4b8e78de92c76fb0915af04d7d2b8babc|6.98|2014-09-26 14:36:00|80.945290274299126|3|7203671181|166|35.414868531832361|0|44|252|-80.995484|45|35.444064|PREMIUM ICE CREAM|0.49|5|HT RASPBERRY SHERBET|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00072036711830|ICE CREAM|FROZEN|-80.945176|80.945291222334149|121|2
35.323246|71ea36770575bf1bf93b6ec106df6589665515e6|1.67|2014-11-18 19:53:00|80.945290274299126|3|7203670851|166|35.414868531832361|0|44|1262|-80.995484|57|35.444064|HALF N HALF WHIPPING CREAM|0.0|3|HIGHLAND CREST HALF&HALF|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00072036708519|MILK|DAIRY|-80.945176|80.945291222334149|121|1
35.323246|c52f659142913119ce26afe7e4bc2c275f531634|1.67|2014-11-19 20:18:00|80.945290274299126|3|7203670851|166|35.414868531832361|0|44|1262|-80.995484|57|35.444064|HALF N HALF WHIPPING CREAM|0.0|3|HIGHLAND CREST HALF&HALF|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00072036708519|MILK|DAIRY|-80.945176|80.945291222334149|121|1
35.323246|80f58468295752bc95d6ceadd99db15c574b8ad2|1.87|2015-01-23 10:43:00|1.4102725052409182|3|7203670851|166|0.6165069451919168|0|1|1262|-80.945176|57|35.323246|HALF N HALF WHIPPING CREAM|0.0|3|HIGHLAND CREST HALF&HALF|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|0.61833652052202714|00072036708519|MILK|DAIRY|-80.945176|1.4127598348062935|166|1
35.323246|e2a0ecf951aa50ddc0cd72baa267af660c51302e|2.29|2014-10-16 10:26:00|80.945290274299126|3|1900008501|166|35.414868531832361|0|44|50|-80.995484|7|35.444064|PEG CANDY|0.29|1|LIFESAVERS PEP-O-MINT PEG|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00019000085030|CANDY|G1 GROCERY|-80.945176|80.945291222334149|121|1
35.323246|5cc662aa959d4e41974fe810789dab2c172d7bd4|6.0|2015-01-06 18:50:00|80.945290274299126|3|7203663118|166|35.414868531832361|0|44|1262|-80.995484|57|35.444064|HALF N HALF WHIPPING CREAM|0.33|3|HT HALF & HALF|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00072036632043|MILK|DAIRY|-80.945176|80.945291222334149|121|3
35.323246|728ad0fdccc146865d413b257955a75b865f0883|3.34|2015-02-05 15:40:00|1.4102725052409182|3|7203643010|166|0.6165069451919168|0|1|252|-80.945176|45|35.323246|PREMIUM ICE CREAM|0.0|5|HT PREM TURTLE PECAN SWIRL IC|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|0.61833652052202714|00072036980144|ICE CREAM|FROZEN|-80.945176|1.4127598348062935|166|1
35.323246|cab45b7701507458813dff7acaae8336c176f23e|5.0|2014-11-01 18:05:00|80.945290274299126|3|20600200000|166|35.414868531832361|0|44|1802|-80.995484|400|35.444064|FFM HAM|2.5|6|HONEY CURED HAM|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00206002000004|FFM MEAT|DELI|-80.945176|80.945291222334149|121|1
35.323246|941179f6979c38fd6c1e26ffd67da84dc0a3ce54|1.49|2014-09-17 13:24:00|80.945290274299126|3|4900002656|166|35.414868531832361|0|44|31|-80.995484|4|35.444064|NON CARBONATED WATER|0.49|1|CB DASANI WATER  1 LITER|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00049000026566|BOTTLED WATER|G1 GROCERY|-80.945176|80.945291222334149|121|1
35.323246|987271b46950da03b43716b44dba32b7652ce9d2|3.95|2014-12-11 21:13:00|80.945290274299126|3|7203663995|166|35.414868505585332|0|44|342|-80.86175|57|35.40953|FRESH MILK|0.0|3|HARRIS TEETER WHOLE MILK|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00072036639950|MILK|DAIRY|-80.945176|80.945319210836331|209|1
35.323246|64edf0ad45267588149ed0cf613543f9a660ef95|3.49|2015-01-14 11:03:00|80.945290274299126|3|7641090137|166|35.414868531832361|0|44|1252|-80.995484|12|35.444064|LUNCH BOX COOKIES|1.75|1|LANCE NEKOT PEANUT BUTTER 8PK|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00076410901398|COOKIES|G1 GROCERY|-80.945176|80.945291222334149|121|1
35.323246|93608f6d79a05beb86027713bdb13286126097d0|1.39|2014-10-29 15:09:00|80.945290274299126|3|8265750067|166|35.414868531832361|0|44|31|-80.995484|4|35.444064|NON CARBONATED WATER|0.39|1|DEER PARK WATER 1LT|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00082657500676|BOTTLED WATER|G1 GROCERY|-80.945176|80.945291222334149|121|1
35.323246|a07a34684ce7b42dd4af4d466633d06f9ad6fa29|1.39|2014-10-28 12:56:00|80.945290274299126|3|8265750067|166|35.414868531832361|0|44|31|-80.995484|4|35.444064|NON CARBONATED WATER|0.39|1|DEER PARK WATER 1LT|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00082657500676|BOTTLED WATER|G1 GROCERY|-80.945176|80.945291222334149|121|1
35.323246|efcd366903514c934d63e32d08a0ff3f59a8fa72|1.39|2014-10-14 11:05:00|80.945290274299126|3|8265750067|166|35.414868531832361|0|44|31|-80.995484|4|35.444064|NON CARBONATED WATER|0.39|1|DEER PARK WATER 1LT|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00082657500676|BOTTLED WATER|G1 GROCERY|-80.945176|80.945291222334149|121|1
35.323246|5f964c9b77a1f20402258dba6021d8cef9219887|1.39|2014-12-23 13:27:00|80.945290274299126|3|8265750067|166|35.414868531832361|0|44|31|-80.995484|4|35.444064|NON CARBONATED WATER|0.39|1|DEER PARK WATER 1LT|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00082657500676|BOTTLED WATER|G1 GROCERY|-80.945176|80.945291222334149|121|1
35.323246|880025674fb64a89767dc70bbbfe04e0b1286758|1.39|2014-10-08 11:09:00|80.945290274299126|3|8265750067|166|35.414868531832361|0|44|31|-80.995484|4|35.444064|NON CARBONATED WATER|0.39|1|DEER PARK WATER 1LT|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00082657500676|BOTTLED WATER|G1 GROCERY|-80.945176|80.945291222334149|121|1
35.323246|610845fe45ed2608bee8b5166364c08a203e58e4|1.39|2014-11-25 12:36:00|80.945290274299126|3|8265750067|166|35.414868531832361|0|44|31|-80.995484|4|35.444064|NON CARBONATED WATER|0.39|1|DEER PARK WATER 1LT|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00082657500676|BOTTLED WATER|G1 GROCERY|-80.945176|80.945291222334149|121|1
35.323246|1d3ffa7698727139fb0795ca4c8159546adcfd57|1.39|2014-11-19 14:38:00|80.945290274299126|3|8265750067|166|35.414868531832361|0|44|31|-80.995484|4|35.444064|NON CARBONATED WATER|0.39|1|DEER PARK WATER 1LT|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00082657500676|BOTTLED WATER|G1 GROCERY|-80.945176|80.945291222334149|121|1
35.323246|3efcc48574fafe9a7b574f66af20ee7bde51b8ef|1.39|2014-11-05 13:27:00|80.945290274299126|3|8265750067|166|35.414868531832361|0|44|31|-80.995484|4|35.444064|NON CARBONATED WATER|0.39|1|DEER PARK WATER 1LT|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00082657500676|BOTTLED WATER|G1 GROCERY|-80.945176|80.945291222334149|121|1
35.323246|feafbb2d6f9b03c8a41d46d54ff33f4df54432a3|1.39|2014-10-31 13:36:00|80.945290274299126|3|8265750067|166|35.414868531832361|0|44|31|-80.995484|4|35.444064|NON CARBONATED WATER|0.39|1|DEER PARK WATER 1LT|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00082657500676|BOTTLED WATER|G1 GROCERY|-80.945176|80.945291222334149|121|1
35.323246|498282b12dcc83318834ddcfc45752641030c525|1.39|2014-10-07 11:00:00|80.945290274299126|3|8265750067|166|35.414868531832361|0|44|31|-80.995484|4|35.444064|NON CARBONATED WATER|0.39|1|DEER PARK WATER 1LT|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00082657500676|BOTTLED WATER|G1 GROCERY|-80.945176|80.945291222334149|121|1
35.323246|677ac3ff6cd904b10d3ba321a535f1aff2d8898f|5.35|2014-09-20 11:04:00|1.4102725052409182|3|20165500000|166|0.6165069451919168|0|1|297|-80.945176|49|35.323246|GROUND BEEF|0.41|2|HT PREMIUM GRND BEEF 80% LEAN|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|0.61833652052202714|00201655000005|BEEF|MEAT|-80.945176|1.4127598348062935|166|1
35.323246|c79e3a3e6c37431f3f4eb13591148293b6152053|11.98|2014-11-18 19:51:00|80.945290274299126|3|1114110029|166|35.414868531832361|0|44|36|-80.995484|10|35.444064|PREMIUM GROUND|2.99|1|EIGHT OCLOCK ORIG GOUND COFFEE|8edfb943511219a6612ce4e5b12b643e5c5dc1ca|6.330899017926867|35.414868532563162|00011141100290|COFFEE|G1 GROCERY|-80.945176|80.945291222334149|121|2
35.103409|9061245f46c18e73ecd4c0fb4bc8420189eacd78|1.69|2014-10-28 06:36:00|1.4132775322775095|4|5200033875|88|0.6126700657242101|0|58|171|-80.992182|20|35.103409|ISOTONIC DRINKS|0.69|1|GATORADE COOL BLUE|90ec89769e7258d49986cbad016276d0b884794c|4.584592257176402|0.61177642288969325|00052000325553|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|ec37be68de8c007fc4a45c9cfef7bd157ac8637f|3.58|2014-09-23 06:40:00|1.4132775322775095|4|4850001775|88|0.6126700657242101|0|58|335|-80.992182|56|35.103409|ORANGE JUICE-REGRIGERATED|0.79|3|TROPICANA PP CALCIUM 12 OZ|90ec89769e7258d49986cbad016276d0b884794c|4.584592257176402|0.61177642288969325|00048500017760|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.992182|1.413580244274486|88|2
35.103409|c1e49bce4c9f35e01e9253e491382ebc5ace0de4|1.45|2014-09-23 06:40:00|1.4132775322775095|4|7203663220|88|0.6126700657242101|0|58|330|-80.992182|55|35.103409|EGGS|0.0|3|HT GRADE A    LARGE EGGS|90ec89769e7258d49986cbad016276d0b884794c|4.584592257176402|0.61177642288969325|00072036632203|EGGS FRESH|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|5c67f116a40f357d30e0f934b6027600b8371e3e|1.45|2014-10-03 06:34:00|1.4132775322775095|4|7203663220|88|0.6126700657242101|0|58|330|-80.992182|55|35.103409|EGGS|0.0|3|HT GRADE A    LARGE EGGS|90ec89769e7258d49986cbad016276d0b884794c|4.584592257176402|0.61177642288969325|00072036632203|EGGS FRESH|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|358c12792d72e9950751f46cbbfce8cbb0366842|4.97|2014-09-25 06:56:00|1.4132775322775095|4|7203658034|88|0.6126700657242101|0|58|358|-80.992182|100|35.103409|REGULAR BACON|1.47|19|HT THICK SLICED BACON|90ec89769e7258d49986cbad016276d0b884794c|4.584592257176402|0.61177642288969325|00072036580320|BACON|CASE READY MEATS|-80.992182|1.413580244274486|88|1
35.103409|abfaae4863968aa2134fb822ba46de6eee0858ed|0.97|2015-02-10 10:04:00|1.4132775322775095|4|7203698758|88|0.6126700657242101|0|58|31|-80.992182|4|35.103409|NON CARBONATED WATER|0.0|1|HT SPRING WATER|90ec89769e7258d49986cbad016276d0b884794c|4.584592257176402|0.61177642288969325|00072036987587|BOTTLED WATER|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|1f1d691b8e0ab414be880f6f299fffe753137b12|0.97|2015-01-28 07:35:00|1.4132775322775095|4|7203671102|88|0.6126700657242101|0|58|1025|-80.992182|162|35.103409|WHITE|0.0|7|HT OLD FASHIONED BREAD|90ec89769e7258d49986cbad016276d0b884794c|4.584592257176402|0.61177642288969325|00072036711021|SLICED BREAD|COMMERCIAL BAKERY|-80.992182|1.413580244274486|88|1
35.43259|ff3e86dad84592e620849f1de8a919a8e71224b7|5.99|2015-02-14 20:10:00|1.4057311447477159|4|3120020300|202|0.6184153580092175|0|52|130|-80.605588|20|35.43259|CRANBERRY JUICE/DRINKS-SHELF|0.0|1|OS CRANBERRY JUICE|93373d6d51d0723a2664eddb34347d298278bb0d|3.6576497896018707|0.6209993146566879|00031200203007|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.605588|1.406832906106031|202|1
35.43259|f03879a0df37bf4aca590fd8fa5b109a77fd843d|0.99|2014-12-24 17:21:00|1.4057311447477159|4|7203695306|202|0.6184153580092175|0|52|1895|-80.605588|450|35.43259|TEA|0.0|6|FFM HALF TEA/LEMONADE|93373d6d51d0723a2664eddb34347d298278bb0d|3.6576497896018707|0.6209993146566879|00072036018878|BEVERAGES|DELI|-80.605588|1.406832906106031|202|1
35.43259|ee06a67937dade55a17675a090330e5396a952a7|2.59|2015-01-10 17:37:00|80.607132136635443|4|7173000720|202|35.485524547245802|0|9|150|-80.662946|23|35.412407|NOODLES/DUMPLINGS-DRY|0.0|1|NO YOLKS DUMPLINGS|93373d6d51d0723a2664eddb34347d298278bb0d|3.6576497896018707|35.47365851958088|00071730007201|PASTA|G1 GROCERY|-80.605588|80.605618668188214|68|1
35.43259|55e9f9356ce33093ca81903254c74070da819a26|8.99|2014-12-24 17:24:00|1.4057311447477159|4|1200050404|202|0.6184153580092175|0|52|31|-80.605588|4|35.43259|NON CARBONATED WATER|2.2|1|AQUAFINA WATER 16.9 OZ 24 PK|93373d6d51d0723a2664eddb34347d298278bb0d|3.6576497896018707|0.6209993146566879|00012000504044|BOTTLED WATER|G1 GROCERY|-80.605588|1.406832906106031|202|1
35.43259|e7a200dda7c725c977dd8b25c9e5dbf4506ff535|1.52|2014-09-14 15:17:00|1.4057311447477159|4||202|0.6184153580092175|0|52|558|-80.605588|64|35.43259|SPECIALTY-VEGETABLES|0.0|4|COO GINGER ROOT, BULK|93373d6d51d0723a2664eddb34347d298278bb0d|3.6576497896018707|0.6209993146566879|00204612000001|FRESH PRODUCE|PRODUCE|-80.605588|1.406832906106031|202|1
35.17739|645ab251a9215994663cfd800a3383dc51807233|3.79|2014-11-15 15:05:00|80.801203185414451|1|980000633|208|35.198878721432052|0|24|45|-80.806073|7|35.106477|PEG GUM|0.0|1|TIC TAC FRUIT BOTTLE|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00009800006304|CANDY|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|350c1feb0242ea2238e3baecfa92a5c71cef601a|6.49|2015-02-07 18:26:00|80.801203185414451|1|89604000100|208|35.198878721432052|0|24|1866|-80.806073|435|35.106477|PIMENTO|0.0|6|PALMETTO JALAPENO PIMENTO CHSE|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00896040001011|SALADS|DELI|-80.80146|80.801479956400485|4|1
35.17739|b0bd16d07d9b733df2faa47c04ec0f490a79b450|2.99|2014-10-19 17:27:00|80.801203185414451|1|1410009840|208|35.198878721432052|0|24|1256|-80.806073|13|35.106477|WHOLESOME CRACKERS|0.99|1|PF BAKED NATURALS ITALIAN HERB|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00014100092292|CRACKERS|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|508ce955dcf3d5db074a819cb0d75753fcc076bd|6.49|2015-02-16 15:07:00|80.801203185414451|1|89604000100|208|35.198878721432052|0|24|1866|-80.806073|435|35.106477|PIMENTO|0.0|6|PALMETTO JALAPENO PIMENTO CHSE|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00896040001011|SALADS|DELI|-80.80146|80.801479956400485|4|1
35.17739|2eb2f0858412f72853ec3757ed676ab2cbb9ad3e|2.69|2015-02-23 15:39:00|80.801203185414451|1|1600026460|208|35.198878721432052|0|24|42|-80.806073|6|35.106477|GRANOLA/YOGURT BARS|0.0|1|NV BAR SWT SLTY PNUT|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00016000277076|BREAKFAST FOODS|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|8eea8fb1ecb471ab2a3bfd8a738300398d7a22bd|2.59|2014-09-23 17:14:00|80.801203185414451|1|79271600032|208|35.198878721432052|0|24|398|-80.806073|69|35.106477|NFS-BATHROOM CLEANERS|0.0|1|CLEAN SHOWER DAILY SHOWER CLEA|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00792716000329|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|3b5b0c85f1e4664c135431d611eb19efa5f2ef1a|1.19|2014-12-16 17:29:00|80.801203185414451|1|7488007017|208|35.198878721432052|0|24|80|-80.806073|34|35.106477|SEASONING PACKETS|0.0|1|SUNBIRD STIR FRY MIX|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00074880070040|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|d66d4ef689784da5fcdb140c956607b900d391be|2.69|2014-12-11 17:27:00|80.801203185414451|1|7512800016|208|35.198878721432052|0|24|1273|-80.806073|50|35.106477|BAG VEG NON STEAM|0.7|5|SAVANNAH SWT CORN HUSHPUPPY|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00075128000126|VEGETABLES-FROZEN|FROZEN|-80.80146|80.801479956400485|4|1
35.17739|6bcec92809a11a4952d3cfcb05bbdb8f0ea8c4d8|2.65|2015-02-09 12:18:00|80.801203185414451|1|8768400095|208|35.198878721432052|0|24|121|-80.806073|20|35.106477|ASEPTIC JUICES|0.15|1|CAPRI SUN FRUIT PUNCH 10 PK|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00087684001073|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|c42e4439202128d3639e3d5078ef43bbf9c1f051|8.27|2014-09-25 17:54:00|80.801203185414451|1|20249700000|208|35.198878721432052|0|24|297|-80.806073|49|35.106477|GROUND BEEF|0.42|2|NY STRIP STEAKBURGER 80% LEAN|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00202497000000|BEEF|MEAT|-80.80146|80.801479956400485|4|1
35.17739|04c758968ddbc63ceea7233080288fdecb694f97|2.77|2015-01-06 09:31:00|80.801203185414451|1|3338353030|208|35.198878721432052|0|24|523|-80.806073|64|35.106477|FRESH POTATOES|0.0|4|RUSSET POTATO 8LB BAG|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00033383530307|FRESH PRODUCE|PRODUCE|-80.80146|80.801479956400485|4|1
35.17739|f64f06512e2c3a522e3f6fbe730786a48c4aacae|4.29|2014-10-22 16:10:00|80.801203185414451|1|2840016014|208|35.198878721432052|0|24|201|-80.806073|31|35.106477|POTATO CHIPS|2.15|1|LAYS WAVY REGULAR|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00028400160209|SNACKS|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|374a6fca733b63433e7400729befb400861f0729|8.58|2014-12-13 17:54:00|80.801203185414451|1|2800028254|208|35.198878721432052|0|24|1134|-80.806073|57|35.106477|CARTON MILK|0.0|3|NESQUICK CHOCOLATE MILK|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00028000282547|MILK|DAIRY|-80.80146|80.801479956400485|4|2
35.17739|12ec76a90b353962ca6689b44ab174378acac85a|5.99|2014-10-14 17:12:00|80.801203185414451|1|1834175105|208|35.198878721432052|0|24|9934|-80.806073|885|35.106477|NFS POP CHARDONNAY|0.0|13|CB-BAREFOOT CHARDONNAY|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00018341751055|POPULAR (4-$7.99)|WINE|-80.80146|80.801479956400485|4|1
35.17739|f7ecaf1db853533aad78f70011e2161c9e4ff8d7|4.29|2014-12-08 16:41:00|80.801203185414451|1|2840016014|208|35.198878721432052|0|24|201|-80.806073|31|35.106477|POTATO CHIPS|0.29|1|LAYS WAVY REGULAR|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00028400160209|SNACKS|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|8da4e63829699ef25f4f0bb4a8e83c4fb6ecfafb|10.0|2014-10-07 22:27:00|80.801203185414451|1|1834175105|208|35.198878721432052|0|24|9934|-80.806073|885|35.106477|NFS POP CHARDONNAY|0.0|13|CB-BAREFOOT CHARDONNAY|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00018341751055|POPULAR (4-$7.99)|WINE|-80.80146|80.801479956400485|4|2
35.17739|04dbbec5af1ee7cff67b1bb72a0fbfe056bbd0ce|6.02|2015-01-29 15:30:00|80.801203185414451|1|20165700000|208|35.198878721432052|0|24|297|-80.806073|49|35.106477|GROUND BEEF|1.34|2|HT GROUND BEEF CHUCK 80% LEAN|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00201657000003|BEEF|MEAT|-80.80146|80.801479956400485|4|1
35.17739|acd76827ce2964f66508ee0f1c1fa0570bb522c0|6.11|2014-10-06 17:08:00|80.801203185414451|1|20165700000|208|35.198878721432052|0|24|297|-80.806073|49|35.106477|GROUND BEEF|0.68|2|HT GROUND BEEF CHUCK 80% LEAN|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00201657000003|BEEF|MEAT|-80.80146|80.801479956400485|4|1
35.17739|29760fc7443b6c9585c5a9087ce562b937cb29ff|4.08|2014-12-10 16:45:00|80.801203185414451|1|20165700000|208|35.198878721432052|0|24|297|-80.806073|49|35.106477|GROUND BEEF|0.45|2|HT GROUND BEEF CHUCK 80% LEAN|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00201657000003|BEEF|MEAT|-80.80146|80.801479956400485|4|1
35.17739|ba8a727ab604857ef04b51f5e85bbc549bfadeac|5.12|2015-02-08 17:55:00|80.801203185414451|1|20165700000|208|35.198878721432052|0|24|297|-80.806073|49|35.106477|GROUND BEEF|0.91|2|HT GROUND BEEF CHUCK 80% LEAN|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00201657000003|BEEF|MEAT|-80.80146|80.801479956400485|4|1
35.17739|8882fc64f2e94270f6590ab594d3cc2e3a3a5da3|6.87|2014-12-09 16:48:00|80.801203185414451|1|20165700000|208|35.198878721432052|0|24|297|-80.806073|49|35.106477|GROUND BEEF|0.77|2|HT GROUND BEEF CHUCK 80% LEAN|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00201657000003|BEEF|MEAT|-80.80146|80.801479956400485|4|1
35.17739|2c3517ab2c0eae1283e7a4efaf31245325b33a5e|3.99|2014-09-11 18:11:00|80.801203185414451|1|7464100992|208|35.198878721432052|0|24|562|-80.806073|64|35.106477|FRESH CUT FRUIT|0.0|4|RED APPLE SLICES 14OZ|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00074641009920|FRESH PRODUCE|PRODUCE|-80.80146|80.801479956400485|4|1
35.17739|5869d0c4632939c4c7f525312914a1bd86d83938|1.67|2015-01-30 18:03:00|80.801203185414451|1|2800008040|208|35.198878721432052|0|24|53|-80.806073|7|35.106477|THEATER BOX|0.0|1|WONKA RUNTS THEATER BOX|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00079200472146|CANDY|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|4c08464f9c33de85087b56c60667738b42a4c100|19.12|2014-12-21 17:11:00|80.801203185414451|1|20128300000|208|35.198878721432052|0|24|296|-80.806073|49|35.106477|RANCHER BEEF|0.0|2|VALUE PK BEEF RIBEYE STK BNLS|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00201283000002|BEEF|MEAT|-80.80146|80.801479956400485|4|1
35.17739|d583c0da8c16b54228bb641312c57e3392ad919b|4.99|2014-11-22 18:02:00|80.801203185414451|1|4950800821|208|35.198878721432052|0|24|1980|-80.806073|480|35.106477|CHOCOLATES|1.0|6|WHITE CHOC PRETZEL CRISPS|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00049508008217|DRY GOODS|DELI|-80.80146|80.801479956400485|4|1
35.17739|b37ec918efd7109b071f7757b266ce8b4b92254a|6.79|2014-12-28 18:50:00|80.801203185414451|1|7064003404|208|35.198878721432052|0|24|252|-80.806073|45|35.106477|PREMIUM ICE CREAM|2.81|5|B BUNNY PREM BIRTHDAY PARTY|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00070640003112|ICE CREAM|FROZEN|-80.80146|80.801479956400485|4|1
35.17739|1f29079fea9073f28b64cc6b9df70e914d469439|4.49|2015-01-11 17:54:00|80.801203185414451|1|5200012125|208|35.198878721432052|0|24|171|-80.806073|20|35.106477|ISOTONIC DRINKS|0.61|1|GATORADE ASTAR RAIN BERRY 6PK|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00052000122152|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|883babbec4cdc094326a0a7a3b7de3ea23044a48|4.49|2015-01-07 17:11:00|80.801203185414451|1|5200012125|208|35.198878721432052|0|24|171|-80.806073|20|35.106477|ISOTONIC DRINKS|0.61|1|GATORADE ASTAR RAIN BERRY 6PK|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00052000122152|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|b6427b1ab853778581a61b5b8df71228d5aa382b|1.99|2014-09-17 11:19:00|80.801203185414451|1|5210000738|208|35.198878721432052|0|24|1245|-80.806073|34|35.106477|SINGLE SPICES|0.0|1|MC PARSLEY FLAKES|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00052100007380|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|d54ded96a3216513040aed00a0ed432e1123a44d|4.49|2015-01-19 17:50:00|80.801203185414451|1|5200012125|208|35.198878721432052|0|24|171|-80.806073|20|35.106477|ISOTONIC DRINKS|0.71|1|GATORADE ASTAR RAIN BERRY 6PK|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00052000122152|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|0af024273552d6bdfa310e9be3638340b80ccc39|4.49|2015-01-05 15:48:00|80.801203185414451|1|5200012125|208|35.198878721432052|0|24|171|-80.806073|20|35.106477|ISOTONIC DRINKS|0.61|1|GATORADE ASTAR RAIN BERRY 6PK|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00052000122152|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|f244ad1b308a4fa70490302cce6829fe8909f0f6|3.49|2014-12-31 18:44:00|80.801203185414451|1|88491212971|208|35.198878721432052|0|24|81|-80.806073|9|35.106477|RTE CEREAL KIDS|0.0|1|POST PEBBLES FRUITY|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00884912129710|CEREAL|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|fcea3ed25aa80cc86da63d23dbc753f3a5fe218d|3.38|2014-10-11 17:12:00|80.801203185414451|1|7203698517|208|35.198878721432052|0|24|426|-80.806073|72|35.106477|NFS-PAPER TOWELS|0.0|1|YH ULT TOWEL 1 ROLL WHITE|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00072036010711|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.80146|80.801479956400485|4|2
35.17739|dd6937c5c62af37dab31f0ef87d820f1903b16e9|1.69|2014-10-07 18:15:00|80.801203185414451|1|7203698517|208|35.198878721432052|0|24|426|-80.806073|72|35.106477|NFS-PAPER TOWELS|0.0|1|YH ULT TOWEL 1 ROLL WHITE|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00072036010711|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|36a8cac03aceddbba76f27283f4238caf45d8b59|3.5|2014-11-17 10:43:00|80.801203185414451|1|7203603041|208|35.198878721432052|0|24|220|-80.806073|34|35.106477|PEPPER|1.0|1|E  HT BLACK PEPPER|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00072036030412|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|8d0f39308a63085dc470b17491e339435a04ba43|3.38|2015-03-04 21:00:00|80.801203185414451|1|7203698517|208|35.198878721432052|0|24|426|-80.806073|72|35.106477|NFS-PAPER TOWELS|0.71|1|YH ULT TOWEL 1 ROLL WHITE|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00072036010711|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.80146|80.801479956400485|4|2
35.17739|5b2a52b8d0f629fbac6ce209b3c1e8dd2626febe|1.17|2014-09-18 14:09:00|80.801203185414451|1|7203628044|208|35.198878721432052|0|24|161|-80.806073|25|35.106477|PEPPERS|0.0|1|HT JALAPENO SLICES|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00072036280442|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|799a42ee43a2407959d868c4471272b51fdf08fd|2.59|2014-09-21 19:20:00|80.801203185414451|1|7203615048|208|35.198878721432052|0|24|1469|-80.806073|278|35.106477|REGULAR CUT FRIES|0.3|5|HT STEAK FRIES|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00072036490223|FROZEN POTATO|FROZEN|-80.80146|80.801479956400485|4|1
35.17739|21070052efd8b6788e39d2bf6d20488bd9f056bb|2.59|2015-02-11 17:32:00|80.801203185414451|1|7203615048|208|35.198878721432052|0|24|1469|-80.806073|278|35.106477|REGULAR CUT FRIES|0.0|5|HT STEAK FRIES|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00072036490223|FROZEN POTATO|FROZEN|-80.80146|80.801479956400485|4|1
35.17739|76f10be7720c0e5eaafbc3763689e1c42b67719e|1.29|2014-11-09 13:34:00|80.801203185414451|1|2200000667|208|35.198878721432052|0|24|48|-80.806073|7|35.106477|REGISTER GUM|0.0|1|WRIGLEY'S JUICY FRUIT 15 PC|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00022000006677|CANDY|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|be8a18210657afab543202b4c6cca850079a06d2|5.98|2015-02-12 19:19:00|80.801203185414451|1|1200081331|208|35.198878721432052|0|24|854|-80.806073|32|35.106477|LIQUID ICED COFFEES|0.2|1|FRAPPUCCINO VANILLA SINGLE|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00012000813313|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.80146|80.801479956400485|4|2
35.17739|501e95fdce77dbd0928adae76456f8ee182fe91e|4.65|2014-12-14 17:05:00|80.801203185414451|1|78616201000|208|35.198878721432052|0|24|31|-80.806073|4|35.106477|NON CARBONATED WATER|1.6500000000000001|1|VIT WATER XXX 20 OZ|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00786162150004|BOTTLED WATER|G1 GROCERY|-80.80146|80.801479956400485|4|3
35.17739|66c655e87e827d490624cd9aa6d4171f05d2f6bb|5.29|2014-11-19 17:24:00|80.801203185414451|1|7104000015|208|35.198878721432052|0|24|332|-80.806073|52|35.106477|STRING/SNACK|0.0|3|POLLY-O-TWISTARELLAS|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00071040065311|CHEESE|DAIRY|-80.80146|80.801479956400485|4|1
35.17739|d166f19a496d7ac4b038239b28e5f9e26d38a49b|4.69|2014-09-10 14:01:00|80.801203185414451|1|6927603205|208|35.198878721432052|0|24|79|-80.806073|273|35.106477|ASIAN SAUCES/SEASONINGS|0.0|1|PATAK PASTE CURRY MILD|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00069276032054|ASIAN PREP. FOODS|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|7dabb3cb8bc578eec498f30c4fba96754d95b759|1.25|2014-10-01 14:53:00|80.801203185414451|1|4900005537|208|35.198878721432052|0|24|54|-80.806073|8|35.106477|DIET|0.26|23|DIET COKE 1.25 LITER BOTTLE|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00049000055399|CARBONATED BEVERAGES|BEVERAGE|-80.80146|80.801479956400485|4|1
35.17739|bb1845164eb69effedeaed47a90e81cae7262203|3.38|2014-12-13 12:34:00|80.801203185414451|1|4900000044|208|35.198878721792063|0|24|55|-80.824767|8|35.116751|REGULAR|0.0|23|CB COKE SINGLE 20 OZ.|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00049000000443|CARBONATED BEVERAGES|BEVERAGE|-80.80146|80.80147936731997|294|2
35.17739|8b4bf6fb8ac4df66851575cb49f4feba5ef3b4f6|2.69|2014-11-13 14:47:00|80.801203185414451|1|5210015742|208|35.198878721432052|0|24|80|-80.806073|34|35.106477|SEASONING PACKETS|0.0|1|MC CHICK BAG N SEASON|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00052100157467|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|ad7bfdac1f5a1b094479404483aafc41e42be650|1.49|2015-02-28 15:39:00|80.801203185414451|1|4900005537|208|35.198878721432052|0|24|54|-80.806073|8|35.106477|DIET|0.49|23|DIET COKE 1.25 LITER BOTTLE|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00049000055399|CARBONATED BEVERAGES|BEVERAGE|-80.80146|80.801479956400485|4|1
35.17739|fadd202a1ffcb1a7baf2a863b02afe68be1a4f6c|1.69|2014-11-07 07:31:00|80.801203185414451|1|4900000044|208|35.198878721432052|0|24|55|-80.806073|8|35.106477|REGULAR|0.0|23|CB COKE SINGLE 20 OZ.|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00049000000443|CARBONATED BEVERAGES|BEVERAGE|-80.80146|80.801479956400485|4|1
35.17739|da0c8af259feec64502944915a8687027867e935|1.69|2014-12-24 11:11:00|80.801203185414451|1|4900000044|208|35.198878721432052|0|24|55|-80.806073|8|35.106477|REGULAR|0.0|23|CB COKE SINGLE 20 OZ.|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00049000000443|CARBONATED BEVERAGES|BEVERAGE|-80.80146|80.801479956400485|4|1
35.17739|4a34d5e1e411dd87382117f2e0916e1501533241|13.99|2014-10-03 17:03:00|80.801203185414451|1|7203695572|208|35.198878721432052|0|24|1653|-80.806073|381|35.106477|CELEBRATION CAKES|0.0|14|1/8 SHEET DL WHITE WHIP TOPPIN|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00072036955722|CAKES|BAKERY|-80.80146|80.801479956400485|4|1
35.17739|9c03692c10a50fc08bd98e028a63f0ee43277b1e|0.97|2014-12-17 17:15:00|80.801203185414451|1|7203637031|208|35.198878721432052|0|24|212|-80.806073|33|35.106477|CONDENSED SOUP|0.17|1|HT SP RS CRM MUSHROOM|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00072036978547|SOUP|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|2dcc8ae709263f366bbe76e6b27a5dc65e687c97|0.97|2014-12-17 17:11:00|80.801203185414451|1|7203637031|208|35.198878721432052|0|24|212|-80.806073|33|35.106477|CONDENSED SOUP|0.17|1|HT SP RS CRM MUSHROOM|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00072036978547|SOUP|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|ab9e5bd5739a8ab095c2169ee352592ceacc1f67|3.88|2014-11-14 11:18:00|80.801203185414451|1|7203637031|208|35.198878721432052|0|24|212|-80.806073|33|35.106477|CONDENSED SOUP|0.0|1|HT SP RS CRM MUSHROOM|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00072036978547|SOUP|G1 GROCERY|-80.80146|80.801479956400485|4|4
35.17739|87510c7f2ac823d5f3e7480f8ffe391224030912|1.69|2015-01-10 16:32:00|80.801203185414451|1|7203688003|208|35.198878721432052|0|24|527|-80.806073|64|35.106477|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00072036880031|FRESH PRODUCE|PRODUCE|-80.80146|80.801479956400485|4|1
35.17739|abe33be81179d75d2c6fa4b014c2494d627da129|1.19|2015-01-27 16:09:00|80.801203185414451|1|7203653022|208|35.198878721432052|0|24|1273|-80.806073|50|35.106477|BAG VEG NON STEAM|0.0|5|HT BABY BUD BROCCOLI FLORETS|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00072036530790|VEGETABLES-FROZEN|FROZEN|-80.80146|80.801479956400485|4|1
35.17739|f7c3e69f02fe709f877c9839f42804db04339329|1.19|2015-01-15 15:10:00|80.801203185414451|1|7203653022|208|35.198878721432052|0|24|1273|-80.806073|50|35.106477|BAG VEG NON STEAM|0.0|5|HT BABY BUD BROCCOLI FLORETS|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00072036530790|VEGETABLES-FROZEN|FROZEN|-80.80146|80.801479956400485|4|1
35.17739|9f758598de5f73a2cfdc7b3fd5193da99e32b0d9|0.73|2014-11-10 12:06:00|80.801203185414451|1||208|35.198878721432052|0|24|524|-80.806073|64|35.106477|FRESH PROD FRESH ONIONS|0.0|4|COO YELLOW ONIONS, LRG|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00204665000003|FRESH PRODUCE|PRODUCE|-80.80146|80.801479956400485|4|1
35.17739|decaa7626b05ab030f28d02c030176036ef976d6|0.47|2014-12-19 17:52:00|80.801203185414451|1||208|35.198878721432052|0|24|524|-80.806073|64|35.106477|FRESH PROD FRESH ONIONS|0.0|4|COO YELLOW ONIONS, LRG|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00204665000003|FRESH PRODUCE|PRODUCE|-80.80146|80.801479956400485|4|1
35.17739|e72128f595709e965ec100edf507b839264be81a|2.99|2015-01-25 18:34:00|80.801203185414451|1|7433610102|208|35.198878721432052|0|24|342|-80.806073|57|35.106477|FRESH MILK|0.0|3|HIGHLAND CREST WHOLE MILK|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00074336879203|MILK|DAIRY|-80.80146|80.801479956400485|4|1
35.17739|c2d0dae31df35b6ebf115a5e7a193be9fa3d5703|11.98|2014-09-23 10:53:00|80.801203185414451|1|7403008182|208|35.198878721432052|0|24|2017|-80.806073|505|35.106477|STRETCHED CURD CHEESE|3.0|6|SORRENTO FRESH MOZZARELLA|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00074030081827|SPECIALTY CHEESE|DELI|-80.80146|80.801479956400485|4|2
35.17739|88284cbbf361842eaca5ce1a4812787bfbc2ab3b|3.59|2014-10-09 17:49:00|80.801203185414451|1|7433610102|208|35.198878721432052|0|24|342|-80.806073|57|35.106477|FRESH MILK|0.0|3|HIGHLAND CREST WHOLE MILK|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00074336879203|MILK|DAIRY|-80.80146|80.801479956400485|4|1
35.17739|0cbaa3bf91ba6172a30f0bafd2beaf5305150ea8|2.29|2014-12-15 16:57:00|80.801203185414451|1|7800023046|208|35.198878721432052|0|24|55|-80.806073|8|35.106477|REGULAR|1.29|23|CHERRY 7 UP 2LTR NR|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00078000005318|CARBONATED BEVERAGES|BEVERAGE|-80.80146|80.801479956400485|4|1
35.17739|a70a3801ff25468f56d558ce350c9643eabec0f9|2.29|2014-12-19 07:30:00|80.801203185414451|1|7800023046|208|35.198878721432052|0|24|55|-80.806073|8|35.106477|REGULAR|1.29|23|CHERRY 7 UP 2LTR NR|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00078000005318|CARBONATED BEVERAGES|BEVERAGE|-80.80146|80.801479956400485|4|1
35.17739|ac5199808197745252ff888cd1ce3c2b0242c258|6.89|2015-01-17 18:48:00|80.801203185414451|1|7790031101|208|35.198878721432052|0|24|1271|-80.806073|41|35.106477|PROTEIN BREAKFAST|0.0|5|J DEAN SAUSAGE BISCUIT 10CT|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00077900311017|BREAKFAST FOODS FROZEN|FROZEN|-80.80146|80.801479956400485|4|1
35.17739|df02ff9d27c69795c39fa3ac7d98620a5a9cb173|2.79|2014-10-24 15:27:00|80.801203185414451|1|7203698374|208|35.198878721432052|0|24|423|-80.806073|72|35.106477|NFS-DISPOSE PLATES/BOWLS|0.79|1|YH ULTRA DESIGNER PLATES|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00072036983756|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|1f19c0be98d1f9ac4d6b34621befeb94c37332d9|3.49|2014-09-27 13:21:00|80.801203185414451|1|65724334603|208|35.198878721432052|0|24|273|-80.806073|43|35.106477|PREMIUM NOVELTIES|0.0|5|PHILLY SWIRL POPPERZ|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00657243346039|FROZEN NOVELTIES|FROZEN|-80.80146|80.801479956400485|4|1
35.17739|4f1e1317e175482ba86a72b020c10624505cf734|1.5|2014-11-25 09:00:00|80.801203185414451|1|7203663107|208|35.198878721432052|0|24|1262|-80.806073|57|35.106477|HALF N HALF WHIPPING CREAM|0.0|3|HT HALF & HALF|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00072036632036|MILK|DAIRY|-80.80146|80.801479956400485|4|1
35.17739|94b9282127d456223196a5aced084c60ed2dc822|2.59|2014-11-07 19:18:00|80.801203185414451|1|7203663996|208|35.198878721432052|0|24|342|-80.806073|57|35.106477|FRESH MILK|0.0|3|HARRIS TEETER WHOLE MILK|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00072036639967|MILK|DAIRY|-80.80146|80.801479956400485|4|1
35.17739|246c01d4716a0b29f7abc9f58c4fede7ad369a35|3.99|2015-01-09 16:38:00|80.801203185414451|1|7127930108|208|35.198878721432052|0|24|555|-80.806073|64|35.106477|PACKAGED SALADS|0.0|4|F.E. BACON CAESAR KIT|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00071279301082|FRESH PRODUCE|PRODUCE|-80.80146|80.801479956400485|4|1
35.17739|7f8bd4451fb03e5b4da1d6633908c0e901a5ee57|3.79|2015-03-04 17:23:00|80.801203185414451|1|7169123097|208|35.198878721432052|0|24|5697|-80.806073|1520|35.106477|RM TAKE ALONG FOOD STORAGE|1.14|18|TAKEALONG TWIST&SEAL 1 CUP|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00071691394549|PLASTIC FOOD STORAGE|GM|-80.80146|80.801479956400485|4|1
35.17739|7158bb248783900b7ff736f3491e69ff9edd1361|4.99|2015-02-19 19:55:00|80.801203185414451|1|7124920730|208|35.198878721432052|0|24|3536|-80.806073|1045|35.106477|SHAMPOO-PREMIUM|1.0|17|S/C LOR ADV HC ULT STRGHT SHAM|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00071249292372|HAIR & SCALP CARE|HBC|-80.80146|80.801479956400485|4|1
35.17739|6bee77e3dcdf630644a68d7222d0b1afbe53e34e|3.99|2015-01-08 14:47:00|80.801203185414451|1|7127930108|208|35.198878721432052|0|24|555|-80.806073|64|35.106477|PACKAGED SALADS|0.0|4|F.E. BACON CAESAR KIT|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00071279301082|FRESH PRODUCE|PRODUCE|-80.80146|80.801479956400485|4|1
35.17739|1787459b6faea0ba8bad5635439396da326cc584|3.99|2014-09-19 17:04:00|80.801203185414451|1|7127930108|208|35.198878721432052|0|24|555|-80.806073|64|35.106477|PACKAGED SALADS|0.0|4|F.E. BACON CAESAR KIT|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00071279301082|FRESH PRODUCE|PRODUCE|-80.80146|80.801479956400485|4|1
35.17739|d5bb74e571064ebdf6c1476335865949e2a50ff3|2.57|2014-09-10 07:58:00|80.801203185414451|1|4410010167|208|35.198878721432052|0|24|341|-80.806073|57|35.106477|CREAMERS|0.0|3|COFFEE DREAM CRMR-FRENCH VAN|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00044100101670|MILK|DAIRY|-80.80146|80.801479956400485|4|1
35.17739|16daa57d6f5b9908f2d2bab0b2e115596eeba344|2.69|2015-03-01 22:54:00|80.801203185414451|1|4400001556|208|35.198878721432052|0|24|87|-80.806073|13|35.106477|CHEESE CRACKERS|0.35|1|CHEESE NIPS CHEDDAR|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00044000034535|CRACKERS|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|1a7a4ce16c764ca93391a3fd294f5af8e928f88d|1.97|2014-11-06 08:15:00|80.801203185414451|1|7203698240|208|35.198878721432052|0|24|442|-80.806073|76|35.106477|NFS-COOKING-STORAGE BAGS|0.0|1|YH RESEALABLE SANDWICH BAGS|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00072036982407|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|9debb0631aeec47a88e49445a7f7ca03d9465962|10.99|2014-12-18 15:02:00|80.801203185414451|1|8224228043|208|35.198878721432052|0|24|9960|-80.806073|887|35.106477|NFS-S/PREM-CAB SAUVIGNON|0.0|13|NOBLE VINES 337 CABERNET SAUV|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00082242280433|SUPER PREMIUM ($11-$14.99)|WINE|-80.80146|80.801479956400485|4|1
35.17739|7681376dec18b018c0b539b6238574756c1a32f3|2.85|2014-12-08 08:43:00|80.801203185414451|1|3040077852|208|35.198878721432052|0|24|427|-80.806073|72|35.106477|NFS-TOILET TISSUE|0.0|1|ANGEL SOFT SOFT/STRONG 4DR|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00030400778520|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|9f8d93afa34b1e1eb80cb24ed568b3ecd243487a|2.39|2015-02-08 12:48:00|80.801203185414451|1|7084781116|208|35.198878721432052|0|24|97|-80.806073|8|35.106477|ENERGY DRINKS|0.0|23|MONSTER ABSOLUTELY ZERO CAN|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00070847000037|CARBONATED BEVERAGES|BEVERAGE|-80.80146|80.801479956400485|4|1
35.17739|36015ba09c43bd838640796c0f9c02efbb844174|4.29|2014-11-08 13:09:00|80.801203185414451|1|2840006399|208|35.198878721432052|0|24|204|-80.806073|31|35.106477|TORTILLA CHIPS|1.79|1|TOSTITOS HINT OF LIME|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00028400064040|SNACKS|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|d773209ad51ae7561a639263851e91b36f4cd7fd|3.99|2014-12-29 16:50:00|80.801203185414451|1|2100067148|208|35.198878721432052|0|24|1441|-80.806073|274|35.106477|MAC AND CHEESE|0.0|1|KRAFT DIN EASY MAC EXTREME|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00021000778539|PREP FOODS DINNERS|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|21e9cd07ae89a0c90def2d24ec6e9d0612ac4092|2.19|2014-11-22 14:11:00|80.801203185414451|1|4900005010|208|35.198878721432052|0|24|55|-80.806073|8|35.106477|REGULAR|0.2|23|CLASSIC COKE 2 LT CONTOUR|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00049000050103|CARBONATED BEVERAGES|BEVERAGE|-80.80146|80.801479956400485|4|1
35.17739|8c77896dc4e71286cb080a72179f5bd79399e303|7.79|2014-12-15 21:00:00|80.801203185414451|1|5400036413|208|35.198878721432052|0|24|427|-80.806073|72|35.106477|NFS-TOILET TISSUE|1.8|1|SCOTT BATH SOFT 12 RL|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00054000364136|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|f0287dc804501d4bcd568d7434ee7d8d24bab880|2.19|2015-01-13 16:23:00|80.801203185414451|1|4900005010|208|35.198878721432052|0|24|55|-80.806073|8|35.106477|REGULAR|0.2|23|CLASSIC COKE 2 LT CONTOUR|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00049000050103|CARBONATED BEVERAGES|BEVERAGE|-80.80146|80.801479956400485|4|1
35.17739|777c1e77f191d303bee5ce0ab39c7710bf258593|2.19|2014-10-31 17:38:00|80.801203185414451|1|4900005010|208|35.198878721432052|0|24|55|-80.806073|8|35.106477|REGULAR|0.2|23|CLASSIC COKE 2 LT CONTOUR|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00049000050103|CARBONATED BEVERAGES|BEVERAGE|-80.80146|80.801479956400485|4|1
35.17739|21beaf7abb9a8862ad3b1c9ceb4c44ef5b71e541|2.19|2014-12-02 16:47:00|80.801203185414451|1|4900005010|208|35.198878721432052|0|24|55|-80.806073|8|35.106477|REGULAR|0.2|23|CLASSIC COKE 2 LT CONTOUR|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00049000050103|CARBONATED BEVERAGES|BEVERAGE|-80.80146|80.801479956400485|4|1
35.17739|9f80d1030f9c399f6692f3829c115cb70143862d|2.19|2014-12-24 15:33:00|80.801203185414451|1|4900005010|208|35.198878721432052|0|24|55|-80.806073|8|35.106477|REGULAR|0.0|23|CLASSIC COKE 2 LT CONTOUR|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00049000050103|CARBONATED BEVERAGES|BEVERAGE|-80.80146|80.801479956400485|4|1
35.17739|1b1b9acda595ff7aac40e7931af91081bbaf86c5|2.19|2015-02-02 15:55:00|80.801203185414451|1|4900005010|208|35.198878721432052|0|24|55|-80.806073|8|35.106477|REGULAR|0.2|23|CLASSIC COKE 2 LT CONTOUR|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00049000050103|CARBONATED BEVERAGES|BEVERAGE|-80.80146|80.801479956400485|4|1
35.17739|5e5dc2047f0627785d7fa130b2931f2fc44464d6|2.19|2014-12-01 07:37:00|80.801203185414451|1|4900005010|208|35.198878721432052|0|24|55|-80.806073|8|35.106477|REGULAR|0.2|23|CLASSIC COKE 2 LT CONTOUR|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00049000050103|CARBONATED BEVERAGES|BEVERAGE|-80.80146|80.801479956400485|4|1
35.17739|2bc45d07c59e1324f2debed6389ea542dd669ff2|2.19|2015-01-20 17:32:00|80.801203185414451|1|4900005010|208|35.198878721432052|0|24|55|-80.806073|8|35.106477|REGULAR|0.2|23|CLASSIC COKE 2 LT CONTOUR|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00049000050103|CARBONATED BEVERAGES|BEVERAGE|-80.80146|80.801479956400485|4|1
35.17739|21de6ba44b99fbec092ab03d1e9f0ef0d09e7f3f|9.98|2014-12-09 20:28:00|80.801203185414451|1|3980001132|208|35.198878721432052|0|24|8433|-80.806073|1769|35.106477|ALKALINE AA|4.0|18|(FE)ER BATTERY E91BP4 SZ AA|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00039800011329|BATTERY & FLASHLIGHT|GM|-80.80146|80.801479956400485|4|2
35.17739|94002e19ccfa1b6cd5c238184701963a90382c2f|1.79|2014-11-24 18:03:00|80.801203185414451|1|7203688032|208|35.198878721432052|0|24|555|-80.806073|64|35.106477|PACKAGED SALADS|0.0|4|HT SHREDDED ICEBERG LETTUCE|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00072036880321|FRESH PRODUCE|PRODUCE|-80.80146|80.801479956400485|4|1
35.17739|2d75dacf90a3eee91c3bf1c7b01836a01dc5365f|3.1|2014-09-24 08:47:00|80.801203185414451|1|3700000445|208|35.198878721432052|0|24|725|-80.806073|66|35.106477|NFS-DISHWASHING LIQUID|0.55|1|DAWN LIQ DISH ORIGINAL 9OZ|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00037000004455|DETERGENTS|G1 GROCERY|-80.80146|80.801479956400485|4|2
35.17739|464f96b95e3875e4605fef7bc1ebcc76d2e2df20|3.49|2014-10-12 17:55:00|80.801203185414451|1|2840024053|208|35.198878721432052|0|24|198|-80.806073|31|35.106477|CORN CHIPS|1.75|1|FRITOS SCOOPS|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00028400240628|SNACKS|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|c64181f64bb820b837c88e41b57882385b68cf7c|2.75|2014-11-19 10:29:00|80.801203185414451|1|1920002522|208|35.198878721432052|0|24|404|-80.806073|69|35.106477|NFS-TOILET BOWL CLEANERS|0.0|1|LYSOL TOILET BOWL CLEANER|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00019200025225|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|711b16f7ce2940b514cffd291530d2bcffa4c6af|1.99|2015-01-10 20:20:00|80.801203185414451|1|3400040568|208|35.198878721432052|0|24|46|-80.806073|7|35.106477|PKG CHOC|0.49|1|HERSHEY MILK 8 PACK|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00034000070152|CANDY|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|ea61fbd3fc3da16086d56aaa5a7a06eaf35cfedd|4.99|2014-11-24 21:14:00|80.801203185414451|1|3500076233|208|35.198878721432052|0|24|4092|-80.806073|1080|35.106477|TOOTHPASTE-WHITENING|1.49|17|COLG OPTIC WH CRYSTL MINT TPST|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00035000763761|ORAL HYGIENE|HBC|-80.80146|80.801479956400485|4|1
35.17739|ec860782a0aed0310d248393825043698214e01b|2.59|2015-02-13 20:34:00|80.801203185414451|1|7203615048|208|35.198878721432052|0|24|1469|-80.806073|278|35.106477|REGULAR CUT FRIES|0.0|5|HT CRINKLE CUT FRIES|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00072036490216|FROZEN POTATO|FROZEN|-80.80146|80.801479956400485|4|1
35.17739|68afd677d3537689961901ec62ff115347aaa78e|5.39|2014-10-22 10:48:00|80.801203185414451|1|2570071016|208|35.198878721432052|0|24|398|-80.806073|69|35.106477|NFS-BATHROOM CLEANERS|1.89|1|SCRUB BUBBLE SHOWER FOAM TRIG|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00025700710165|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|a27267576757807963a0e6cad032e1a44ad025e5|4.59|2014-12-23 21:03:00|80.801203185414451|1|2420006040|208|35.198878721432052|0|24|389|-80.806073|66|35.106477|NFS-LAUNDRY DETERGENTS|0.6|1|PUREX HE LIQUID DETERGENT|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00024200023508|DETERGENTS|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|4bfea2bb97a6b0cf726b5006e687df9f7293836e|4.59|2014-11-09 16:19:00|80.801203185414451|1|2420006040|208|35.198878721432052|0|24|389|-80.806073|66|35.106477|NFS-LAUNDRY DETERGENTS|1.25|1|PUREX HE LIQUID DETERGENT|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00024200023508|DETERGENTS|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|4481398270643aed46f556043f73cf0a56d67aaa|13.99|2014-10-24 19:59:00|80.801203185414451|1|1820005990|208|35.198878721432052|0|24|456|-80.806073|82|35.106477|DOMESTIC SUPER PREM 12PK&>|0.0|16|MICHELOB ULTRA 12PK 12OZ BTL|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00018200059902|DOMESTIC BEER|BEER|-80.80146|80.801479956400485|4|1
35.17739|8b8801d566a7cff08e8e9559abff41537a4603cb|2.49|2014-10-06 07:30:00|80.801203185414451|1|1410008550|208|35.198878721432052|0|24|87|-80.806073|13|35.106477|CHEESE CRACKERS|0.0|1|PP GF FLAVOR BLAST ORIGINAL|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00014100085485|CRACKERS|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|c6cd337a55e995b3cc3bff994457699e1d60e272|5.59|2015-01-12 11:10:00|80.801203185414451|1|20600100000|208|35.198878721432052|0|24|1802|-80.806073|400|35.106477|FFM HAM|0.0|6|VIRGINIA BAKED HAM|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00206001000005|FFM MEAT|DELI|-80.80146|80.801479956400485|4|1
35.17739|f6b728c545d17a632e90619d848ef5fc5ea65d01|1.79|2014-12-11 21:12:00|80.801203185414451|1|7339000393|208|35.198878721432052|0|24|48|-80.806073|7|35.106477|REGISTER GUM|0.0|1|MENTOS RED FRUIT GUM 15CT|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00073390003937|CANDY|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|5985356c6364cc604619c6e1213281b78c5e451a|5.39|2014-12-18 10:58:00|80.801203185414451|1|3450015193|208|35.198878721432052|0|24|312|-80.806073|51|35.106477|BUTTER|1.89|3|LOL BUTTER HALF STICKS|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00034500151818|BUTTER & MARGARINE|DAIRY|-80.80146|80.801479956400485|4|1
35.17739|e96dfd1b108f39f6e34797c7bbe87f631c6dfe44|7.78|2015-01-15 15:13:00|80.801203185414451|1|3700029213|208|35.198878721432052|0|24|393|-80.806073|68|35.106477|NFS-AIR FRESHENERS|1.78|1|FEBREZE SR GAIN ISLAND FRESH|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00037000905011|FRESHENERS/DEODORIZERS|G1 GROCERY|-80.80146|80.801479956400485|4|2
35.17739|55434be3d809d41348286084cbfb3506e0036e13|8.99|2015-02-28 20:34:00|80.801203185414451|1|8383700626|208|35.198878721432052|0|24|9952|-80.806073|886|35.106477|NFS-PREM-PINOT NOIR|0.0|13|CASTLE ROCK PINOT NOIR|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00083837006261|PREMIUM ($8-$10.99)|WINE|-80.80146|80.801479956400485|4|1
35.17739|6031472ba9edc3b0337b815194dae2a4eda3a7f7|2.97|2014-10-19 17:31:00|80.801203185414451|1|3400000031|208|35.198878721432052|0|24|47|-80.806073|7|35.106477|REGISTER BARS|0.0|1|YORK PEPPERMINT PATTIES|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00034000003303|CANDY|G1 GROCERY|-80.80146|80.801479956400485|4|3
35.17739|9df0290af7243c074c7cef3a3e573267ce0d6086|6.99|2015-01-21 18:38:00|80.801203185414451|1|1820005989|208|35.198878721432052|0|24|455|-80.806073|82|35.106477|DOMESTIC PREMIUM 12PK&>|0.0|16|MICHELOB ULTRA 6PK 12OZ  BTL|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00018200059896|DOMESTIC BEER|BEER|-80.80146|80.801479956400485|4|1
35.17739|3fc7969fd4c72bf16e057aabd56bc638d36755bd|6.99|2014-09-27 13:22:00|80.801203185414451|1|1820005989|208|35.198878721432052|0|24|455|-80.806073|82|35.106477|DOMESTIC PREMIUM 12PK&>|0.0|16|MICHELOB ULTRA 6PK 12OZ  BTL|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00018200059896|DOMESTIC BEER|BEER|-80.80146|80.801479956400485|4|1
35.17739|7c97544693133618a7cd5318726b7b69e6d904a9|6.99|2014-12-18 19:23:00|80.801203185414451|1|1820005989|208|35.198878721432052|0|24|455|-80.806073|82|35.106477|DOMESTIC PREMIUM 12PK&>|0.0|16|MICHELOB ULTRA 6PK 12OZ  BTL|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00018200059896|DOMESTIC BEER|BEER|-80.80146|80.801479956400485|4|1
35.17739|5f99565170adae83e31760a2ef07b328802b98bf|6.99|2014-10-30 16:07:00|80.801203185414451|1|1820005989|208|35.198878721432052|0|24|455|-80.806073|82|35.106477|DOMESTIC PREMIUM 12PK&>|0.0|16|MICHELOB ULTRA 6PK 12OZ  BTL|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00018200059896|DOMESTIC BEER|BEER|-80.80146|80.801479956400485|4|1
35.17739|06a38cc4419a29dec0c2b7f0aecfc2014383bfc2|6.99|2015-03-01 17:38:00|80.801203185414451|1|1820005989|208|35.198878721432052|0|24|455|-80.806073|82|35.106477|DOMESTIC PREMIUM 12PK&>|0.0|16|MICHELOB ULTRA 6PK 12OZ  BTL|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00018200059896|DOMESTIC BEER|BEER|-80.80146|80.801479956400485|4|1
35.17739|b37c734adf2e36933aab96fa4a769b722fe6c2f1|6.99|2014-11-10 14:53:00|80.801203185414451|1|1820005989|208|35.198878721432052|0|24|455|-80.806073|82|35.106477|DOMESTIC PREMIUM 12PK&>|0.0|16|MICHELOB ULTRA 6PK 12OZ  BTL|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00018200059896|DOMESTIC BEER|BEER|-80.80146|80.801479956400485|4|1
35.17739|b64be9f9789297b24e10655dde679cc829d4c3ed|6.99|2014-11-07 23:00:00|80.801203185414451|1|1820005989|208|35.198878721432052|0|24|455|-80.806073|82|35.106477|DOMESTIC PREMIUM 12PK&>|0.0|16|MICHELOB ULTRA 6PK 12OZ  BTL|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00018200059896|DOMESTIC BEER|BEER|-80.80146|80.801479956400485|4|1
35.17739|43788f5abe0557171cddabdf5d379c66f74919b9|6.99|2015-02-13 19:55:00|80.801203185414451|1|1820005989|208|35.198878721432052|0|24|455|-80.806073|82|35.106477|DOMESTIC PREMIUM 12PK&>|0.0|16|MICHELOB ULTRA 6PK 12OZ  BTL|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00018200059896|DOMESTIC BEER|BEER|-80.80146|80.801479956400485|4|1
35.17739|3c135447285329addd4b7731bce693dd05d4d781|6.99|2014-12-16 13:47:00|80.801203185414451|1|1820005989|208|35.198878721432052|0|24|455|-80.806073|82|35.106477|DOMESTIC PREMIUM 12PK&>|0.0|16|MICHELOB ULTRA 6PK 12OZ  BTL|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00018200059896|DOMESTIC BEER|BEER|-80.80146|80.801479956400485|4|1
35.17739|5117968442744ceb016c1d66810cacf643e19f19|6.99|2015-02-08 14:57:00|80.801203185414451|1|1820005989|208|35.198878721432052|0|24|455|-80.806073|82|35.106477|DOMESTIC PREMIUM 12PK&>|0.0|16|MICHELOB ULTRA 6PK 12OZ  BTL|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00018200059896|DOMESTIC BEER|BEER|-80.80146|80.801479956400485|4|1
35.17739|37f0e046412e0940af276a815c297952c0c36c23|5.59|2014-11-20 10:18:00|80.801203185414451|1|3700016943|208|35.198878721432052|0|24|403|-80.806073|69|35.106477|NFS-RUG CLEANERS|0.0|1|SWIFFER DUSTER 360 STARTER KIT|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00037000169437|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.80146|80.801479956400485|4|1
35.17739|ecded972a8b12df187ebe5dc0a123f7bd578d916|1.69|2014-12-14 13:52:00|80.801203185414451|1|1200000129|208|35.198878721432052|0|24|55|-80.806073|8|35.106477|REGULAR|0.0|23|CB DR PEPPER 20 OZ NR SINGLE|93fa34aa28db18148cf336458cbadb7ee99bce0e|1.4848191852233257|35.194272495053255|00078000082401|CARBONATED BEVERAGES|BEVERAGE|-80.80146|80.801479956400485|4|1
35.603432|d5178e476aff61d82026dfa9ccffa79c6ca9ecb4|1.25|2015-01-06 17:35:00|80.891462859624312|4||274|35.677211999422255|0|45|522|-80.995484|64|35.444064|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|94b81c3502b84162b847c537fabd1c2f8dbb5748|5.098031121419033|35.636605227883024|00204664000004|FRESH PRODUCE|PRODUCE|-80.895009|80.895200431290206|121|1
35.175855|34290a82e7d4c075cc9620a175407cef533e5c46|4.55|2014-11-04 08:44:00|80.850140887259911|4|4400002244|218|35.188411584468334|0|50|1251|-80.85753|12|35.116638|WHOLESOME COOKIES|1.05|1|NEWTONS FRUIT THIN CRNBRRY OAT|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00044000012618|COOKIES|G1 GROCERY|-80.85013|80.850139978467453|204|1
35.175855|3ee0466ed028e8f914142a9e8daa740cf615b6bc|0.5|2015-01-07 16:14:00|80.850140887259911|4||218|35.188411584468334|0|50|524|-80.85753|64|35.116638|FRESH PROD FRESH ONIONS|0.0|4|COO YELLOW ONIONS, LRG|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00204665000003|FRESH PRODUCE|PRODUCE|-80.85013|80.850139978467453|204|1
35.175855|05eb10d63f5b044862b96c5edc050cf3fb1cd2f2|2.69|2014-11-26 14:18:00|80.850140887259911|4|70935100013|218|35.188411584468334|0|50|556|-80.85753|64|35.116638|PACKAGED VEGETABLES|0.19|4|APIO BROCCOLI & CARROTS|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00709351000256|FRESH PRODUCE|PRODUCE|-80.85013|80.850139978467453|204|1
35.175855|9840f0227ba6aafd574c6424c7cfe5040ec01336|2.69|2014-12-20 16:31:00|80.850140887259911|4|70935100013|218|35.188411584468334|0|50|556|-80.85753|64|35.116638|PACKAGED VEGETABLES|0.19|4|APIO BROCCOLI & CARROTS|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00709351000256|FRESH PRODUCE|PRODUCE|-80.85013|80.850139978467453|204|1
35.175855|a45fa190715ecf73e991eb5c8e789907341bafde|3.99|2014-11-08 12:42:00|80.850140887259911|4|75928333445|218|35.188411584468334|0|50|286|-80.85753|194|35.116638|MEATLESS|0.0|5|BOCA ALL AMERICAN BURGER|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00759283673219|MEATLESS-FROZEN|FROZEN|-80.85013|80.850139978467453|204|1
35.175855|d83486e0b7581632a67e8e5a3c661a6f1ffc880f|2.89|2015-02-19 14:14:00|80.850140887259911|4|7203697887|218|35.188411584468334|0|50|61|-80.85753|9|35.116638|RTE CEREAL ADULT|0.92|1|HT CER CRUNCH GRAN RAISIN BRAN|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00072036978899|CEREAL|G1 GROCERY|-80.85013|80.850139978467453|204|1
35.175855|31b3160285271062ece611eb5bd38ba3a5eb7a7c|2.19|2014-11-28 16:48:00|80.850140887259911|4|7203608066|218|35.188411586986213|0|50|1220|-80.849471|275|35.161696|PASTA SC PREMIUM|0.0|1|HTO PASTA SC TOM BASIL|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00072036080660|PASTA SAUCES|G1 GROCERY|-80.85013|80.850132216771257|35|1
35.175855|4306dbd95a9a2b437c1e85ccc5ccc8d71f9b29b1|2.89|2015-02-16 08:48:00|80.850140887259911|4|7203655029|218|35.188411584468334|0|50|331|-80.85753|52|35.116638|NATURAL SLICED|1.22|3|HT SWISS 2% SLICES CHEESE|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00072036983954|CHEESE|DAIRY|-80.85013|80.850139978467453|204|1
35.175855|93180059eb5a72c610869df68cc1437ebba598ad|8.58|2014-12-10 16:16:00|80.850140887259911|4|2898905534|218|35.188411584468334|0|50|286|-80.85753|194|35.116638|MEATLESS|1.91|5|MSF  GRILL PRIME|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00028989055347|MEATLESS-FROZEN|FROZEN|-80.85013|80.850139978467453|204|2
35.175855|c7780fd8de595f5e26e0cf2c3bb2bfc79fb58980|8.58|2014-12-04 12:52:00|80.850140887259911|4|2898905534|218|35.188411584468334|0|50|286|-80.85753|194|35.116638|MEATLESS|1.91|5|MSF  GRILL PRIME|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00028989055347|MEATLESS-FROZEN|FROZEN|-80.85013|80.850139978467453|204|2
35.175855|cd47a54811e6d569d416c7f38126c1e721030738|1.99|2014-10-20 19:04:00|80.850140887259911|4|930000011|218|35.188411584468334|0|50|161|-80.85753|25|35.116638|PEPPERS|0.0|1|MT OLV JALAPENO DICED|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00009300000161|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.85013|80.850139978467453|204|1
35.175855|76e0ad0fea8990902331b420ac912dca3a8052b4|4.69|2014-10-19 13:51:00|80.850140887259911|4|3736300612|218|35.188411584468334|0|50|1279|-80.85753|48|35.116638|SINGLE SERVE FLAVOR|0.0|5|MICH ANGELO VEG LASAGNA|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00037363581259|FROZEN MEALS|FROZEN|-80.85013|80.850139978467453|204|1
35.175855|c189110cd3c104b078a002459365d2138f833700|4.69|2015-01-22 15:50:00|80.850140887259911|4|3736300612|218|35.188411584468334|0|50|1279|-80.85753|48|35.116638|SINGLE SERVE FLAVOR|0.0|5|MICH ANGELO VEG LASAGNA|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00037363581259|FROZEN MEALS|FROZEN|-80.85013|80.850139978467453|204|1
35.175855|72bd7e91b47e36dc56e0204ae8fbac710b5bc8f9|4.69|2015-03-03 14:08:00|80.850140887259911|4|3736300612|218|35.188411584468334|0|50|1279|-80.85753|48|35.116638|SINGLE SERVE FLAVOR|0.0|5|MICH ANGELO VEG LASAGNA|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00037363581259|FROZEN MEALS|FROZEN|-80.85013|80.850139978467453|204|1
35.175855|0e63944170d7b9a5b55eeb14d1bf6a36ac9fc0ff|4.69|2014-09-11 15:43:00|80.850140887259911|4|3736300612|218|35.188411584468334|0|50|1279|-80.85753|48|35.116638|SINGLE SERVE FLAVOR|1.35|5|MICH ANGELO VEG LASAGNA|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00037363581259|FROZEN MEALS|FROZEN|-80.85013|80.850139978467453|204|1
35.175855|1bccaf342354a534b27c836d3d6440fa9640477f|4.69|2014-10-07 16:09:00|80.850140887259911|4|3736300612|218|35.188411584468334|0|50|1279|-80.85753|48|35.116638|SINGLE SERVE FLAVOR|1.35|5|MICH ANGELO VEG LASAGNA|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00037363581259|FROZEN MEALS|FROZEN|-80.85013|80.850139978467453|204|1
35.175855|42ffd4f98394c8b6b34e219e62efd493b1fab536|7.7|2014-12-29 12:31:00|80.850140887259911|4|4812127620|218|35.188411584468334|0|50|1037|-80.85753|164|35.116638|ENGLISH MUFFINS|1.92|7|THOMAS 100% WHEAT ENG MUFN PP|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00048121184070|BREAKFAST|COMMERCIAL BAKERY|-80.85013|80.850139978467453|204|2
35.175855|6bb154bcef360d0bbaeea2dc87c6a2cfe684984f|3.99|2014-11-20 15:22:00|80.850140887259911|4|2840007134|218|35.188411584468334|0|50|204|-80.85753|31|35.116638|TORTILLA CHIPS|0.0|1|SIMPLY TOSTITOS BLUE|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00028400071345|SNACKS|G1 GROCERY|-80.85013|80.850139978467453|204|1
35.175855|28779a08987f5574e41fbbfe3d9004c712e280b7|3.99|2015-01-01 09:34:00|80.850140887259911|4|2840007134|218|35.188411584468334|0|50|204|-80.85753|31|35.116638|TORTILLA CHIPS|0.0|1|SIMPLY TOSTITOS BLUE|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00028400071345|SNACKS|G1 GROCERY|-80.85013|80.850139978467453|204|1
35.175855|fa33c597c3b4eb9bf5f74f7c599b91cee38473e4|1.69|2015-01-03 12:20:00|80.850140887259911|4|7203633026|218|35.188411584468334|0|50|200|-80.85753|31|35.116638|MICROWAVE POPCORN|0.0|1|HT MICROWAVE POPCORN|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00072036330260|SNACKS|G1 GROCERY|-80.85013|80.850139978467453|204|1
35.175855|7994c2617392bcdd1637b9cf40f93af32d3761cb|0.67|2015-02-05 15:22:00|80.850140887259911|4|7203641111|218|35.188411584468334|0|50|242|-80.85753|39|35.116638|CANNED BEANS|0.0|1|HT PEAS BLACKEYE|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00072036411143|VEGETABLES-CAN/JAR|G1 GROCERY|-80.85013|80.850139978467453|204|1
35.175855|351103b59bb1f84bc9168337018368c5bf29db72|8.99|2014-09-14 16:53:00|80.850140887259911|4|8308590302|218|35.188411584468334|0|50|9957|-80.85753|886|35.116638|NFS-PREM-OTHER RED|0.0|13|RUFFINO CHIANTI|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00083085903022|PREMIUM ($8-$10.99)|WINE|-80.85013|80.850139978467453|204|1
35.175855|4ffc18bccfb8cb134f1a4897f4799f92163eb60d|8.58|2015-01-31 14:37:00|80.850140887259911|4|2840006399|218|35.188411584468334|0|50|204|-80.85753|31|35.116638|TORTILLA CHIPS|2.14|1|TOSTITOS HINT OF LIME|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00028400064040|SNACKS|G1 GROCERY|-80.85013|80.850139978467453|204|2
35.175855|0267346e8c65ad4129741f82ec7bb4c454b1d9e6|3.99|2014-11-26 16:30:00|80.850140887259911|4|7203602701|218|35.188411584468334|0|50|1878|-80.85753|435|35.116638|HUMMUS|0.5|6|FFM ARTISAN RED PEPPER HUMMUS|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00072036027030|SALADS|DELI|-80.85013|80.850139978467453|204|1
35.175855|9391551b40af62e34e01b9c40201c947860ff4e5|2.55|2015-01-27 18:39:00|1.4094857484078087|4|7203636026|218|0.6139344869541099|0|26|54|-80.85013|8|35.175855|DIET|0.25|23|HT DIET TONIC WITH QUININE|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|0.61471665291522548|00072036360410|CARBONATED BEVERAGES|BEVERAGE|-80.85013|1.4111009691654428|218|3
35.175855|76c527e7e8620ee7b6c7e832c9ee4ec5d30b3235|1.7|2014-11-29 15:16:00|80.850140887259911|4|7203636026|218|35.188411584468334|0|50|54|-80.85753|8|35.116638|DIET|0.7|23|HT DIET TONIC WITH QUININE|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00072036360410|CARBONATED BEVERAGES|BEVERAGE|-80.85013|80.850139978467453|204|2
35.175855|aca69d1ecf207e5cf2da8ceb9a61b441f7ed8a0c|1.7|2014-10-12 14:30:00|80.850140887259911|4|7203636026|218|35.188411586463133|0|50|54|-80.844274|8|35.204336|DIET|0.0|23|HT DIET TONIC WITH QUININE|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00072036360410|CARBONATED BEVERAGES|BEVERAGE|-80.85013|80.850134957668416|61|2
35.175855|5ea60d3334f89fdca8902cf57a636bcb649d7cd3|2.55|2015-01-15 13:21:00|80.850140887259911|4|7203636026|218|35.188411584468334|0|50|54|-80.85753|8|35.116638|DIET|0.0|23|HT DIET TONIC WITH QUININE|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00072036360410|CARBONATED BEVERAGES|BEVERAGE|-80.85013|80.850139978467453|204|3
35.175855|ad52861782f7386e9100ac8da88a2b052e4d504f|1.7|2014-09-30 16:54:00|80.850140887259911|4|7203636026|218|35.188411584468334|0|50|54|-80.85753|8|35.116638|DIET|0.0|23|HT DIET TONIC WITH QUININE|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00072036360410|CARBONATED BEVERAGES|BEVERAGE|-80.85013|80.850139978467453|204|2
35.175855|cbe5429e4db37fb29f600963cbbe5964c6e67dea|1.7|2015-02-07 10:52:00|80.850140887259911|4|7203636026|218|35.188411584468334|0|50|54|-80.85753|8|35.116638|DIET|0.0|23|HT DIET TONIC WITH QUININE|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00072036360410|CARBONATED BEVERAGES|BEVERAGE|-80.85013|80.850139978467453|204|2
35.175855|1f856f2ffc40c408d0030d87603efedb0335594d|0.69|2014-09-21 18:40:00|80.850140887259911|4|71070842240|218|35.188411584468334|0|50|580|-80.85753|136|35.116638|OTHER MERCH DRESSINGS|0.0|4|ORGANIC BALSAMIC VIN DRESSING|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00710708422409|OTHER MERCHANDISE|PRODUCE|-80.85013|80.850139978467453|204|1
35.175855|20f231a1bb6b0bea12b47dafbf7040274d14c232|4.79|2014-12-17 20:38:00|80.850140887259911|4|18685200031|218|35.188411584468334|0|50|275|-80.85753|45|35.116638|SUPER PREMIUM ICE CREAM|0.0|5|TALENTI  BLACK RASB.CHO.CHP. .|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00186852000617|ICE CREAM|FROZEN|-80.85013|80.850139978467453|204|1
35.175855|0fb3fa784226df5ced600c534e15475eb38ef813|5.69|2014-11-12 14:57:00|80.850140887259911|4|1450000711|218|35.188411584468334|0|50|1274|-80.85753|50|35.116638|BAG VEG PROTEIN|0.0|5|BE VOILA SHRIMP SCAMPI|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00014500011725|VEGETABLES-FROZEN|FROZEN|-80.85013|80.850139978467453|204|1
35.175855|d64d88e89cc77303df24fbcc07f42f6cb15ee992|1.79|2014-11-14 09:00:00|1.4094857484078087|4|7203663157|218|0.6139344869541099|0|26|1134|-80.85013|57|35.175855|CARTON MILK|0.0|3|HARRIS TEETER FF SKIM MILK|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|0.61471665291522548|00072036631565|MILK|DAIRY|-80.85013|1.4111009691654428|218|1
35.175855|c4c815c1d73e668dcded4a92623c74f2ac5e5b80|3.49|2014-12-27 11:16:00|1.4094857484078087|4|4589307223|218|0.6139344869541099|0|26|3198|-80.85013|1015|35.175855|HAND & BODY PRICE|0.0|17|SUAVE VIT E LOTION|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|0.61471665291522548|00045893072253|HAND & BODY LOTION/SUN CARE|HBC|-80.85013|1.4111009691654428|218|1
35.175855|5a80718f041088295ec3e36a2ede2e915c459518|7.98|2014-12-09 19:09:00|80.850140887259911|4|3400008752|218|35.188411584468334|0|50|46|-80.85753|7|35.116638|PKG CHOC|0.0|1|MOUNDS SNACK BARS|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00034000020102|CANDY|G1 GROCERY|-80.85013|80.850139978467453|204|2
35.175855|c89e15f262d349e8be6e509338b914c9093c3c9d|3.99|2015-01-20 19:36:00|80.850140887259911|4|3400008752|218|35.188411584468334|0|50|46|-80.85753|7|35.116638|PKG CHOC|0.0|1|MOUNDS SNACK BARS|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00034000020102|CANDY|G1 GROCERY|-80.85013|80.850139978467453|204|1
35.175855|d051a25a26eca7addb46198018fcf3efc56adf1a|3.99|2014-12-21 11:37:00|80.850140887259911|4|7020052202|218|35.188411584468334|0|50|582|-80.85753|136|35.116638|DIPS-REFRIG. & DRY|0.99|4|MARZ RANCH VEGGIE DIP|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00070200522008|OTHER MERCHANDISE|PRODUCE|-80.85013|80.850139978467453|204|1
35.175855|63a8de99708f8704cfb2b46d07f52c0b117b2a75|13.99|2015-01-21 19:29:00|80.850140887259911|4|8834510053|218|35.188411584468334|0|50|459|-80.85753|83|35.116638|IMPORT BEER|0.0|16|NEWCASTLE 12PK 12OZ BTL|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00088345100531|IMPORT BEER|BEER|-80.85013|80.850139978467453|204|1
35.175855|c541342286a217d5c2474eb9c06b316168496969|4.99|2014-12-24 09:23:00|80.850140887259911|4|7336070341|218|35.188411584468334|0|50|30|-80.85753|4|35.116638|CARBONATED WATER|0.0|1|LACROIX WTR CRAN RSP 12PK|9987f22e8e8dc6794b75e0bc0bddb5bb2dcba1f6|0.8676298467081957|35.186025810841215|00073360323416|BOTTLED WATER|G1 GROCERY|-80.85013|80.850139978467453|204|1
35.444064|677d2be2a35a5fce74596f37c5a2a3fcc88a54ae|6.99|2015-02-28 16:40:00|1.4102725052409182|4|7203627074|121|0.6186156170875914|0|1|152|-80.995484|24|35.444064|NFS-CAT FOOD DRY|0.0|1|HT YOURPET 4 FLAVOR CAT FOOD|9a21f9e0433081fdad6b71eabdc616d46b30304a|2.1745380689868767|0.61833652052202714|00072036270740|PET FOOD/SUPPLIES|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|8a09cd6c5b9b5baf8c4dbf146e2680c87613c796|3.99|2015-03-04 18:45:00|1.4102725052409182|4|1600027534|121|0.6186156170875914|0|1|81|-80.995484|9|35.444064|RTE CEREAL KIDS|0.0|1|GM LUCKY CHARMS  11.5OZ|9a21f9e0433081fdad6b71eabdc616d46b30304a|2.1745380689868767|0.61833652052202714|00016000275348|CEREAL|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|c09a3d9f0997ef12cfc488c4b11d2a82a647566b|3.49|2015-03-02 17:25:00|1.4102725052409182|4|88491212971|121|0.6186156170875914|0|1|81|-80.995484|9|35.444064|RTE CEREAL KIDS|0.0|1|POST PEBBLES FRUITY|9a21f9e0433081fdad6b71eabdc616d46b30304a|2.1745380689868767|0.61833652052202714|00884912129710|CEREAL|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|73123c4cb4c4bf5a3143ca386e72bff50fac3eac|3.49|2014-11-15 17:52:00|1.4102725052409182|4|88491212971|121|0.6186156170875914|0|1|81|-80.995484|9|35.444064|RTE CEREAL KIDS|0.0|1|POST PEBBLES FRUITY|9a21f9e0433081fdad6b71eabdc616d46b30304a|2.1745380689868767|0.61833652052202714|00884912129710|CEREAL|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|d06ed4a24dd89e95d97736bfb12f6ebcb6584770|6.57|2015-01-02 18:43:00|80.995508130988839|4|7203698771|121|35.475534533245657|0|40|176|-80.8955|72|35.4437|NFS-DISPOSE CUPS|0.0|1|YH FOAM CUPS 10 OZ|9a21f9e0433081fdad6b71eabdc616d46b30304a|2.1745380689868767|35.466476270328783|00072036987716|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.995484|80.995501392718978|272|3
35.444064|aa5a72529577a4aec01634ec8f1882f2c5284f2f|11.99|2014-09-27 19:33:00|1.4102725052409182|4|71981200314|121|0.6186156170875914|0|1|5861|-80.995484|1538|35.444064|COLANDERS|0.0|18|"OXO 8"" STRAINER"|9a21f9e0433081fdad6b71eabdc616d46b30304a|2.1745380689868767|0.61833652052202714|00719812003146|KITCHEN GADGETS|GM|-80.995484|1.413637875046387|121|1
35.17335|8a7211914c93e3933b18e067a1a3b3010b9f89c8|3.59|2014-11-23 14:05:00|80.709059419360486|4|4900006520|174|35.192035539366074|0|31|54|-80.739|8|35.141204|DIET|0.6|23|COKE LIFE 12 OZ 6PK CANS|9a958617c18962a2c524840f610ee4e85097e55b|1.2911257893178383|35.187384292804154|00049000065206|CARBONATED BEVERAGES|BEVERAGE|-80.70901|80.709020763162584|171|1
35.17335|df8318585b3164719a573661fd775d8ae3fd85fc|0.85|2015-01-27 14:25:00|80.709059419360486|4||174|35.192035539366074|0|31|522|-80.739|64|35.141204|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|9a958617c18962a2c524840f610ee4e85097e55b|1.2911257893178383|35.187384292804154|00204664000004|FRESH PRODUCE|PRODUCE|-80.70901|80.709020763162584|171|1
35.17335|2dae5f454cf69e83d1e885969bec4f1a50b6a4ed|3.19|2015-02-27 20:24:00|80.709059419360486|4|5000062231|174|35.192035539366074|0|31|326|-80.739|54|35.141204|COOKIES/BROWNIES-REFRIGERATED|0.0|3|NESTLE WHT CHOC CHIP MACADAMIA|9a958617c18962a2c524840f610ee4e85097e55b|1.2911257893178383|35.187384292804154|00050000009237|DOUGH PRODUCTS|DAIRY|-80.70901|80.709020763162584|171|1
35.17335|de1194ba81d51381599c1d8a32efd9eadd6ca1aa|2.29|2014-12-15 20:26:00|80.709059419360486|4|7800023046|174|35.192035540108023|0|31|55|-80.80146|8|35.17739|REGULAR|1.29|23|CHERRY SUNDROP 2 LTR|9a958617c18962a2c524840f610ee4e85097e55b|1.2911257893178383|35.187384292804154|00078000232462|CARBONATED BEVERAGES|BEVERAGE|-80.70901|80.70901862195754|208|1
35.17335|86bb7a641aca519a6b0a915f2d7473cb19f077df|5.99|2015-02-13 17:58:00|80.709059419360486|4|7756725423|174|35.192035539366074|0|31|252|-80.739|45|35.141204|PREMIUM ICE CREAM|2.99|5|BREYERS BUTTER PECAN I/C|9a958617c18962a2c524840f610ee4e85097e55b|1.2911257893178383|35.187384292804154|00077567254405|ICE CREAM|FROZEN|-80.70901|80.709020763162584|171|1
35.17335|d0dc3fd9b7198a6e27cc194cc8166222014e0b21|2.99|2015-01-09 19:03:00|80.709059419360486|4|8201110007|174|35.192035539046451|0|31|1250|-80.709466|12|35.124987|SPECIALTY COOKIES|0.0|1|MURRAY GINGER SNAPS|9a958617c18962a2c524840f610ee4e85097e55b|1.2911257893178383|35.187384292804154|00082011100078|COOKIES|G1 GROCERY|-80.70901|80.709021564038693|157|1
35.17335|6df88ceee9de5c0864f9ee4de349fb94695cc49f|4.59|2014-11-08 17:11:00|80.709059419360486|4|5000088600|174|35.192035539366074|0|31|341|-80.739|57|35.141204|CREAMERS|2.09|3|I/O COFFEEMATE PUMPKIN SPICE|9a958617c18962a2c524840f610ee4e85097e55b|1.2911257893178383|35.187384292804154|00050000886005|MILK|DAIRY|-80.70901|80.709020763162584|171|1
35.17335|fd545cf4d115bf35e15e72c7eae75b5ceb23bdff|3.34|2015-01-05 20:22:00|80.709059419360486|4|7203643010|174|35.192035539366074|0|31|252|-80.739|45|35.141204|PREMIUM ICE CREAM|0.0|5|HT PREM CHOCOLATE IC|9a958617c18962a2c524840f610ee4e85097e55b|1.2911257893178383|35.187384292804154|00072036430113|ICE CREAM|FROZEN|-80.70901|80.709020763162584|171|1
35.17335|7da8086a47b3dc23962f85701f242c1df00bb6d5|2.89|2015-03-04 21:04:00|1.4094857484078087|4|7203603037|174|0.6138907664563474|0|26|1253|-80.70901|12|35.17335|ALL OTHER COOKIES|0.39|1|HT GINGER SNAPS|9a958617c18962a2c524840f610ee4e85097e55b|1.2911257893178383|0.61471665291522548|00072036030368|COOKIES|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|f68c6033625caf82615985dcc1eacd9f0b4c16d4|0.79|2014-12-24 17:42:00|1.4094857484078087|4|7203641055|174|0.6138907664563474|0|26|257|-80.70901|39|35.17335|TOMATOES|0.0|1|HT TOMATOES PETITE DICED|9a958617c18962a2c524840f610ee4e85097e55b|1.2911257893178383|0.61471665291522548|00072036410726|VEGETABLES-CAN/JAR|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|b8bcdf5e0997b9ea36581f73e39a993c9856cf24|2.99|2015-02-28 18:16:00|80.709059419360486|4|67791671581|174|35.192035539366074|0|31|7002|-80.739|1600|35.141204|VALENTINE PARTY GOOD/DECORTN|2.24|18|I/O VAL PRNT BCKET W/RIBN HNDL|9a958617c18962a2c524840f610ee4e85097e55b|1.2911257893178383|35.187384292804154|00677916715818|SEASONAL MERCHANDISE|GM|-80.70901|80.709020763162584|171|1
35.17335|72220d87caf8b3b55dbdfd6a8bce99218d997229|5.49|2015-01-16 16:58:00|80.709059419360486|4|73866500003|174|35.192035540108023|0|31|1511|-80.80146|65|35.17739|CHARCOAL/L NFS-FIREWOOD|0.0|1|CUSTIS BUNDLED FIREWOOD|9a958617c18962a2c524840f610ee4e85097e55b|1.2911257893178383|35.187384292804154|00738665000034|CHARCOAL/LOGS/ACCESSORIES|G1 GROCERY|-80.70901|80.70901862195754|208|1
35.17335|baf4447452b4b0c483514208010d111b1d84b371|1.69|2014-10-25 13:49:00|1.4094857484078087|4|4430010632|174|0.6138907664563474|0|26|1212|-80.70901|272|35.17335|HISP BEANS/PEPPERS|0.69|1|ROSARITA REFRIED BEANS TRAD|9a958617c18962a2c524840f610ee4e85097e55b|1.2911257893178383|0.61471665291522548|00044300106321|HISPANIC PREP. FOODS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|da477994fe7ed689d84fd19f441bfcd7d045b5d7|3.19|2014-11-21 20:28:00|1.4094857484078087|4|2340036004|174|0.6138907664563474|0|26|393|-80.70901|68|35.17335|NFS-AIR FRESHENERS|0.69|1|RENUZIT SUPER ODOR BREEZE|9a958617c18962a2c524840f610ee4e85097e55b|1.2911257893178383|0.61471665291522548|00023400360437|FRESHENERS/DEODORIZERS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|775d28d1055c05b9947e48296b0f193f4134d92c|2.99|2015-02-14 18:31:00|80.709059419360486|4|3485602884|174|35.192035539366074|0|31|1200|-80.739|6|35.141204|FRUIT SNACKS|0.0|1|WELCH'S FRUIT SNACKS MIX FRUIT|9a958617c18962a2c524840f610ee4e85097e55b|1.2911257893178383|35.187384292804154|00034856028888|BREAKFAST FOODS|G1 GROCERY|-80.70901|80.709020763162584|171|1
35.412407|2dd716b5e07790cbc631b18daa2780a26f2d44c8|6.79|2014-11-15 12:27:00|1.4102725052409182|4|2500005838|68|0.6180630982062877|0|1|55|-80.662946|8|35.412407|REGULAR|0.0|23|MINUTE MAID L'ADE 12OZ 12PK CN|9b262db65caaf7ba34428646a041c88af769ee95|3.131160616213855|0.61833652052202714|00025000058387|CARBONATED BEVERAGES|BEVERAGE|-80.662946|1.40783399205839|68|1
35.412407|8879fe7dbd9d33b585fee28400c218c50483d77e|5.98|2014-10-04 19:37:00|1.4102725052409182|4|3620021922|68|0.6180630982062877|0|1|1219|-80.662946|275|35.412407|PASTA SC CORE|0.0|1|BERTOLLI SC ALFREDO GARLIC|9b262db65caaf7ba34428646a041c88af769ee95|3.131160616213855|0.61833652052202714|00036200219195|PASTA SAUCES|G1 GROCERY|-80.662946|1.40783399205839|68|2
35.23102|0643babf8812d793ec3e9ffcd72caf75b1420e08|1.49|2014-12-14 12:59:00|80.843945456961976|4|7203670302|205|35.239786191835215|0|59|728|-80.810056|72|35.219587|NFS-PLASTIC FLATWARE|0.49|1|YH OCCASIONS FS FORKS|9c98831eb38af2cc1c78c82fb474f7f8eedd18c2|0.6057226865682583|35.232478750868765|00072036703019|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.8438|80.843800365254637|401|1
35.23102|b6873dc11017714984fd5e2327ca38f89a76f420|1.99|2014-12-08 18:51:00|1.4094857484078087|4||205|0.6148972978359727|0|26|535|-80.8438|64|35.23102|FRESH GREENS|0.0|4|SPINACH, BUNCH (RPC)|9c98831eb38af2cc1c78c82fb474f7f8eedd18c2|0.6057226865682583|0.61471665291522548|00204090000005|FRESH PRODUCE|PRODUCE|-80.8438|1.4109904898237917|205|1
35.23102|4d2a041237ce4b1e16a4ee0730f4585d4a7fc781|3.35|2014-10-18 12:45:00|80.843945456961976|4||205|35.239786191835215|0|59|500|-80.810056|64|35.219587|FRESH APPLES|1.26|4|HONEY CRISP APPLE|9c98831eb38af2cc1c78c82fb474f7f8eedd18c2|0.6057226865682583|35.232478750868765|00233283000003|FRESH PRODUCE|PRODUCE|-80.8438|80.843800365254637|401|1
35.23102|3049b6f5700de73b33880e853665c2150c7f0777|7.98|2014-11-14 16:03:00|1.4094857484078087|4|20405400000|205|0.6148972978359727|0|26|504|-80.8438|64|35.23102|FRESH BERRIES|1.99|4|RED RASPBERRIES 6 OZ|9c98831eb38af2cc1c78c82fb474f7f8eedd18c2|0.6057226865682583|0.61471665291522548|00715756100019|FRESH PRODUCE|PRODUCE|-80.8438|1.4109904898237917|205|2
35.23102|91e852f999d0544eb96cb0c0e4b4371b12c4d58b|3.49|2014-09-13 18:51:00|1.4094857484078087|4|7203695248|205|0.6148972978359727|0|26|1611|-80.8438|371|35.23102|PITA'S AND FLAT BREADS|0.99|14|FFM WHEAT PITA POCKET|9c98831eb38af2cc1c78c82fb474f7f8eedd18c2|0.6057226865682583|0.61471665291522548|00072036952516|BREAD|BAKERY|-80.8438|1.4109904898237917|205|1
35.23102|566ad816a55da3ba684e298376bb00958b9fa48a|1.89|2014-10-20 17:45:00|1.4094857484078087|4|5100005977|205|0.6148972978359727|0|26|212|-80.8438|33|35.23102|CONDENSED SOUP|0.22|1|CAMP HLTHY REQ CREAM MUSHROOM|9c98831eb38af2cc1c78c82fb474f7f8eedd18c2|0.6057226865682583|0.61471665291522548|00051000060075|SOUP|G1 GROCERY|-80.8438|1.4109904898237917|205|1
35.23102|6e0a8a47c9265feb3fb41e43a8c7fc83181e2db8|4.99|2014-12-14 13:55:00|1.4094857484078087|4|71575620002|205|0.6148972978359727|0|26|504|-80.8438|64|35.23102|FRESH BERRIES|0.0|4|STRAWBERRIES 1LB CLAM|9c98831eb38af2cc1c78c82fb474f7f8eedd18c2|0.6057226865682583|0.61471665291522548|00665290001184|FRESH PRODUCE|PRODUCE|-80.8438|1.4109904898237917|205|1
35.23102|6daaff798f8dc8598146c2e3332540ebbded9d48|3.58|2014-12-14 13:56:00|1.4094857484078087|4|5100001047|205|0.6148972978359727|0|26|212|-80.8438|33|35.23102|CONDENSED SOUP|0.24|1|CAMP COND 25% LS CRM MUSHROOM|9c98831eb38af2cc1c78c82fb474f7f8eedd18c2|0.6057226865682583|0.61471665291522548|00051000166814|SOUP|G1 GROCERY|-80.8438|1.4109904898237917|205|2
35.41832|cc2a0c6f6e8080645cbaf0190731500e23292c8e|4.69|2014-10-10 21:42:00|80.749667378538092|4|4900002468|190|35.485348167703414|0|3|54|-80.737839|8|35.297134|DIET|1.19|23|DIET COKE .5 LITER/6 PK.|9d78b966e64db8ad75c69a1189d9076c6f16c118|4.631487974860437|35.465179900649026|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.746334|80.746434487896622|258|1
35.41832|1f60da3b9c0f2852d98668ecbe4ced161a9c7da2|7.99|2015-01-20 19:31:00|80.749667378538092|4|1820017993|190|35.485348167703414|0|3|458|-80.737839|82|35.297134|CRAFT BEER|0.0|16|SHOCK TOP SEASONAL 6PK|9d78b966e64db8ad75c69a1189d9076c6f16c118|4.631487974860437|35.465179900649026|00018200179938|DOMESTIC BEER|BEER|-80.746334|80.746434487896622|258|1
35.41832|da9e5b42a360c10b9c9c8307b413b390b5f36bb6|4.85|2014-12-10 18:45:00|80.749667378538092|4|7790011553|190|35.485348167703414|0|3|361|-80.737839|105|35.297134|BREAKFAST SAUSAGE|1.51|19|JIMMY DEAN SAGE SAUSAGE|9d78b966e64db8ad75c69a1189d9076c6f16c118|4.631487974860437|35.465179900649026|00077900116339|BREAKFAST SAUSAGE|CASE READY MEATS|-80.746334|80.746434487896622|258|1
35.41832|3d6a4d3beddf8f85601ce7d4a2feb3f080f6cef3|3.39|2014-10-22 18:30:00|80.749667378538092|4|5000062261|190|35.485348167703414|0|3|326|-80.737839|54|35.297134|COOKIES/BROWNIES-REFRIGERATED|0.39|3|I/O NES SCOTCHIE|9d78b966e64db8ad75c69a1189d9076c6f16c118|4.631487974860437|35.465179900649026|00050000622610|DOUGH PRODUCTS|DAIRY|-80.746334|80.746434487896622|258|1
35.41832|26acb07824b51980a9a39dfb096f870603c4747d|7.19|2014-10-31 16:19:00|80.749667378538092|4|7080004118|190|35.485348216650557|0|3|358|-80.762919|100|35.442529|REGULAR BACON|3.6|19|SMITHFIELD CHERRYWOOD BACON|9d78b966e64db8ad75c69a1189d9076c6f16c118|4.631487974860437|35.465179900649026|00070800041268|BACON|CASE READY MEATS|-80.746334|80.746348474010929|471|1
35.41832|e83d8ee7c025aa421da9a9c91dfdf47d3c084962|12.99|2014-11-26 11:18:00|80.749667378538092|4|4460031182|190|35.485348167703414|0|3|385|-80.737839|65|35.297134|NFS-CHARCOAL|1.81|1|KINGSFORD CHARCOAL|9d78b966e64db8ad75c69a1189d9076c6f16c118|4.631487974860437|35.465179900649026|00044600304519|CHARCOAL/LOGS/ACCESSORIES|G1 GROCERY|-80.746334|80.746434487896622|258|1
35.41832|316eb4751ab3b371aefbd18ea8347e534c9ac90e|2.35|2014-12-23 22:29:00|80.749667378538092|4|2150004209|190|35.485348167703414|0|3|71|-80.737839|11|35.297134|GROC CONDIMENTS MARINADE|0.0|1|LAWRYS MARINADE STEAK & CHOP|9d78b966e64db8ad75c69a1189d9076c6f16c118|4.631487974860437|35.465179900649026|00021500042178|CONDIMENTS|G1 GROCERY|-80.746334|80.746434487896622|258|1
35.41832|11be5e547b7fa03ac9aa243425814b5b1f58c221|11.99|2014-10-11 20:27:00|80.749667378538092|4|7203663048|190|35.485348167703414|0|3|297|-80.737839|49|35.297134|GROUND BEEF|1.0|2|93% LEAN GROUND BEEF 2 LB|9d78b966e64db8ad75c69a1189d9076c6f16c118|4.631487974860437|35.465179900649026|00072036630483|BEEF|MEAT|-80.746334|80.746434487896622|258|1
35.41832|a94aa0b6a05744e0ba1695499b02156e139c6559|2.87|2014-10-24 18:38:00|80.749667378538092|4|7203602031|190|35.485348167703414|0|3|387|-80.737839|65|35.297134|NFS-REMAIN CHAR/LOGS/ACC|0.0|1|HT LIGHTER FLUID CAN|9d78b966e64db8ad75c69a1189d9076c6f16c118|4.631487974860437|35.465179900649026|00072036020314|CHARCOAL/LOGS/ACCESSORIES|G1 GROCERY|-80.746334|80.746434487896622|258|1
35.41832|0ceede84be5aa132442ead987291c13218af8a4f|7.19|2014-11-21 18:19:00|80.749667378538092|4|7080004118|190|35.485348167703414|0|3|845|-80.737839|100|35.297134|NATURAL/ORGANIC BACON|3.6|19|SMFD NATURAL HICKORY BACON|9d78b966e64db8ad75c69a1189d9076c6f16c118|4.631487974860437|35.465179900649026|00070800023103|BACON|CASE READY MEATS|-80.746334|80.746434487896622|258|1
35.41832|af8593df08ec21f5001d92bd8cbad642c3f28ddd|12.99|2014-11-14 21:01:00|80.749667378538092|4|8470409132|190|35.485348031672174|0|3|9983|-80.810056|889|35.219587|NFS-SPARKLING|0.0|13|CB-KORBEL BRUT|9d78b966e64db8ad75c69a1189d9076c6f16c118|4.631487974860437|35.465179900649026|00084704091328|SPARKLING|WINE|-80.746334|80.746527852685446|401|1
35.41832|f6e2b96a175ed6a77cb99e86fb35bc757a06d6e7|2.49|2015-01-26 08:23:00|1.4102725052409182|4|1200001643|190|0.6181662995249579|0|1|97|-80.746334|8|35.41832|ENERGY DRINKS|0.5|23|MTN DEW AMP TALL  BOY|9d78b966e64db8ad75c69a1189d9076c6f16c118|4.631487974860437|0.61833652052202714|00012000016431|CARBONATED BEVERAGES|BEVERAGE|-80.746334|1.409289387215043|190|1
35.103409|5e862da6eaf9169fde69a2f56841c8d4153c1850|11.99|2014-09-25 16:48:00|1.4132775322775095|4|2301286481|88|0.6126700657242101|0|58|1477|-80.992182|485|35.103409|SUSHI HYBRID|0.0|6|"CHEF SAMPLER ""A"""|9f081a637214777df021a9077adc6364bb79a5be|3.902154818395855|0.61177642288969325|00023012864811|SUSHI|DELI|-80.992182|1.413580244274486|88|1
35.103409|e9a81a19321ee4d2e0af4495609a87b268a100d7|1.0|2014-11-25 12:28:00|1.4132775322775095|4|4000000435|88|0.6126700657242101|0|58|47|-80.992182|7|35.103409|REGISTER BARS|0.2|1|(FE)DOVE MILK CHOC SINGLES|9f081a637214777df021a9077adc6364bb79a5be|3.902154818395855|0.61177642288969325|00040000459842|CANDY|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|b4f09d301f0842b459673577d4c22183cfac4ba7|2.79|2014-10-19 14:16:00|1.4132775322775095|3|1800065680|88|0.6126700657242101|0|58|1270|-80.992182|41|35.103409|SWEET BREAKFAST|0.0|5|PILLSBURY TSTR STRDL BLUEBERRY|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00018000655304|BREAKFAST FOODS FROZEN|FROZEN|-80.992182|1.413580244274486|88|1
35.103409|2ee73994ea14754273b246395daaf52e3962dfda|10.76|2015-02-16 10:56:00|1.4132775322775095|3|1450000253|88|0.6126700657242101|0|58|1272|-80.992182|50|35.103409|BAG VEG STEAM|2.76|5|BE STEAMFRESH PREM GRN BEANS|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00014500011572|VEGETABLES-FROZEN|FROZEN|-80.992182|1.413580244274486|88|4
35.103409|ded3aac93bfa0d7eeca78d3f0cf754363ba29df4|12.99|2014-12-12 19:30:00|1.4132775322775095|3|8769200129|88|0.6126700657242101|0|58|458|-80.992182|82|35.103409|CRAFT BEER|0.0|16|SAM ADAMS REBEL IPA 12PK BTL|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00087692001294|DOMESTIC BEER|BEER|-80.992182|1.413580244274486|88|1
35.103409|d808fd2d06106be5d6040ab8d17f18b5c6f6ca09|3.49|2014-09-14 19:45:00|1.4132775322775095|3|2840023981|88|0.6126700657242101|0|58|203|-80.992182|31|35.103409|CHEESE SNACKS|0.99|1|CHEETOS JUMBO PUFFS|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00028400239875|SNACKS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|5c490f99ab06640f05562db4c7a0aa99adf61fe7|3.29|2015-01-05 21:17:00|1.4132775322775095|3|2840004768|88|0.6126700657242101|0|58|202|-80.992182|31|35.103409|PRETZELS|0.29|1|ROLD GOLD 3 CHEESE PRETZEL THN|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00028400232043|SNACKS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|8e73874d083399fccc7ec3122eb8a07a121abf87|3.98|2014-11-23 13:59:00|1.4132775322775095|3|3900004504|88|0.6126700657242101|0|58|114|-80.992182|14|35.103409|PUMPKIN|0.4|1|LIBBY SOLID PACK PUMPKIN|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00039000045049|DESSERTS/GELS/SYRUPS|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|fcba8a6861dd38cb07d5494c011a9ed7b20a291b|6.98|2015-01-26 18:59:00|1.4132775322775095|3|7017715419|88|0.6126700657242101|0|58|233|-80.992182|37|35.103409|BLACK TEA|0.49|1|TWININGS TEA BLK IRISH BREAKFS|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00070177154240|TEA|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|254afe11a5d8d75fdc072f34ba2ef4cba46b27b3|2.29|2015-01-10 16:59:00|1.4132775322775095|3|5210004620|88|0.6126700657242101|0|58|18|-80.992182|3|35.103409|CAKE DECORATIONS & ICING|0.0|1|CAKE MATE BLACK GEL|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00052100046419|BAKING SUPPLIES|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|1d9f757756483978a9e52e16f13d50b491bfb287|6.79|2015-02-06 17:16:00|1.4132775322775095|3|5233633181|88|0.6126700657242101|0|58|3589|-80.992182|1050|35.103409|HAIR STYLING GLUE|1.8|17|GOT 2B GLUED SPIKE GEL 33145|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00052336331457|HAIR STYLING|HBC|-80.992182|1.413580244274486|88|1
35.103409|f2e27076b12ba9d71e26c4a9cbb66ef40c67ace9|6.79|2014-11-09 09:55:00|1.4132775322775095|3|5233633181|88|0.6126700657242101|0|58|3589|-80.992182|1050|35.103409|HAIR STYLING GLUE|1.0|17|GOT 2B GLUED SPIKE GEL 33145|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00052336331457|HAIR STYLING|HBC|-80.992182|1.413580244274486|88|1
35.103409|e9115bec3c0b4905ddb152de25aab95e26806d52|3.5|2015-02-13 19:37:00|1.4132775322775095|3|20496000000|88|0.6126700657242101|0|58|755|-80.992182|87|35.103409|NFS-BALLOONS|0.0|9|*BALLOONS|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00204960000005|FLORAL|FLORAL|-80.992182|1.413580244274486|88|1
35.103409|7d3ef2d81ce26ec75a3e3cc39a6184b55ca6e742|2.39|2015-01-04 12:06:00|1.4132775322775095|3|5210004680|88|0.6126700657242101|0|58|734|-80.992182|3|35.103409|NFS-CANDLES/BIRTHDAY SUP|0.0|1|MC DECORATING TIPS|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00052100046808|BAKING SUPPLIES|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|e52c7779f92b3c6f4c0323c58779fd1c4e889bd9|6.98|2014-11-26 20:00:00|1.4132775322775095|3|7017706776|88|0.6126700657242101|0|58|230|-80.992182|37|35.103409|HERBAL TEA|1.98|1|TWININGS TEA HERB CHAMOMILE|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00070177067762|TEA|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|8cfab0f243db06126464dd52b3cb49c1e3f02bb5|3.39|2014-11-03 20:11:00|1.4132775322775095|3|5000012734|88|0.6126700657242101|0|58|341|-80.992182|57|35.103409|CREAMERS|0.0|3|COFFEEMATE FF HAZELNUT|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00050000127344|MILK|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|b72f13c5c26f901600202a241545b58041130c57|3.39|2014-11-22 19:08:00|1.4132775322775095|3|5000012734|88|0.6126700657242101|0|58|341|-80.992182|57|35.103409|CREAMERS|0.89|3|COFFEEMATE FF HAZELNUT|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00050000127344|MILK|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|65860b2be3a838d4fc3ad873508335aba960809c|3.39|2015-01-18 12:24:00|1.4132775322775095|3|5000012734|88|0.6126700657242101|0|58|341|-80.992182|57|35.103409|CREAMERS|0.89|3|COFFEEMATE FF HAZELNUT|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00050000127344|MILK|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|8f31b5680b433e6b34172e547b204974d4b92525|3.39|2014-12-29 19:03:00|1.4132775322775095|3|5000012734|88|0.6126700657242101|0|58|341|-80.992182|57|35.103409|CREAMERS|0.89|3|COFFEEMATE FF HAZELNUT|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00050000127344|MILK|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|764e472673103c47cd1c406ad347e8366ebd4c58|6.7|2015-02-19 18:49:00|1.4132775322775095|3|5000012734|88|0.6126700657242101|0|58|341|-80.992182|57|35.103409|CREAMERS|0.0|3|COFFEEMATE FF HAZELNUT|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00050000127344|MILK|DAIRY|-80.992182|1.413580244274486|88|2
35.103409|5924667a39e53badc7864f8104b99d21695170c3|3.39|2014-12-07 18:41:00|1.4132775322775095|3|5000012734|88|0.6126700657242101|0|58|341|-80.992182|57|35.103409|CREAMERS|0.0|3|COFFEEMATE FF HAZELNUT|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00050000127344|MILK|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|ef99df1812c94db3d64cb2e7199c6819f8be00a6|3.35|2015-02-15 18:34:00|1.4132775322775095|3|5000012734|88|0.6126700657242101|0|58|341|-80.992182|57|35.103409|CREAMERS|0.0|3|COFFEEMATE FF HAZELNUT|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00050000127344|MILK|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|901c391b86429f3687a3aad8a7242fd094d992d7|10.49|2014-12-03 23:41:00|1.4132775322775095|3|79849310320|88|0.6126700657242101|0|58|36|-80.992182|10|35.103409|PREMIUM GROUND|3.5|1|CARIBOU BLEND  GROUND COFFEE|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00798493103659|COFFEE|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|def7392617139aadaa3a56f3fe09d285551b7e30|2.29|2014-11-27 13:04:00|1.4132775322775095|3|5210004620|88|0.6126700657242101|0|58|18|-80.992182|3|35.103409|CAKE DECORATIONS & ICING|0.79|1|MC GREEN GEL|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00052100046303|BAKING SUPPLIES|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|e9a8d5c658607e003f246ec02aba252fa78ec3a4|9.29|2014-09-27 18:39:00|1.4132775322775095|3|7192101639|88|0.6126700657242101|0|58|284|-80.992182|892|35.103409|SUPER PREMIUM PIZZA|0.0|5|DIGIORNO 12in S/ C  PEPPERONI|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00071921016395|FROZEN PIZZA|FROZEN|-80.992182|1.413580244274486|88|1
35.103409|5264d0c1a85cf7a4855116e426db2c4f92181b81|4.99|2014-11-10 19:28:00|1.4132775322775095|3|7790019206|88|0.6126700657242101|0|58|487|-80.992182|105|35.103409|PRECOOKED B/FAST SAUSAGE|1.65|19|JIMMY DEAN TURKEY CRUMBLES|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00077900196317|BREAKFAST SAUSAGE|CASE READY MEATS|-80.992182|1.413580244274486|88|1
35.103409|0d7af25720b9d271ba5aa3aaeca2c1ed98138c2a|5.49|2015-01-03 19:43:00|1.4132775322775095|3|7447100078|88|0.6126700657242101|0|58|66|-80.992182|10|35.103409|GROUND CAN|0.0|1|MEDAGLIA D'ORO CAFFE' ESPRESSO|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00074471000784|COFFEE|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|64cc661751d6f2813c6675aad1214e282ddde2ed|1.63|2015-01-08 18:47:00|1.4132775322775095|3||88|0.6126700657242101|0|58|561|-80.992182|64|35.103409|FR PROD ORGANIC PRODUCE|0.0|4|COO ORG YUKON GOLD POTATOES|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00294727000003|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|1
35.103409|65f407af2c9b499c20e06503058f763e6057b06f|13.99|2015-01-25 18:18:00|1.4132775322775095|3|2124212009|88|0.6126700657242101|0|58|458|-80.992182|82|35.103409|CRAFT BEER|0.0|16|REDHOOK SAMPLER 12PK|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00021242120097|DOMESTIC BEER|BEER|-80.992182|1.413580244274486|88|1
35.103409|8b650e26fbae6dec5c71a7d7595da920b049365a|12.99|2015-02-22 19:01:00|1.4132775322775095|3|2124212009|88|0.6126700657242101|0|58|458|-80.992182|82|35.103409|CRAFT BEER|0.0|16|REDHOOK SAMPLER 12PK|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00021242120097|DOMESTIC BEER|BEER|-80.992182|1.413580244274486|88|1
35.103409|7d65de7006fff311c135a84e83d98784ed0519e2|13.99|2015-01-23 20:28:00|1.4132775322775095|3|2124212009|88|0.6126700657242101|0|58|458|-80.992182|82|35.103409|CRAFT BEER|0.0|16|REDHOOK SAMPLER 12PK|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00021242120097|DOMESTIC BEER|BEER|-80.992182|1.413580244274486|88|1
35.103409|49e11f202e0bdfd51ff709bb7bb9ed570569604f|25.98|2014-12-31 18:42:00|1.4132775322775095|3|2124212009|88|0.6126700657242101|0|58|458|-80.992182|82|35.103409|CRAFT BEER|0.0|16|REDHOOK SAMPLER 12PK|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00021242120097|DOMESTIC BEER|BEER|-80.992182|1.413580244274486|88|2
35.103409|005585bca4409333284da6ef21b516eb5ae9375f|12.99|2014-12-27 20:12:00|1.4132775322775095|3|2124212009|88|0.6126700657242101|0|58|458|-80.992182|82|35.103409|CRAFT BEER|0.0|16|REDHOOK SAMPLER 12PK|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00021242120097|DOMESTIC BEER|BEER|-80.992182|1.413580244274486|88|1
35.103409|16aac4894b4dd063ea66c374c23b9f9473052327|3.15|2014-09-22 19:04:00|1.4132775322775095|3|4127102564|88|0.6126700657242101|0|58|341|-80.992182|57|35.103409|CREAMERS|0.0|3|ITNAT'L HAZELNUT|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00041271025682|MILK|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|33e783b0304e38fddf4fd0d51c3a5f295f415a9d|7.99|2014-10-29 19:00:00|1.4132775322775095|3|71280812982|88|0.6126700657242101|0|58|458|-80.992182|82|35.103409|CRAFT BEER|0.0|16|HIGHLAND GAELIC ALE 6PK|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00712808129820|DOMESTIC BEER|BEER|-80.992182|1.413580244274486|88|1
35.103409|34b0cb54591eef139c5c30169ef0c7d4d64da1dd|3.89|2014-09-23 19:14:00|1.4132775322775095|3|3800039125|88|0.6126700657242101|0|58|74|-80.992182|9|35.103409|RTE CEREAL ALL FAMILY|0.9|1|KELLOGG RICE KRISPIES 9|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00038000318443|CEREAL|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|42f18068b2a5119850cbf6a20c8f74f03c858884|3.0|2014-11-25 21:58:00|1.4132775322775095|3|5000039758|88|0.6126700657242101|0|58|1147|-80.992182|229|35.103409|HOT COCOA MIX|1.0|1|NESTLE HOT COCOA RCH CHOCOLATE|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00050000397587|COCOAS CREAMERS SYRUPS|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|d46f6ee42650aa09709157d2cc03ab48f4919ca1|5.69|2014-10-02 19:15:00|1.4132775322775095|3|1101776290|88|0.6126700657242101|0|58|4895|-80.992182|1240|35.103409|FOOT ODOR/WETNESS|0.0|17|ODOR DESTROYERS DEOD SPRAY|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00011017762904|FOOT CARE|HBC|-80.992182|1.413580244274486|88|1
35.103409|7af27c9be2b388658e3c148b4ec11fdcae45302e|2.79|2015-01-16 06:38:00|1.4132775322775095|3|1600015110|88|0.6126700657242101|0|58|205|-80.992182|31|35.103409|REMAINING SNACKS|0.0|1|CHEX SNACK MIX - CHEDDAR|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00016000158405|SNACKS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|c4a4232a797e72f38cdd8edb2463855227c61a8e|11.99|2015-01-09 21:28:00|1.4132775322775095|3|8869286023|88|0.6126700657242101|0|58|9948|-80.992182|886|35.103409|NFS-PREM-CAB SAUVIGNON|0.0|13|STERLING VINTERS CAB SAUV|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00088692860232|PREMIUM ($8-$10.99)|WINE|-80.992182|1.413580244274486|88|1
35.103409|9ea686bb084809f7ec293fcc8e097bb6bcb612de|6.74|2014-10-21 19:01:00|1.4132775322775095|3|20319700000|88|0.6126700657242101|0|58|641|-80.992182|137|35.103409|PREMIUM PORK|1.2|2|VALUE PK PORK BUTT CNTRY RIB|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00203197000000|PORK|MEAT|-80.992182|1.413580244274486|88|1
35.103409|0870dae4dc54fabc1d4adb6f1b07265534364f48|1.01|2014-12-09 19:45:00|1.4132775322775095|3||88|0.6126700657242101|0|58|524|-80.992182|64|35.103409|FRESH PROD FRESH ONIONS|0.12|4|COO HONEY SWEET ONIONS|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00204166000007|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|1
35.103409|18894497084c5972b78de4579c5d992384e3dc56|5.55|2014-09-23 17:23:00|1.4132775322775095|3|20899600000|88|0.6126700657242101|0|58|1419|-80.992182|201|35.103409|SMART CHICKEN ORGANIC|0.0|2|SMART ORGANIC CHICKEN WINGS|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00208996000008|POULTRY|MEAT|-80.992182|1.413580244274486|88|1
35.103409|fae5c9695d349a89bac6744083c8ad593bc074b4|1.19|2014-10-04 22:14:00|1.4132775322775095|3|2146659306|88|0.6126700657242101|0|58|1730|-80.992182|392|35.103409|CANDLES|0.0|14|NUMBER 6 CANDLE|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00021466593066|DECORATING|BAKERY|-80.992182|1.413580244274486|88|1
35.103409|441e9e270c280b2572667839c0f71d839e6edc93|1.78|2014-10-27 19:44:00|1.4132775322775095|3||88|0.6126700657242101|0|58|561|-80.992182|64|35.103409|FR PROD ORGANIC PRODUCE|0.26|4|ORG TOMATOES|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00294799000000|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|1
35.103409|cf76e1b4954f690e929c46ea5edf88794e906f7f|0.5|2015-01-26 17:39:00|1.4132775322775095|3||88|0.6126700657242101|0|58|509|-80.992182|64|35.103409|FRESH CITRUS-REMAINING|0.0|4|COO LIMES, LRG|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00204048000002|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|1
35.103409|f76a76a0d86d5e6415a51669d58d4efae056e23d|17.99|2014-11-23 20:56:00|1.4132775322775095|3|7289000152|88|0.6126700657242101|0|58|459|-80.992182|83|35.103409|IMPORT BEER|0.0|16|HEINEKEN 18PK BTLS|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00072890001528|IMPORT BEER|BEER|-80.992182|1.413580244274486|88|1
35.103409|6271e872a063a715015701699e46c6ed1e556fe1|20.99|2014-09-14 20:36:00|1.4132775322775095|3|7289000152|88|0.6126700657242101|0|58|459|-80.992182|83|35.103409|IMPORT BEER|0.0|16|HEINEKEN 18PK BTLS|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00072890001528|IMPORT BEER|BEER|-80.992182|1.413580244274486|88|1
35.103409|d38089740f81da88cb22188082dc7f895ac23a4d|20.99|2014-09-21 20:39:00|1.4132775322775095|3|7289000152|88|0.6126700657242101|0|58|459|-80.992182|83|35.103409|IMPORT BEER|0.0|16|HEINEKEN 18PK BTLS|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00072890001528|IMPORT BEER|BEER|-80.992182|1.413580244274486|88|1
35.103409|2205034c9ce9e5ec2f788a7a0a912817ed33b4cd|17.99|2014-11-16 20:56:00|1.4132775322775095|3|7289000152|88|0.6126700657242101|0|58|459|-80.992182|83|35.103409|IMPORT BEER|0.0|16|HEINEKEN 18PK BTLS|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00072890001528|IMPORT BEER|BEER|-80.992182|1.413580244274486|88|1
35.103409|c22ff17155af3acac40555d11657ebc1fb798c08|17.99|2014-11-21 20:18:00|1.4132775322775095|3|7289000152|88|0.6126700657242101|0|58|459|-80.992182|83|35.103409|IMPORT BEER|0.0|16|HEINEKEN 18PK BTLS|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00072890001528|IMPORT BEER|BEER|-80.992182|1.413580244274486|88|1
35.103409|7518796e5361869d435ec68b0fb9259e3262a8bf|12.99|2014-10-23 21:38:00|1.4132775322775095|3|7289000016|88|0.6126700657242101|0|58|459|-80.992182|83|35.103409|IMPORT BEER|0.0|16|HEINEKEN 12PK 12OZ BOTTLES|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00072890000163|IMPORT BEER|BEER|-80.992182|1.413580244274486|88|1
35.103409|3c8c8b71797aba4b7450f5d99eb4a5ef18195ff7|12.99|2014-09-25 20:58:00|1.4132775322775095|3|7289000016|88|0.6126700657242101|0|58|459|-80.992182|83|35.103409|IMPORT BEER|0.0|16|HEINEKEN 12PK 12OZ BOTTLES|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00072890000163|IMPORT BEER|BEER|-80.992182|1.413580244274486|88|1
35.103409|fb109c79b60c33d84930a76a8e2791aba5148afe|24.99|2015-02-13 19:34:00|1.4132775322775095|3|7203696866|88|0.6126700657242101|0|58|740|-80.992182|87|35.103409|NFS-ROSE BQT|5.0|9|15 STEM ROSE BOUQUET|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00072036968661|FLORAL|FLORAL|-80.992182|1.413580244274486|88|1
35.103409|6b43f2d1530f722f0055372e08fec8579c45733f|12.99|2014-12-05 16:59:00|1.4132775322775095|3|8769201103|88|0.6126700657242101|0|58|458|-80.992182|82|35.103409|CRAFT BEER|0.0|16|SAM ADAMS SEASONAL 12PK|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00087692011033|DOMESTIC BEER|BEER|-80.992182|1.413580244274486|88|1
35.103409|f39af4d3b70534755dc1b8c0d3aa3171fc86b4c5|12.99|2014-12-06 22:26:00|1.4132775322775095|3|8769201103|88|0.6126700657242101|0|58|458|-80.992182|82|35.103409|CRAFT BEER|0.0|16|SAM ADAMS SEASONAL 12PK|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00087692011033|DOMESTIC BEER|BEER|-80.992182|1.413580244274486|88|1
35.103409|14c2855f86d3924f0506739b499547121da0dc62|4.95|2014-10-23 23:44:00|1.4132775322775095|3||88|0.6126700657242101|0|58|507|-80.992182|64|35.103409|FRESH ORANGES|0.19|4|NAVEL ORANGE, FL XL|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00204385000000|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|5
35.103409|0ab767f5ec0ee35627b18f2c99837da3c9af9ec5|7.65|2015-01-05 16:43:00|1.4132775322775095|3|76211120604|88|0.6126700657242101|0|58|36|-80.992182|10|35.103409|PREMIUM GROUND|0.0|1|STARBUCKS ESPRESSO ROAST COFFE|9f937055dc5c535198e99d38d3df13f059d7f21a|1.6769912711007346|0.61177642288969325|00762111206039|COFFEE|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.024464|1535d1f5a0d5aa45b6b33f65bb40ff730864cf3d|6.98|2014-09-26 11:27:00|80.848351720559364|2|3700022205|317|35.07123342569227|0|25|725|-80.848528|66|35.053394|NFS-DISHWASHING LIQUID|0.98|1|DAWN LIQ DISH ANTIBAC APPLE BL|a311a6dd70f5cdc114c30718fa3e271280055e47|3.2316545129474337|35.082633588753836|00037000222026|DETERGENTS|G1 GROCERY|-80.847383|80.847399919491735|11|2
35.024464|44040c6ec452f9de81bfd5e9093d881911f1a4ef|2.85|2014-12-21 18:31:00|80.848351720559364|2|4400000055|317|35.07123342538214|0|25|88|-80.8062|13|35.037115|FLAKED SODA CRACKERS|0.35|1|NABISCO PREMIUMS|a311a6dd70f5cdc114c30718fa3e271280055e47|3.2316545129474337|35.082633588753836|00044000000578|CRACKERS|G1 GROCERY|-80.847383|80.847401153554344|27|1
35.024464|24b9c8216f9e62918c700123fa64a860805c3ce5|7.35|2015-01-09 16:04:00|80.848351720559364|2|4470002268|317|35.071233421678031|0|25|358|-80.816172|100|35.059823|REGULAR BACON|3.68|19|OSCAR MAYER SLICED BACON|a311a6dd70f5cdc114c30718fa3e271280055e47|3.2316545129474337|35.082633588753836|00044700019887|BACON|CASE READY MEATS|-80.847383|80.847412094841218|66|1
35.024464|f795aef978a6bc82ee0606f390c8dad1d4004b6e|6.99|2014-09-30 19:17:00|1.41290891556208|2|4667716953|317|0.6112922155462233|0|33|6123|-80.847383|1546|35.024464|BULB-3 WAYS|0.0|18|PHILIPS 50/150W L/L 3WAY 3PK|a311a6dd70f5cdc114c30718fa3e271280055e47|3.2316545129474337|0.61055446569467375|00046677169534|LIGHT BULBS/ELECTRICAL|GM|-80.847383|1.4110530249708906|317|1
35.024464|ad56eba8003a32e7028528064ba01b11d7535417|3.69|2014-09-25 18:34:00|80.848351720559364|2|5783616826|317|35.07123342538214|0|25|532|-80.8062|64|35.037115|FRESH CUCUMBERS|0.0|4|MINI SEEDLESS CUCUMBERS|a311a6dd70f5cdc114c30718fa3e271280055e47|3.2316545129474337|35.082633588753836|00069905861062|FRESH PRODUCE|PRODUCE|-80.847383|80.847401153554344|27|1
35.024464|581208179b80dc1422b232bfbbffd321212b1a72|1.99|2014-09-18 20:19:00|80.848351720559364|2||317|35.07123342569227|0|25|535|-80.848528|64|35.053394|FRESH GREENS|0.0|4|SPINACH, BUNCH (RPC)|a311a6dd70f5cdc114c30718fa3e271280055e47|3.2316545129474337|35.082633588753836|00204090000005|FRESH PRODUCE|PRODUCE|-80.847383|80.847399919491735|11|1
35.024464|00d605c63b0573b8ff92a5d412433526888c0703|2.75|2015-02-08 18:16:00|80.848351720559364|2|2066200020|317|35.07123342538214|0|25|1219|-80.8062|275|35.037115|PASTA SC CORE|0.0|1|NEWMANS SC RST TOM GARLIC|a311a6dd70f5cdc114c30718fa3e271280055e47|3.2316545129474337|35.082633588753836|00020662004611|PASTA SAUCES|G1 GROCERY|-80.847383|80.847401153554344|27|1
35.024464|98ca4811de02a6a8e189877ca6ae64a10e527297|1.69|2014-09-12 13:43:00|80.848351720559364|2|7203688040|317|35.07123342538214|0|25|561|-80.8062|64|35.037115|FR PROD ORGANIC PRODUCE|0.19|4|ORG HT BABY CARROTS 1LB BAG|a311a6dd70f5cdc114c30718fa3e271280055e47|3.2316545129474337|35.082633588753836|00072036880406|FRESH PRODUCE|PRODUCE|-80.847383|80.847401153554344|27|1
35.024464|ccae1545be360d37b9514eb6048dff9e90ebecb5|8.99|2014-10-11 15:47:00|80.848351720559364|2|2301290142|317|35.07123342538214|0|25|1477|-80.8062|485|35.037115|SUSHI HYBRID|0.0|6|CRUNCHY DRAGON ROLL SP|a311a6dd70f5cdc114c30718fa3e271280055e47|3.2316545129474337|35.082633588753836|00023012901424|SUSHI|DELI|-80.847383|80.847401153554344|27|1
35.024464|4d776c1195240083a45d14cd429127bb069843f2|9.99|2014-09-17 10:12:00|80.848351720559364|2|8500001868|317|35.071233421678031|0|25|9944|-80.816172|885|35.059823|NFS POP OTHER RED|0.0|13|BAREFOOT SWEET RED 1.5L|a311a6dd70f5cdc114c30718fa3e271280055e47|3.2316545129474337|35.082633588753836|00085000018682|POPULAR (4-$7.99)|WINE|-80.847383|80.847412094841218|66|1
35.024464|255c555591b8dd14062c4630690977b673f1c9c9|3.69|2014-09-20 17:57:00|80.848351720559364|2|20892500000|317|35.07123342538214|0|25|658|-80.8062|137|35.037115|FRESH PORK SAUSAGE|0.0|2|PORK ITALIAN SWEET SAUSAGE|a311a6dd70f5cdc114c30718fa3e271280055e47|3.2316545129474337|35.082633588753836|00208925000000|PORK|MEAT|-80.847383|80.847401153554344|27|1
35.024464|62844e829c2fff73d063265ab49183ed86dd7aaa|4.99|2014-09-30 10:51:00|80.848351720559364|2|70708210032|317|35.07123342538214|0|25|232|-80.8062|37|35.037115|WELLNESS TEA|0.0|1|OREGON CHAI ORG TEA ORIG LIQ|a311a6dd70f5cdc114c30718fa3e271280055e47|3.2316545129474337|35.082633588753836|00707082100320|TEA|G1 GROCERY|-80.847383|80.847401153554344|27|1
35.024464|db0ac43c36abcb273d99ee1632243db6b936833f|0.68|2014-10-24 19:01:00|80.848351720559364|2||317|35.071233421678031|0|25|534|-80.816172|64|35.059823|FRESH CHILI PEPPERS|0.0|4|COO ORANGE HABANERO CHILI|a311a6dd70f5cdc114c30718fa3e271280055e47|3.2316545129474337|35.082633588753836|00204711000001|FRESH PRODUCE|PRODUCE|-80.847383|80.847412094841218|66|1
35.024464|3ef46d04ab0ba6024032a671fb973057215a634e|0.84|2014-09-11 19:44:00|80.848351720559364|2||317|35.07123342538214|0|25|534|-80.8062|64|35.037115|FRESH CHILI PEPPERS|0.0|4|COO ORANGE HABANERO CHILI|a311a6dd70f5cdc114c30718fa3e271280055e47|3.2316545129474337|35.082633588753836|00204711000001|FRESH PRODUCE|PRODUCE|-80.847383|80.847401153554344|27|1
35.024464|fc82908f077e2a08b38d0083e24f1088d55e92e4|0.6|2014-09-13 18:48:00|80.848351720559364|2||317|35.07123342538214|0|25|530|-80.8062|64|35.037115|FRESH CABBAGE|0.0|4|COO GREEN CABBAGE|a311a6dd70f5cdc114c30718fa3e271280055e47|3.2316545129474337|35.082633588753836|00204069000005|FRESH PRODUCE|PRODUCE|-80.847383|80.847401153554344|27|1
35.024464|dc2f244667c7200d80be1538ea26c693d43e8321|11.99|2015-01-31 14:41:00|80.848351720559364|2|82471033315|317|35.07123342569227|0|25|663|-80.848528|154|35.053394|FISH FILLETS/STEAKS PKGD|3.02|12|PIER 33 VP SALMON PORTION|a311a6dd70f5cdc114c30718fa3e271280055e47|3.2316545129474337|35.082633588753836|00824710333155|FISH FILLETS/STEAKS|SEAFOOD|-80.847383|80.847399919491735|11|1
35.066546|b6cafdc6e0a84d6c6b113e7850b4a9887ee26cea|4.99|2014-10-24 17:35:00|1.4091206135396188|4|71575620002|45|0.6120266850020475|0|47|504|-80.771677|64|35.066546|FRESH BERRIES|2.5|4|STRAWBERRIES 1LB CLAM|a51527394aa27f93b542347e6fb696426cf7ee2e|0.5958199724277814|0.61242566243833529|00715756200023|FRESH PRODUCE|PRODUCE|-80.771677|1.409731706007376|45|1
35.066546|5e8682f4fda87e4f1f63e97d19f2dd8317a77ce7|3.89|2015-02-05 19:26:00|1.4091206135396188|4|5210007139|45|0.6120266850020475|0|47|1246|-80.771677|34|35.066546|SPICE BLENDS|0.0|1|MC GARLIC POWDER CALIFORNIA|a51527394aa27f93b542347e6fb696426cf7ee2e|0.5958199724277814|0.61242566243833529|00052100071398|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.771677|1.409731706007376|45|1
35.066546|94bab397fd2e35c4f54e95292366592ca5483163|2.99|2014-10-07 16:48:00|80.782094729586973|4|2066200020|45|35.075168873237558|0|27|1219|-80.739|275|35.141204|PASTA SC CORE|0.7|1|NEWMANS SC TOM BASIL BOMBOLINA|a51527394aa27f93b542347e6fb696426cf7ee2e|0.5958199724277814|35.102887530186244|00020662000286|PASTA SAUCES|G1 GROCERY|-80.771677|80.771686751411735|171|1
35.066546|fc101bebbaa639c6d1733710120904069ff469c9|5.6|2014-10-03 08:48:00|80.782094729586973|4|20563700000|45|35.075168876008178|0|27|1823|-80.8062|410|35.037115|BH HAM|0.0|6|BOARS HEAD SWEET SLICE HAM|a51527394aa27f93b542347e6fb696426cf7ee2e|0.5958199724277814|35.102887530186244|00205637000007|BH MEAT|DELI|-80.771677|80.771681874226886|27|1
35.066546|463c0b80d394d0a44aecf324c945b9a802e74f53|9.49|2014-10-22 08:51:00|80.782094729586973|4|20598400000|45|35.075168876008178|0|27|1822|-80.8062|410|35.037115|BH CHICKEN|0.0|6|BOARS HEAD EVERROAST CKN BRST|a51527394aa27f93b542347e6fb696426cf7ee2e|0.5958199724277814|35.102887530186244|00205984000002|BH MEAT|DELI|-80.771677|80.771681874226886|27|1
35.066546|63db6e3a15ba413c7b86f768ade074e00a899bb6|9.99|2014-10-02 19:10:00|1.4091206135396188|4|7203695262|45|0.6120266850020475|0|47|1671|-80.771677|383|35.066546|CHEESE CAKE|1.0|14|FRESH MADE MARBLE CHEESCAKE|a51527394aa27f93b542347e6fb696426cf7ee2e|0.5958199724277814|0.61242566243833529|00072036950758|PASTRY CASE|BAKERY|-80.771677|1.409731706007376|45|1
35.123768|58b869d94cf201b5fdcd14b392899867a4c2bff1|2.89|2015-03-08 11:18:00|80.6036218474908|2|2100065894|473|35.242502025096968|0|34|1441|-80.62331|274|35.140781|MAC AND CHEESE|0.0|1|KRAFT DIN MAC CHS FAMILY|a7e5886834041f364131cb2d24f4d9fcee198054|8.204234815178278|35.262263711360632|00021000658947|PREP FOODS DINNERS|G1 GROCERY|-80.654118|80.654164116708827|39|1
35.123768|7cee7e304143d5a237fc6046e130c4751193bb5f|7.99|2015-01-03 09:46:00|80.6036218474908|2|2100061161|473|35.242502025096968|0|34|314|-80.62331|52|35.140781|CHEESE-PROCESSED-OTHER|0.0|3|KRAFT VELVEETA CHEESE|a7e5886834041f364131cb2d24f4d9fcee198054|8.204234815178278|35.262263711360632|00021000611614|CHEESE|DAIRY|-80.654118|80.654164116708827|39|1
35.123768|54ca5c61c9024e324959e384bc1358718512f6a7|2.19|2015-01-17 08:23:00|80.6036218474908|2|7418226090|473|35.242501995622476|0|34|722|-80.64817|73|35.04711|NFS-HAND SOAPS|1.19|1|SS HAND SOAP PUMP COCONUT GING|a7e5886834041f364131cb2d24f4d9fcee198054|8.204234815178278|35.262263711360632|00074182270919|PERSONAL SOAP/BATH ADDITIVES|G1 GROCERY|-80.654118|80.65423027034474|129|1
35.123768|025fd5476411f366e44da8b681ae715b87500784|0.55|2015-01-25 13:41:00|80.6036218474908|2||473|35.242502025096968|0|34|522|-80.62331|64|35.140781|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|a7e5886834041f364131cb2d24f4d9fcee198054|8.204234815178278|35.262263711360632|00204664000004|FRESH PRODUCE|PRODUCE|-80.654118|80.654164116708827|39|1
35.123768|03e3c0539ac7c38c6d92b1f787aa5ae4939f9795|1.69|2014-12-10 12:23:00|80.6036218474908|2|4900000044|473|35.242502025096968|0|34|55|-80.62331|8|35.140781|REGULAR|0.0|23|CB COKE SINGLE 20 OZ.|a7e5886834041f364131cb2d24f4d9fcee198054|8.204234815178278|35.262263711360632|00049000000443|CARBONATED BEVERAGES|BEVERAGE|-80.654118|80.654164116708827|39|1
35.123768|36127ac8bac02ee56f77d506f0a520b5de78d8bd|2.79|2015-01-05 18:30:00|80.6036218474908|2|7225001130|473|35.242502025096968|0|34|1033|-80.62331|163|35.140781|HAMBURGER|0.0|7|MERITA 8PK HAMBURGER BUNS|a7e5886834041f364131cb2d24f4d9fcee198054|8.204234815178278|35.262263711360632|00072250011303|BUNS/ROLLS|COMMERCIAL BAKERY|-80.654118|80.654164116708827|39|1
35.123768|4366eeca888a9dce58278afd2c930d857325ba6c|4.59|2015-01-04 06:43:00|80.6036218474908|2|1340945132|473|35.242501995622476|0|34|68|-80.64817|11|35.04711|BARBECUE SAUCES|0.0|1|SWEET BABY RAY 40 BBQ BRW SUGR|a7e5886834041f364131cb2d24f4d9fcee198054|8.204234815178278|35.262263711360632|00013409515372|CONDIMENTS|G1 GROCERY|-80.654118|80.65423027034474|129|1
35.123768|d58cb76605282188be8f3560bf69df8603b31208|1.39|2015-02-07 18:31:00|80.6036218474908|2|2200000488|473|35.242501955318176|0|34|48|-80.771677|7|35.066546|REGISTER GUM|0.0|1|(FE)ORBIT SPEARMINT GUM 14 PC|a7e5886834041f364131cb2d24f4d9fcee198054|8.204234815178278|35.262263711360632|00022000004840|CANDY|G1 GROCERY|-80.654118|80.654282110916768|45|1
35.123768|6744f4a215a0dc5379786620fd55686ab0db3c71|1.9|2014-12-29 09:37:00|80.6036218474908|2|61300871771|473|35.242501995622476|0|34|99|-80.64817|32|35.04711|LIQUID TEA|0.15|1|GOLDEN BEAR LEMONADE|a7e5886834041f364131cb2d24f4d9fcee198054|8.204234815178278|35.262263711360632|00613008734862|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.654118|80.65423027034474|129|2
35.123768|f5b8eea1c079dacfe9088bb77d15e222713f54e7|34.99|2015-01-15 14:18:00|80.6036218474908|2|87126000460|473|35.242502027701576|0|34|740|-80.709466|87|35.124987|NFS-ROSE BQT|15.0|9|DZ COLOR ROSE BQT    ELITE|a7e5886834041f364131cb2d24f4d9fcee198054|8.204234815178278|35.262263711360632|00871260004608|FLORAL|FLORAL|-80.654118|80.654152653161049|157|1
35.384824|7c0c77060b067fb0577777e44526a813fbb98a0f|3.29|2015-02-27 17:58:00|80.779636304526477|4|7203695076|476|35.410690199773462|0|17|1609|-80.782849|371|35.372142|TAKE & BAKE BREAD|0.0|14|TAKE & BAKE SMALL WHEAT FRENCH|a92fb6c7128277df7eefa7b7c6fb6d7df1dc798a|1.787291953670539|35.392509581117899|00072036950765|BREAD|BAKERY|-80.784334|80.784337966121981|122|1
35.384824|7ba022e31f8051ffaa8dfda94d71ae956e60c8d8|1.25|2014-09-22 20:05:00|80.779636304526477|4|2550020188|476|35.410690199773462|0|17|67|-80.782849|10|35.372142|SOLUBLE INSTANT|0.25|1|FOLGER INST CRYST SNGL SRV REG|a92fb6c7128277df7eefa7b7c6fb6d7df1dc798a|1.787291953670539|35.392509581117899|00025500201887|COFFEE|G1 GROCERY|-80.784334|80.784337966121981|122|1
35.384824|121b2f426d5b08125e4bb1dc702a1367669251ff|1.95|2014-10-25 19:04:00|80.779636304526477|4|5480003077|476|35.410690199773462|0|17|138|-80.782849|38|35.372142|RICE MICROWAVE|0.0|1|UNCLE BEN RR RED BEANS N RICE.|a92fb6c7128277df7eefa7b7c6fb6d7df1dc798a|1.787291953670539|35.392509581117899|00054800420056|RICE GRAINS AND BEANS|G1 GROCERY|-80.784334|80.784337966121981|122|1
35.384824|bc6d2c0c696fb8e7581262b0c9ce1156ddbc5dff|6.99|2015-02-16 16:02:00|1.4102725052409182|4|7203602601|476|0.61758168403871|0|1|1981|-80.784334|480|35.384824|CHIPS|2.0|6|HTT 18OZ MULTI GRAIN PITA CHIP|a92fb6c7128277df7eefa7b7c6fb6d7df1dc798a|1.787291953670539|0.61833652052202714|00072036026040|DRY GOODS|DELI|-80.784334|1.4099526123308008|476|1
35.384824|9135828e7050a9e0356561d912fc5b03bd865e1d|4.88|2014-12-07 13:47:00|80.779636304526477|4||476|35.410690199773462|0|17|501|-80.782849|64|35.372142|FRESH PEARS|0.0|4|BOSC PEARS|a92fb6c7128277df7eefa7b7c6fb6d7df1dc798a|1.787291953670539|35.392509581117899|00204413000002|FRESH PRODUCE|PRODUCE|-80.784334|80.784337966121981|122|1
35.384824|d814fe52bf5a97d1924ead6aee28183aa741414e|4.49|2014-11-03 19:12:00|80.779636304526477|4|7203676180|476|35.410690199773462|0|17|122|-80.782849|19|35.372142|HONEY|0.0|1|HT TRADER EUCALYPTUS HONEY|a92fb6c7128277df7eefa7b7c6fb6d7df1dc798a|1.787291953670539|35.392509581117899|00072036982759|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.784334|80.784337966121981|122|1
35.384824|2442d9db385a80c8de746d822c52fa23fd1c89c4|5.99|2014-09-10 19:50:00|80.779636304526477|4|2550081121|476|35.410690199773462|0|17|37|-80.782849|10|35.372142|PODS/CUPS/SINGLES|0.0|1|FOLGERS SINGLES REGULAR 19 BAG|a92fb6c7128277df7eefa7b7c6fb6d7df1dc798a|1.787291953670539|35.392509581117899|00025500811215|COFFEE|G1 GROCERY|-80.784334|80.784337966121981|122|1
35.384824|7e4c89325951db4faf8ef0dcf3e3926a0f5c0420|1.89|2014-12-09 16:04:00|80.779636304526477|4|7203695050|476|35.410690156457811|0|17|1605|-80.810056|371|35.219587|PAR BAKED (BREAD)|0.0|14|SMALL HONEY WHEAT FRENCH|a92fb6c7128277df7eefa7b7c6fb6d7df1dc798a|1.787291953670539|35.392509581117899|00072036950505|BREAD|BAKERY|-80.784334|80.784392207145885|401|1
35.006282|6c6de6a0afdca0f8e2bffc055b5c7a45938ca56e|1.04|2015-03-01 11:34:00|80.562862110758871|4||60|35.07927644082752|0|21|522|-80.760919|64|35.024332|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|b15bee016b63ffedcec519af3d65454b98ce4d6b|5.043740853804177|35.054042368968126|00204664000004|FRESH PRODUCE|PRODUCE|-80.562829|80.562892216644201|343|1
35.006282|4e8940a612b0e9b1fd96118866eff9268599821d|4.19|2015-01-18 12:56:00|80.562862110758871|4|2900007325|60|35.07927644082752|0|21|1149|-80.760919|21|35.024332|PEANUTS|1.19|1|PLANTERS D/R PEANUTS|b15bee016b63ffedcec519af3d65454b98ce4d6b|5.043740853804177|35.054042368968126|00029000073258|NUTS|G1 GROCERY|-80.562829|80.562892216644201|343|1
35.006282|23fc752f84880cad5222ee72bfa69090e0eee61c|9.98|2014-12-24 18:24:00|1.4091206135396188|4|7203688079|60|0.6109748797816256|0|47|523|-80.562829|64|35.006282|FRESH POTATOES|0.0|4|HT WHITE POTATO 5LB BAG|b15bee016b63ffedcec519af3d65454b98ce4d6b|5.043740853804177|0.61242566243833529|00072036880796|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|2
35.006282|f927f99304dce02e23377616145ea6fb9f352fc0|1.89|2014-10-15 15:21:00|80.562862110758871|4|31254662380|60|35.079276385136232|0|21|4207|-80.758228|1200|34.95459|COUGH DROP-ADULT|0.0|17|HALLS STRAWBERRY     -62380|b15bee016b63ffedcec519af3d65454b98ce4d6b|5.043740853804177|35.054042368968126|00312546623804|COUGH/COLD/SINUS|HBC|-80.562829|80.562955986428719|182|1
35.603432|129b3222dc5ee24e8809bc5e1bf43489050a1389|13.99|2014-11-26 17:04:00|1.4102725052409182|3|8066095615|274|0.6213971134099097|0|1|459|-80.895009|83|35.603432|IMPORT BEER|0.0|16|CORONA EXTRA 12PK 12OZ BTL|b2d96d6d4691710b170baf365e42ee5579b41978|2.7571517018135867|0.61833652052202714|00080660956152|IMPORT BEER|BEER|-80.895009|1.4118842554804456|274|1
35.603432|794380a51169167e3ff0ef0463d16639d16990d0|1.95|2014-12-07 12:20:00|1.4102725052409182|3|930000011|274|0.6213971134099097|0|1|161|-80.895009|25|35.603432|PEPPERS|0.0|1|MT OLV BANANA PEPPER MILD FP|b2d96d6d4691710b170baf365e42ee5579b41978|2.7571517018135867|0.61833652052202714|00009300001021|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.895009|1.4118842554804456|274|1
35.603432|d7da80b30bf1e71358848444b448839e936ef82a|11.58|2014-12-26 17:35:00|1.4102725052409182|3|4400000665|274|0.6213971134099097|0|1|1254|-80.895009|12|35.603432|FUDGE ENROBED|2.6|1|NABISCO MALLOMARS|b2d96d6d4691710b170baf365e42ee5579b41978|2.7571517018135867|0.61833652052202714|00044000006747|COOKIES|G1 GROCERY|-80.895009|1.4118842554804456|274|2
35.603432|22f9bc45e45aaf8845be53ad11d213680bdf7cae|3.69|2014-12-24 14:07:00|1.4102725052409182|3|71514172928|274|0.6213971134099097|0|1|330|-80.895009|55|35.603432|EGGS|0.0|3|EGGLAND BEST GRADE A EX-LG EGG|b2d96d6d4691710b170baf365e42ee5579b41978|2.7571517018135867|0.61833652052202714|00715141729283|EGGS FRESH|DAIRY|-80.895009|1.4118842554804456|274|1
35.603432|075972359cd9291dc4b8d916bde5562d36b5edc5|2.29|2015-03-08 13:18:00|1.4102725052409182|3|7203663996|274|0.6213971134099097|0|1|342|-80.895009|57|35.603432|FRESH MILK|0.0|3|HARRIS TEETER WHOLE MILK|b2d96d6d4691710b170baf365e42ee5579b41978|2.7571517018135867|0.61833652052202714|00072036639967|MILK|DAIRY|-80.895009|1.4118842554804456|274|1
35.603432|51a3db6338a4a5e9c576c16cf4bfa06cbbc6e753|6.57|2015-03-06 22:39:00|1.4102725052409182|3|1200000496|274|0.6213971134099097|0|1|54|-80.895009|8|35.603432|DIET|0.52|23|DIET PEPSI 2 LTR NR|b2d96d6d4691710b170baf365e42ee5579b41978|2.7571517018135867|0.61833652052202714|00012000002311|CARBONATED BEVERAGES|BEVERAGE|-80.895009|1.4118842554804456|274|3
35.603432|cabe0da21cd1d40ad884661dc8ae9514156bdf09|23.98|2014-11-30 14:35:00|1.4102725052409182|3|3125900923|274|0.6213971134099097|0|1|9936|-80.895009|885|35.603432|NFS POP MERLOT|0.0|13|YELLOW TAIL MERLOT 1.5L|b2d96d6d4691710b170baf365e42ee5579b41978|2.7571517018135867|0.61833652052202714|00031259009230|POPULAR (4-$7.99)|WINE|-80.895009|1.4118842554804456|274|2
35.341927|49212c5b7fedbad2a3fc9cee3c1abf71e8c2f60e|1.29|2014-09-25 13:14:00|80.779636304526477|4|8379152001|220|35.388384739568522|0|17|1981|-80.780702|480|35.318911|CHIPS|0.18|6|DIRTY POTATO CHIP BBQ|b4ac9585d5997003eaa1b9e6290fb6ec1349617b|3.2101177698257164|35.392509581117899|00083791520049|DRY GOODS|DELI|-80.764523|80.764540821253263|167|1
35.341927|bbb882b0bb8e6a4d10488ff48954d2f4ee22688c|7.99|2015-02-08 12:58:00|1.4102725052409182|4|1820012989|220|0.6168329901494819|0|1|457|-80.764523|82|35.341927|DOMESTIC SINGLES/SIX PACKS|0.0|16|MICHELOB ULTRA LIME CACTUS 6PK|b4ac9585d5997003eaa1b9e6290fb6ec1349617b|3.2101177698257164|0.61833652052202714|00018200129896|DOMESTIC BEER|BEER|-80.764523|1.4096068451526882|220|1
35.341927|50d09383e58fa64547de50a09598ac54f32fee5c|9.38|2014-10-01 17:19:00|1.4102725052409182|4|74236526435|220|0.6168329901494819|0|1|345|-80.764523|57|35.341927|ORGANIC MILK|0.0|3|HORIZON WHOLE  DHA|b4ac9585d5997003eaa1b9e6290fb6ec1349617b|3.2101177698257164|0.61833652052202714|00742365264474|MILK|DAIRY|-80.764523|1.4096068451526882|220|2
35.341927|96333a6b73efa33d8f36bf9b8ce3e0e2e04fb335|5.19|2015-02-10 18:09:00|80.779636304526477|4|74236526435|220|35.388384739086376|0|17|345|-80.737839|57|35.297134|ORGANIC MILK|0.0|3|HORIZON WHOLE  DHA|b4ac9585d5997003eaa1b9e6290fb6ec1349617b|3.2101177698257164|35.392509581117899|00742365264474|MILK|DAIRY|-80.764523|80.764542620517034|258|1
35.341927|247e7e51a071516e5e6e3e935a0aafcbb9a189c1|9.78|2014-11-09 12:37:00|80.779636304526477|4|74236526435|220|35.388384739086376|1|17|345|-80.737839|57|35.297134|ORGANIC MILK|0.0|3|HORIZON WHOLE  DHA|b4ac9585d5997003eaa1b9e6290fb6ec1349617b|3.2101177698257164|35.392509581117899|00742365264474|MILK|DAIRY|-80.764523|80.764542620517034|258|2
35.341927|5d5a3924be5bb1f43832f0f91523a28a815632de|17.99|2014-10-02 17:22:00|1.4102725052409182|4|1820096292|220|0.6168329901494819|0|1|456|-80.764523|82|35.341927|DOMESTIC SUPER PREM 12PK&>|0.0|16|BUD LIGHT LIME 18PK BOTTLES|b4ac9585d5997003eaa1b9e6290fb6ec1349617b|3.2101177698257164|0.61833652052202714|00018200962929|DOMESTIC BEER|BEER|-80.764523|1.4096068451526882|220|1
35.341927|cecd802d84f5121ef4529aed98661bd3d5404dec|17.99|2014-10-03 18:34:00|1.4102725052409182|4|1820096292|220|0.6168329901494819|0|1|456|-80.764523|82|35.341927|DOMESTIC SUPER PREM 12PK&>|0.0|16|BUD LIGHT LIME 18PK BOTTLES|b4ac9585d5997003eaa1b9e6290fb6ec1349617b|3.2101177698257164|0.61833652052202714|00018200962929|DOMESTIC BEER|BEER|-80.764523|1.4096068451526882|220|1
35.341927|4df3d669926eecc29da99c5ad68b6849962238f8|13.38|2015-01-14 10:53:00|1.4102725052409182|4|20298800000|220|0.6168329901494819|0|1|652|-80.764523|141|35.341927|FRESH LAMB PRIMALS|0.0|2|LAMB LOIN CHOP|b4ac9585d5997003eaa1b9e6290fb6ec1349617b|3.2101177698257164|0.61833652052202714|00202988000007|LAMB|MEAT|-80.764523|1.4096068451526882|220|1
35.341927|fd447756e0273a708994de7c5e41974a14be2b6b|8.97|2015-02-01 13:38:00|80.779636304526477|4|7203671072|220|35.388384739086376|0|17|317|-80.737839|52|35.297134|CHUNK AND BAR CHEESE|0.0|3|HT EXTRA SHARP CHEDDAR CHEESE|b4ac9585d5997003eaa1b9e6290fb6ec1349617b|3.2101177698257164|35.392509581117899|00072036710734|CHEESE|DAIRY|-80.764523|80.764542620517034|258|1
35.23102|b8ffde7c625d71f2d286ae8f7b71c0c411b36a25|1.7|2014-11-20 22:03:00|80.843945456961976|4|7203636026|205|35.233525626650305|0|59|55|-80.80146|8|35.17739|REGULAR|0.35|23|HT CLUB SODA|b98d7ebe997751130de4e0245b89435f1e7ca0a4|0.17313276225630675|35.232478750868765|00072036360274|CARBONATED BEVERAGES|BEVERAGE|-80.8438|80.843801122560265|208|2
35.23102|7d065f2b6eb21f32909842fd0fea1a0c4e2d01df|1.7|2014-12-08 15:48:00|80.843945456961976|4|7203636026|205|35.233525626150509|0|59|55|-80.825175|8|35.152722|REGULAR|0.7|23|HT CLUB SODA|b98d7ebe997751130de4e0245b89435f1e7ca0a4|0.17313276225630675|35.232478750868765|00072036360274|CARBONATED BEVERAGES|BEVERAGE|-80.8438|80.843802239207946|160|2
35.23102|739073c3705ff6ae430f9cbbbabc8d00261959bb|2.59|2014-09-22 20:44:00|80.843945456961976|4|7047041381|205|35.233525626650305|0|59|687|-80.80146|61|35.17739|BLENDED|0.0|3|YOPLAIT HARVEST PEACH 4PK|b98d7ebe997751130de4e0245b89435f1e7ca0a4|0.17313276225630675|35.232478750868765|00070470434834|YOGURT|DAIRY|-80.8438|80.843801122560265|208|1
35.23102|108c1b706df3ab1d4421ac283fbbf859b1f85aee|5.39|2015-02-16 19:47:00|80.843945456961976|4|74759961699|205|35.233525626650305|0|59|1147|-80.80146|229|35.17739|HOT COCOA MIX|0.0|1|GHIRADELLI DOUBLE CHOC COCOA|b98d7ebe997751130de4e0245b89435f1e7ca0a4|0.17313276225630675|35.232478750868765|00747599616990|COCOAS CREAMERS SYRUPS|G1 GROCERY|-80.8438|80.843801122560265|208|1
35.23102|bc8b0874f5d0ea27e8a07b3cd47ce1fd75db1963|2.79|2015-02-15 18:46:00|80.843945456961976|4|7225001131|205|35.233525626150509|0|59|1034|-80.825175|163|35.152722|HOT DOG|0.0|7|MERITA 8PK HOTDOG BUN|b98d7ebe997751130de4e0245b89435f1e7ca0a4|0.17313276225630675|35.232478750868765|00072250011310|BUNS/ROLLS|COMMERCIAL BAKERY|-80.8438|80.843802239207946|160|1
35.23102|20249307209c1bbb1bc503c890b532738d6fd212|1.97|2014-12-07 19:09:00|80.843945456961976|4|7203631016|205|35.233525626119864|0|59|1245|-80.849471|34|35.161696|SINGLE SPICES|0.0|1|E  HT CINNAMON|b98d7ebe997751130de4e0245b89435f1e7ca0a4|0.17313276225630675|35.232478750868765|00072036310163|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.8438|80.84380229003186|35|1
35.23102|b89e219f616495c408ff59c8c57a3e93f97582dd|5.33|2014-12-22 22:15:00|80.843945456961976|4|20337700000|205|35.233525626816629|0|59|641|-80.810056|137|35.219587|PREMIUM PORK|0.0|2|PORK LOIN CHOPS BNLS THIN|b98d7ebe997751130de4e0245b89435f1e7ca0a4|0.17313276225630675|35.232478750868765|00203377000004|PORK|MEAT|-80.8438|80.843800104392102|401|1
35.23102|9bfe36f3851bcfd068458c8d14f8e52363aaf3a0|3.19|2014-12-21 13:56:00|80.843945456961976|4|74759961274|205|35.233525626119864|0|59|16|-80.849471|3|35.161696|BAKING CHOCOLATE/CHIPS/MORSELS|0.69|1|GHIRADELLI SEMI SWT CHOC CH|b98d7ebe997751130de4e0245b89435f1e7ca0a4|0.17313276225630675|35.232478750868765|00747599640155|BAKING SUPPLIES|G1 GROCERY|-80.8438|80.84380229003186|35|1
35.23102|cffdf4ef0118078e233cb730771e61d17e4bf710|3.49|2014-12-16 21:41:00|80.843945456961976|4|4400001473|205|35.233525626119864|0|59|1248|-80.849471|12|35.161696|SANDWICH COOKIES|0.49|1|WHITE FUDGE OREO|b98d7ebe997751130de4e0245b89435f1e7ca0a4|0.17313276225630675|35.232478750868765|00044000014735|COOKIES|G1 GROCERY|-80.8438|80.84380229003186|35|1
35.23102|ac4fd0bb08a2c62761cc715e7a550aea0e865096|0.29|2014-11-08 12:17:00|80.843945456961976|4||205|35.233525626150509|0|59|502|-80.825175|64|35.152722|FRESH BANANAS|0.0|4|BANANAS, YELLOW|b98d7ebe997751130de4e0245b89435f1e7ca0a4|0.17313276225630675|35.232478750868765|00204011000008|FRESH PRODUCE|PRODUCE|-80.8438|80.843802239207946|160|1
35.23102|a1bd089aace1f31c80dfdc67839345a6e895e31f|4.99|2015-01-25 13:24:00|80.843945456961976|4|8265750406|205|35.233525626650305|0|59|31|-80.80146|4|35.17739|NON CARBONATED WATER|1.49|1|(U)DEER PARK WATER 24PK .5LT|b98d7ebe997751130de4e0245b89435f1e7ca0a4|0.17313276225630675|35.232478750868765|00082657504063|BOTTLED WATER|G1 GROCERY|-80.8438|80.843801122560265|208|1
35.123768|e6524805da82410db32b47180904f32bbf9fbe06|3.49|2015-02-09 18:36:00|80.632521683083056|4|3010000133|473|35.180478696713905|0|39|88|-80.62331|13|35.140781|FLAKED SODA CRACKERS|0.99|1|ZESTA ORIGINAL|bcc27d42065e355e7ff3438266e55b6324731957|3.9185723887938253|35.177497916598789|00030100001331|CRACKERS|G1 GROCERY|-80.654118|80.654140009823365|39|1
35.123768|f8021a1a33bba0c661892b5039e35e9f9e211574|3.19|2015-02-25 19:35:00|80.632521683083056|4|7225001120|473|35.180478682646807|0|39|1026|-80.64817|162|35.04711|WHEAT|0.0|7|MERITA 100% WHEAT BREAD 20OZ|bcc27d42065e355e7ff3438266e55b6324731957|3.9185723887938253|35.177497916598789|00072250011204|SLICED BREAD|COMMERCIAL BAKERY|-80.654118|80.654171582541338|129|1
35.123768|07d35856521e021241899d5d2f9ae890a075a96e|4.49|2015-02-20 16:45:00|80.632521683083056|4|7336077201|473|35.180478696713905|0|39|30|-80.62331|4|35.140781|CARBONATED WATER|0.0|1|LACROIX CUR CHRY LIME 8PK|bcc27d42065e355e7ff3438266e55b6324731957|3.9185723887938253|35.177497916598789|00073360772023|BOTTLED WATER|G1 GROCERY|-80.654118|80.654140009823365|39|1
35.123768|0bc013802d50dbf2a10b551ddf80d99d7ac861d1|6.78|2015-01-07 18:32:00|80.632521683083056|4|7196000500|473|35.180478696713905|0|39|187|-80.62331|29|35.140781|SALMON-CANNED|0.39|1|ROYAL PINK SALMON 14.75 OZ|bcc27d42065e355e7ff3438266e55b6324731957|3.9185723887938253|35.177497916598789|00071960005008|SEAFOOD-CANNED|G1 GROCERY|-80.654118|80.654140009823365|39|2
35.123768|5cf0dcc1d0d3d695c61c248e8b9a9d6db55ea895|3.19|2014-11-26 19:33:00|80.632521683083056|4|7203655010|473|35.180478680891419|0|39|317|-80.562829|52|35.006282|CHUNK AND BAR CHEESE|0.0|3|HT EXTRA SHARP CHEDDAR CHEESE|bcc27d42065e355e7ff3438266e55b6324731957|3.9185723887938253|35.177497916598789|00072036559951|CHEESE|DAIRY|-80.654118|80.65417429309008|60|1
35.123768|9b24eb3f8126f60473cd4b4ee0a48607539eb208|4.99|2015-02-16 14:24:00|80.632521683083056|4|76235737516|473|35.180478696713905|0|39|577|-80.62331|136|35.140781|OTHER MERCH FR MSC JUICE|0.0|4|EVOLUTION COCONUT WATER GREENS|bcc27d42065e355e7ff3438266e55b6324731957|3.9185723887938253|35.177497916598789|00762357375162|OTHER MERCHANDISE|PRODUCE|-80.654118|80.654140009823365|39|1
35.123768|8be719a054addab2e29b03333de7c927452f1cfe|4.99|2014-10-27 18:45:00|80.632521683083056|4|7203688080|473|35.180478680891419|0|39|523|-80.562829|64|35.006282|FRESH POTATOES|2.5|4|HT YUKON GOLD 5 LB BAG|bcc27d42065e355e7ff3438266e55b6324731957|3.9185723887938253|35.177497916598789|00072036880802|FRESH PRODUCE|PRODUCE|-80.654118|80.65417429309008|60|1
35.123768|138a5f8e2c29256264daf47ba657203f73985fb9|4.99|2015-02-18 15:57:00|80.632521683083056|4|7203688080|473|35.180478696713905|0|39|523|-80.62331|64|35.140781|FRESH POTATOES|0.0|4|HT YUKON GOLD 5 LB BAG|bcc27d42065e355e7ff3438266e55b6324731957|3.9185723887938253|35.177497916598789|00072036880802|FRESH PRODUCE|PRODUCE|-80.654118|80.654140009823365|39|1
35.123768|1ee824f24d20643bef6f223fc5be4f71945a1acb|2.78|2014-12-28 19:50:00|80.632521683083056|4|5210094269|473|35.180478696713905|0|39|80|-80.62331|34|35.140781|SEASONING PACKETS|0.78|1|MC WHITE CHICKEN CHILI SEAS|bcc27d42065e355e7ff3438266e55b6324731957|3.9185723887938253|35.177497916598789|00052100007809|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.654118|80.654140009823365|39|2
35.123768|241540be9c5cf2f1e555a061b5a40480c7ef6ef9|2.0|2015-02-06 17:37:00|80.632521683083056|4|4000000435|473|35.180478680891419|0|39|47|-80.562829|7|35.006282|REGISTER BARS|0.0|1|(FE)M&M PEANUT CANDY|bcc27d42065e355e7ff3438266e55b6324731957|3.9185723887938253|35.177497916598789|00040000000327|CANDY|G1 GROCERY|-80.654118|80.65417429309008|60|2
35.123768|0f50e561b90e2eaf3275582811d3b39286f3ddb9|3.39|2014-12-15 16:39:00|80.632521683083056|4||473|35.180478696713905|0|39|500|-80.62331|64|35.140781|FRESH APPLES|0.0|4|RED DEL APPLE, WA  48|bcc27d42065e355e7ff3438266e55b6324731957|3.9185723887938253|35.177497916598789|00233284000002|FRESH PRODUCE|PRODUCE|-80.654118|80.654140009823365|39|1
35.123768|75a5bc99b9585e50a88308f3412cee661ea9496f|19.99|2015-02-14 09:05:00|80.632521683083056|4|20496500000|473|35.180478682646807|0|39|751|-80.64817|87|35.04711|NFS-BOUQUETS|0.0|9|*BOUQUETS|bcc27d42065e355e7ff3438266e55b6324731957|3.9185723887938253|35.177497916598789|00204965000000|FLORAL|FLORAL|-80.654118|80.654171582541338|129|1
35.123768|3ff24bbf3a801cb5533bfb0cf4569c3b4712cb4d|19.98|2014-12-13 08:52:00|80.632521683083056|4|7203696996|473|35.180478682646807|0|39|751|-80.64817|87|35.04711|NFS-BOUQUETS|0.0|9|9.99 DUOCHROMATIC BQT  SS|bcc27d42065e355e7ff3438266e55b6324731957|3.9185723887938253|35.177497916598789|00072036969965|FLORAL|FLORAL|-80.654118|80.654171582541338|129|2
35.585842|3bf27b9279fee911929affaf569dc37aa33c46a0|3.79|2015-02-01 15:48:00|1.4102725052409182|4|4950800600|99|0.6210901099944839|0|1|1981|-80.875654|480|35.585842|CHIPS|1.8|6|SALT & PEPPER PRETZEL CRISPS|bd5b046a04a6e26c8fae21d6cbf74ab665225c11|2.7742842793455997|0.61833652052202714|00049508100034|DRY GOODS|DELI|-80.875654|1.411546447003722|99|1
35.585842|fa211845eec1063a02375e3f19ffcb0b4f88045e|5.1|2015-02-06 21:10:00|1.4102725052409182|4|4369505631|99|0.6210901099944839|0|1|1276|-80.875654|279|35.585842|FROZEN SANDWICHES|2.12|5|LEAN POCKETS 3 CHSE & BROCCOLI|bd5b046a04a6e26c8fae21d6cbf74ab665225c11|2.7742842793455997|0.61833652052202714|00043695083187|FROZEN SANDWICH AND SNACKS|FROZEN|-80.875654|1.411546447003722|99|2
35.585842|7a75228bb97550b6c94153ae3d2a066e2c926a74|3.99|2015-02-17 13:47:00|1.4102725052409182|4|7203670859|99|0.6210901099944839|0|1|1280|-80.875654|48|35.585842|MULTI SERVE MEALS|0.99|5|HTT CHICKEN FRIED RICE|bd5b046a04a6e26c8fae21d6cbf74ab665225c11|2.7742842793455997|0.61833652052202714|00072036708618|FROZEN MEALS|FROZEN|-80.875654|1.411546447003722|99|1
35.585842|d3bd53c8329da6bc8138f280dfe8d21e8753977e|9.98|2014-11-01 16:07:00|1.4102725052409182|4|2410044068|99|0.6210901099944839|0|1|87|-80.875654|13|35.585842|CHEESE CRACKERS|2.99|1|CHEEZ-IT HOT AND SPICY|bd5b046a04a6e26c8fae21d6cbf74ab665225c11|2.7742842793455997|0.61833652052202714|00024100789092|CRACKERS|G1 GROCERY|-80.875654|1.411546447003722|99|2
35.585842|060f062552d3ae958953d9238cd7a59646177e31|3.29|2015-01-28 17:08:00|80.891462859624312|4|2840004768|99|35.625992185896969|0|45|202|-80.8955|31|35.4437|PRETZELS|0.79|1|ROLD GOLD PRETZEL THINS|bd5b046a04a6e26c8fae21d6cbf74ab665225c11|2.7742842793455997|35.636605227883024|00028400231879|SNACKS|G1 GROCERY|-80.875654|80.875731234810701|272|1
35.585842|0062e4ad37d00b25abf017df02448b4a8fa6398c|2.29|2014-10-04 19:47:00|80.891462859624312|4|7203695175|99|35.625992234825418|0|45|1607|-80.895009|371|35.603432|FROZEN DOUGH (BREAD)|0.0|14|FRESH LRG FRENCH BREAD|bd5b046a04a6e26c8fae21d6cbf74ab665225c11|2.7742842793455997|35.636605227883024|00072036951755|BREAD|BAKERY|-80.875654|80.875658641592082|274|1
35.585842|b1e5c6c73600e10f9cafaed9dbf668d36b87415e|2.15|2014-10-08 19:04:00|1.4102725052409182|4|3800030110|99|0.6210901099944839|0|1|44|-80.875654|6|35.585842|TOASTER PASTRIES-SHELF STABLE|0.0|1|KELL POPTART CONFETTI CUPCAKE|bd5b046a04a6e26c8fae21d6cbf74ab665225c11|2.7742842793455997|0.61833652052202714|00038000713422|BREAKFAST FOODS|G1 GROCERY|-80.875654|1.411546447003722|99|1
35.585842|b95c9a91fdaf597eb7c6a0f8f2347e8c9977802a|1.99|2014-10-15 09:55:00|80.891462859624312|4||99|35.625992234825418|0|45|540|-80.895009|64|35.603432|FRESH CELERY|0.3|4|COO CELERY (RPC) 24'S|bd5b046a04a6e26c8fae21d6cbf74ab665225c11|2.7742842793455997|35.636605227883024|00204070000001|FRESH PRODUCE|PRODUCE|-80.875654|80.875658641592082|274|1
35.585842|082f52d2f1dab8c9b1e5c14c9a9ce4569422e739|4.99|2014-11-26 16:51:00|80.891462859624312|4|7790019206|99|35.625992234825418|0|45|487|-80.895009|105|35.603432|PRECOOKED B/FAST SAUSAGE|0.0|19|JIMMY DEAN TURKEY CRUMBLES|bd5b046a04a6e26c8fae21d6cbf74ab665225c11|2.7742842793455997|35.636605227883024|00077900196317|BREAKFAST SAUSAGE|CASE READY MEATS|-80.875654|80.875658641592082|274|1
35.585842|2a55997938b5525326e37fefa15e862bcfe0a257|3.89|2014-10-13 09:42:00|80.891462859624312|4|7535511201|99|35.625992234825418|0|45|128|-80.895009|20|35.603432|APPLE JUICE-SHELF|0.4|1|OLD ORHRD ORGANIC APL JUICE|bd5b046a04a6e26c8fae21d6cbf74ab665225c11|2.7742842793455997|35.636605227883024|00075355112012|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.875654|80.875658641592082|274|1
35.585842|fe714653927c22f5f890221fe43892ea9ee822e9|1.99|2015-02-09 15:46:00|1.4102725052409182|4|7205860615|99|0.6210901099944839|0|1|1211|-80.875654|272|35.585842|HISP SALSA/DIPS|0.74|1|MRS WAGES MIX GUACAMOLE|bd5b046a04a6e26c8fae21d6cbf74ab665225c11|2.7742842793455997|0.61833652052202714|00072058606152|HISPANIC PREP. FOODS|G1 GROCERY|-80.875654|1.411546447003722|99|1
35.585842|3c51047ef0c02b0b86c14721f1b2bbe0683f32c3|3.99|2014-10-15 09:57:00|80.891462859624312|4|7430500116|99|35.625992234825418|0|45|82|-80.895009|11|35.603432|VINEGAR|0.0|1|BRAGG ORG VINEGAR APPLE CIDER|bd5b046a04a6e26c8fae21d6cbf74ab665225c11|2.7742842793455997|35.636605227883024|00074305001161|CONDIMENTS|G1 GROCERY|-80.875654|80.875658641592082|274|1
35.585842|e0b0a4b8776823fe8091339def87c5c8263d3f1b|3.99|2014-12-18 09:20:00|80.891462859624312|4|7430500116|99|35.625992234825418|0|45|82|-80.895009|11|35.603432|VINEGAR|0.0|1|BRAGG ORG VINEGAR APPLE CIDER|bd5b046a04a6e26c8fae21d6cbf74ab665225c11|2.7742842793455997|35.636605227883024|00074305001161|CONDIMENTS|G1 GROCERY|-80.875654|80.875658641592082|274|1
35.585842|790c953e9143d17d684f2950ddb1c7420aa7cd9d|5.99|2015-02-11 16:18:00|1.4102725052409182|4|7756725423|99|0.6210901099944839|0|1|252|-80.875654|45|35.585842|PREMIUM ICE CREAM|2.99|5|BREYERS CHOCOLATE I/C|bd5b046a04a6e26c8fae21d6cbf74ab665225c11|2.7742842793455997|0.61833652052202714|00077567254207|ICE CREAM|FROZEN|-80.875654|1.411546447003722|99|1
35.585842|d72a6cdd4ec1d512616a29c0568964db92153e2c|3.34|2014-11-18 19:58:00|1.4102725052409182|4|7203643010|99|0.6210901099944839|0|1|252|-80.875654|45|35.585842|PREMIUM ICE CREAM|0.0|5|HT PREM COOKIES & CREAM IC|bd5b046a04a6e26c8fae21d6cbf74ab665225c11|2.7742842793455997|0.61833652052202714|00072036430229|ICE CREAM|FROZEN|-80.875654|1.411546447003722|99|1
35.585842|05a1076f29748315f0e8f6f1aa40bf5d245e2643|3.34|2015-01-29 21:23:00|1.4102725052409182|4|7203643010|99|0.6210901099944839|0|1|252|-80.875654|45|35.585842|PREMIUM ICE CREAM|0.84|5|HT PREM MOOSE TRACKS IC|bd5b046a04a6e26c8fae21d6cbf74ab665225c11|2.7742842793455997|0.61833652052202714|00072036430328|ICE CREAM|FROZEN|-80.875654|1.411546447003722|99|1
35.585842|23c0c440e207d36e40dcbb9016176821d041b2b3|3.33|2015-03-06 21:27:00|1.4102725052409182|4|7203643010|99|0.6210901099944839|0|1|252|-80.875654|45|35.585842|PREMIUM ICE CREAM|0.0|5|HT PREM MOOSE TRACKS IC|bd5b046a04a6e26c8fae21d6cbf74ab665225c11|2.7742842793455997|0.61833652052202714|00072036430328|ICE CREAM|FROZEN|-80.875654|1.411546447003722|99|1
35.585842|9fd64a0b560acf359a7d0ecf146b01403d4eb9f9|6.99|2014-10-18 19:45:00|1.4102725052409182|4|7192196239|99|0.6210901099944839|0|1|284|-80.875654|892|35.585842|SUPER PREMIUM PIZZA|1.99|5|DIGIORNO ITALIAN CHICKEN PARM|bd5b046a04a6e26c8fae21d6cbf74ab665225c11|2.7742842793455997|0.61833652052202714|00071921843830|FROZEN PIZZA|FROZEN|-80.875654|1.411546447003722|99|1
35.585842|27b10e41842fd9668bc1adc39606620367af3a89|6.99|2015-01-08 10:02:00|80.891462859624312|4|3700088942|99|35.625992234825418|0|45|4092|-80.895009|1080|35.603432|TOOTHPASTE-WHITENING|2.0|17|CREST 3DW BRILLIANCE TOOTHPAST|bd5b046a04a6e26c8fae21d6cbf74ab665225c11|2.7742842793455997|35.636605227883024|00037000889427|ORAL HYGIENE|HBC|-80.875654|80.875658641592082|274|1
35.585842|98e71ebbe1b28b7c3c51722c3672af6035ee73e7|3.49|2014-11-15 13:29:00|1.4102725052409182|4|7797508161|99|0.6210901099944839|0|1|204|-80.875654|31|35.585842|TORTILLA CHIPS|0.99|1|SOH RESTURNT STYLE TORTILLA CH|bd5b046a04a6e26c8fae21d6cbf74ab665225c11|2.7742842793455997|0.61833652052202714|00077975081785|SNACKS|G1 GROCERY|-80.875654|1.411546447003722|99|1
35.585842|6c21629cd421e32fb69a328d64afac21c69eda5d|1.27|2014-09-15 18:49:00|1.4102725052409182|4|5963500189|99|0.6210901099944839|0|1|1461|-80.875654|40|35.585842|FROZEN GARLIC TOAST AND BRD|0.0|5|FURLANI TEXAS TOAST|bd5b046a04a6e26c8fae21d6cbf74ab665225c11|2.7742842793455997|0.61833652052202714|00059635001890|FROZEN DOUGH|FROZEN|-80.875654|1.411546447003722|99|1
35.585842|e3b3f89481fd11f3f7dbd0a755e75ddd68a2e61d|3.35|2014-10-20 19:00:00|1.4102725052409182|4|7203656080|99|0.6210901099944839|0|1|318|-80.875654|52|35.585842|SHREDDED/GRATED CHEESE|0.0|3|HT SHRED SHARP CHED CHEESE 2%|bd5b046a04a6e26c8fae21d6cbf74ab665225c11|2.7742842793455997|0.61833652052202714|00072036590466|CHEESE|DAIRY|-80.875654|1.411546447003722|99|1
35.03469|95b22f07a8b1386946a05a30eee175051f01d50f|4.39|2014-12-17 17:23:00|80.970593795509558|2|4400002796|82|35.068500512103562|0|4|90|-80.837892|13|34.937113|SNACK CRACKERS|2.2|1|TRISCUIT ORIGINAL|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00044000027957|CRACKERS|G1 GROCERY|-80.97058|80.970597291516128|372|1
35.03469|78f91ab607d2d860498e20c3be72547d41fa5649|3.79|2014-12-19 07:28:00|80.970593795509558|2|4850002013|82|35.068500514562629|0|4|335|-80.994596|56|35.061685|ORANGE JUICE-REGRIGERATED|0.79|3|TROPICANA PP W/CALCIUM|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00048500305690|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.97058|80.970587132420093|475|1
35.03469|25fc9617d520409cd3f946db623f0fe0d01317ba|1.29|2014-10-18 16:44:00|80.970593795509558|2|85382600333|82|35.068500514562629|0|4|104|-80.994596|16|35.061685|APPLESAUCE-CUPS|0.0|1|D HAPPY SQZ ORG POM BLUE APPLE|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00853826003331|FRUIT-CAN/JAR|G1 GROCERY|-80.97058|80.970587132420093|475|1
35.03469|b21ea8fbc0c9ac0fe0beee3eb7bcd2d4d14dd214|1.59|2015-02-15 09:34:00|1.4132775322775095|2|85382600333|82|0.6114706929155321|0|58|104|-80.97058|16|35.03469|APPLESAUCE-CUPS|0.8|1|D HAPPY SQZ ORG POM BLUE APPLE|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|0.61177642288969325|00853826003331|FRUIT-CAN/JAR|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|62b1e0b45bd0b4c581868133c4e069782d8dd213|7.99|2015-01-04 19:06:00|1.4132775322775095|2|7560904128|82|0.6114706929155321|0|58|3249|-80.97058|1020|35.03469|FACIAL CLEANSER|2.0|17|OLAY REGEN CLEANSER|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|0.61177642288969325|00075609601477|FACIAL CLEANSER & MOISTURIZER|HBC|-80.97058|1.4132032182494703|82|1
35.03469|4cbe1e4e90979a6252106b048ade217491749310|3.39|2015-01-24 20:20:00|80.970593795509558|2|7460900007|82|35.068500514562629|0|4|71|-80.994596|11|35.061685|GROC CONDIMENTS MARINADE|0.0|1|D  KCM MARINADE CARIBBEAN JERK|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00074609054399|CONDIMENTS|G1 GROCERY|-80.97058|80.970587132420093|475|1
35.03469|0a5e868a36a1a3d6483c34a75c1fcc5cde365c02|4.85|2014-10-24 17:41:00|1.4132775322775095|2|7790011553|82|0.6114706929155321|0|58|361|-80.97058|105|35.03469|BREAKFAST SAUSAGE|0.0|19|JIMMY DEAN MILD SAUSAGE|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|0.61177642288969325|00077900115530|BREAKFAST SAUSAGE|CASE READY MEATS|-80.97058|1.4132032182494703|82|1
35.03469|40b18ba8261be9743e952bfff1dcd8f6a35e4a50|7.99|2014-11-02 08:53:00|80.970593795509558|2|7560904128|82|35.068500514562629|0|4|3249|-80.994596|1020|35.061685|FACIAL CLEANSER|0.0|17|OLAY REGEN CLEANSER|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00075609601477|FACIAL CLEANSER & MOISTURIZER|HBC|-80.97058|80.970587132420093|475|1
35.03469|494cb21414da22543e454b7c686bc104710e8f21|1.59|2014-11-28 18:28:00|80.970593795509558|2|8190000008|82|35.068500514562629|0|4|1218|-80.994596|273|35.061685|ASIAN OTHER|0.0|1|KOALA COOKIE CHOCOLATE|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00081900000086|ASIAN PREP. FOODS|G1 GROCERY|-80.97058|80.970587132420093|475|1
35.03469|7b337f40a4cad71c4bb4797ed05ce87f9a906a06|3.89|2014-11-26 13:53:00|80.970593795509558|2|2100012277|82|35.068500514562629|0|4|320|-80.994596|53|35.061685|COTTAGE CHEESE|0.0|3|BREAKSTONE 2% COTTAGE CHEESE|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00021000123544|CULTURES|DAIRY|-80.97058|80.970587132420093|475|1
35.03469|59b918768b4f1dc4f8921b131d461dbfae098519|10.99|2014-11-30 12:22:00|80.970593795509558|2|3329300300|82|35.068500159096104|0|4|9983|-80.8955|889|35.4437|NFS-SPARKLING|0.0|13|FREIXENET CORDON NEGRO BRUT|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00033293003007|SPARKLING|WINE|-80.97058|80.970769520619641|272|1
35.03469|3b529cfa47ace592509510f03575601c5a681ca5|1.99|2015-03-03 18:53:00|80.970593795509558|2|3000016920|82|35.068500514562629|0|4|721|-80.994596|31|35.061685|RICE SNACKS|0.0|1|QUAKER RICE CRISP BUTR POPCRN|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00030000319772|SNACKS|G1 GROCERY|-80.97058|80.970587132420093|475|1
35.03469|11f60a95194da7b74e261ac6b6f2904d60b28724|6.99|2014-11-14 18:53:00|80.970593795509558|2|3913116852|82|35.068500514562629|0|4|254|-80.994596|892|35.061685|PREMIUM PIZZA|0.0|5|BELLATORIA ULTIMATE PEPPERONI|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00039131168525|FROZEN PIZZA|FROZEN|-80.97058|80.970587132420093|475|1
35.03469|e742b6a44a3b11101a3222c13d6a6c16e0eea6e5|6.99|2015-02-05 18:34:00|80.970593795509558|2|3913116852|82|35.068500514562629|0|4|254|-80.994596|892|35.061685|PREMIUM PIZZA|0.0|5|BELLATORIA ULTIMATE PEPPERONI|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00039131168525|FROZEN PIZZA|FROZEN|-80.97058|80.970587132420093|475|1
35.03469|da024cc3dc523181bd143e97e7660a729945bafc|1.59|2014-09-19 11:46:00|80.970593795509558|2|78616201000|82|35.068500508622286|0|4|31|-80.992182|4|35.103409|NON CARBONATED WATER|0.59|1|VIT WATER XXX 20 OZ|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00786162150004|BOTTLED WATER|G1 GROCERY|-80.97058|80.970605500300422|88|1
35.03469|2df3a4c7c82194ce4114caf0a7be32ab93dac341|9.99|2014-12-21 16:01:00|80.970593795509558|2|8500001443|82|35.068500514562629|0|4|9938|-80.994596|885|35.061685|NFS POP PINOT GRS/GRIGIO|0.0|13|CB-BAREFOOT PINOT GRIGIO 1.5L|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00085000014431|POPULAR (4-$7.99)|WINE|-80.97058|80.970587132420093|475|1
35.03469|1dcd246a936421fd0597356c503ed07ccec32adf|10.99|2014-11-16 12:37:00|80.970593795509558|2|8500001443|82|35.068500514562629|0|4|9938|-80.994596|885|35.061685|NFS POP PINOT GRS/GRIGIO|0.0|13|CB-BAREFOOT PINOT GRIGIO 1.5L|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00085000014431|POPULAR (4-$7.99)|WINE|-80.97058|80.970587132420093|475|1
35.03469|7971f952c9ad629a976d433e28c5a05d2b795a0d|10.99|2015-01-14 20:39:00|80.970593795509558|2|8500001443|82|35.068500514562629|0|4|9938|-80.994596|885|35.061685|NFS POP PINOT GRS/GRIGIO|0.0|13|CB-BAREFOOT PINOT GRIGIO 1.5L|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00085000014431|POPULAR (4-$7.99)|WINE|-80.97058|80.970587132420093|475|1
35.03469|635fdad3acabd123567cb9cf5be32df0b3abc863|9.99|2014-10-02 19:25:00|80.970593795509558|2|8500001443|82|35.068500514562629|0|4|9938|-80.994596|885|35.061685|NFS POP PINOT GRS/GRIGIO|0.0|13|CB-BAREFOOT PINOT GRIGIO 1.5L|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00085000014431|POPULAR (4-$7.99)|WINE|-80.97058|80.970587132420093|475|1
35.03469|0c762e24f1b50e77c06f49302e34f6a5d7358576|10.99|2014-10-12 17:58:00|80.970593795509558|2|8500001443|82|35.068500514562629|0|4|9938|-80.994596|885|35.061685|NFS POP PINOT GRS/GRIGIO|0.0|13|CB-BAREFOOT PINOT GRIGIO 1.5L|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00085000014431|POPULAR (4-$7.99)|WINE|-80.97058|80.970587132420093|475|1
35.03469|e7988b6192904afe3c526518828ea0b9119752b5|9.99|2014-10-07 17:29:00|1.4132775322775095|2|8500001443|82|0.6114706929155321|0|58|9938|-80.97058|885|35.03469|NFS POP PINOT GRS/GRIGIO|0.0|13|CB-BAREFOOT PINOT GRIGIO 1.5L|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|0.61177642288969325|00085000014431|POPULAR (4-$7.99)|WINE|-80.97058|1.4132032182494703|82|1
35.03469|cca30f4ea781de3c892b38de4b625db27b2dbcd6|9.99|2014-11-11 17:50:00|80.970593795509558|2|8500001443|82|35.068500514562629|0|4|9938|-80.994596|885|35.061685|NFS POP PINOT GRS/GRIGIO|0.0|13|CB-BAREFOOT PINOT GRIGIO 1.5L|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00085000014431|POPULAR (4-$7.99)|WINE|-80.97058|80.970587132420093|475|1
35.03469|b71a4974571c02bdefe46b2c66a94a84538f697d|9.99|2014-12-08 15:22:00|80.970593795509558|2|8500001443|82|35.068500514562629|0|4|9938|-80.994596|885|35.061685|NFS POP PINOT GRS/GRIGIO|0.0|13|CB-BAREFOOT PINOT GRIGIO 1.5L|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00085000014431|POPULAR (4-$7.99)|WINE|-80.97058|80.970587132420093|475|1
35.03469|5980327028a882ad05cc18b6fd552c68f4b554ac|3.58|2014-10-17 20:25:00|80.970593795509558|2|4850001775|82|35.068500514562629|0|4|335|-80.994596|56|35.061685|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA 50 W/CALCIUM 12 OZ|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00048500019047|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.97058|80.970587132420093|475|2
35.03469|415682e7e8dffaea8935a2b1ba002c0a50cd4a1d|2.5|2014-09-17 17:45:00|1.4132775322775095|2|81851201703|82|0.6114706929155321|0|58|43|-80.97058|6|35.03469|INSTANT BREAKFAST-POWDERED|0.51|1|SPROUT RSE STWBRY BAN SMOOTHIE|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|0.61177642288969325|00818512017016|BREAKFAST FOODS|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|0d43919605bc3fb1484b34cef6aabf566b968df5|8.99|2014-11-09 08:01:00|80.970593795509558|2|8380407471|82|35.068500514562629|0|4|9983|-80.994596|889|35.061685|NFS-SPARKLING|0.0|13|COOKS STOWAWAYS BRUT 4PK|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00083804074712|SPARKLING|WINE|-80.97058|80.970587132420093|475|1
35.03469|c0de0b09d69ce80cb568d1b3c829c5706389e6fd|8.99|2015-01-09 17:34:00|80.970593795509558|2|8380407471|82|35.068500514562629|0|4|9983|-80.994596|889|35.061685|NFS-SPARKLING|0.0|13|COOKS STOWAWAYS BRUT 4PK|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00083804074712|SPARKLING|WINE|-80.97058|80.970587132420093|475|1
35.03469|7db13019378821741315254aa16be1bb1a9f550a|8.99|2014-12-30 17:40:00|1.4132775322775095|2|8380407471|82|0.6114706929155321|0|58|9983|-80.97058|889|35.03469|NFS-SPARKLING|0.0|13|COOKS STOWAWAYS BRUT 4PK|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|0.61177642288969325|00083804074712|SPARKLING|WINE|-80.97058|1.4132032182494703|82|1
35.03469|e965b2c61b3eff3a6659a95f481ea6c9a7d3155d|8.99|2015-03-01 18:35:00|1.4132775322775095|2|8380407471|82|0.6114706929155321|0|58|9983|-80.97058|889|35.03469|NFS-SPARKLING|0.0|13|COOKS STOWAWAYS BRUT 4PK|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|0.61177642288969325|00083804074712|SPARKLING|WINE|-80.97058|1.4132032182494703|82|1
35.03469|7039c8df5f1434fac92d6fdaee979feeb6cec0bd|5.99|2014-09-20 11:43:00|80.970593795509558|2|73127991266|82|35.068500514562629|0|4|184|-80.994596|28|35.061685|SALAD DRESSINGS-LIQUID|0.0|1|T LISH DRS VIN CHIPOTLE|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00731279912663|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.97058|80.970587132420093|475|1
35.03469|a725cc5545887813d9115ec0b45a59bd4358da53|8.49|2014-12-18 18:19:00|80.970593795509558|2|2301290136|82|35.068500514562629|0|4|1477|-80.994596|485|35.061685|SUSHI HYBRID|0.0|6|CRUNCHY ROLL SP|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00023012901363|SUSHI|DELI|-80.97058|80.970587132420093|475|1
35.03469|49d3aa36f34144b5c72f6c3dbab46d8d2bd3566b|8.99|2014-09-27 17:10:00|80.970593795509558|2|1820017993|82|35.068500514562629|0|4|458|-80.994596|82|35.061685|CRAFT BEER|0.0|16|SHOCK TOP SEASONAL 6PK|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00018200179938|DOMESTIC BEER|BEER|-80.97058|80.970587132420093|475|1
35.03469|20e5868a2bc659fcfef40592ced54f3b0025dd65|10.99|2015-02-14 10:05:00|80.970593795509558|2|20499400000|82|35.068500514562629|0|4|755|-80.994596|87|35.061685|NFS-BALLOONS|2.0|9|"*AD - 36"" Jumbo Balloon"|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00204994000002|FLORAL|FLORAL|-80.97058|80.970587132420093|475|1
35.03469|79d24d5d9772efabcdc4604ccd41bc215ebe4736|3.65|2014-10-31 07:32:00|80.970593795509558|2|3010003012|82|35.068500514562629|0|4|91|-80.994596|13|35.061685|SPRAYED BUTTER CRACKERS|0.65|1|KEELBER CLUB ORIGINAL|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00030100100577|CRACKERS|G1 GROCERY|-80.97058|80.970587132420093|475|1
35.03469|037709c740416996b82317eb86f4784be92f43a0|2.79|2014-10-16 07:24:00|80.970593795509558|2|7203620074|82|35.068500514562629|0|4|128|-80.994596|20|35.061685|APPLE JUICE-SHELF|0.79|1|HT APPLE JUICE - PLST|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00072036200723|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.97058|80.970587132420093|475|1
35.03469|84695777ccf508f3c9b174d0d6e3821dad8d38ae|5.99|2014-12-27 20:15:00|80.970593795509558|2|82927451375|82|35.068500514562629|0|4|152|-80.994596|24|35.061685|NFS-CAT FOOD DRY|1.0|1|MEOW MIX HAIRBALL CONTROL FORM|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00851599000397|PET FOOD/SUPPLIES|G1 GROCERY|-80.97058|80.970587132420093|475|1
35.03469|518e784646d40b45ef7748a3b14270c625e790a5|1.49|2014-10-07 11:43:00|80.970593795509558|2|1200080008|82|35.068500508622286|0|4|55|-80.992182|8|35.103409|REGULAR|0.5|23|PEPSI 1.5L|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00012000800085|CARBONATED BEVERAGES|BEVERAGE|-80.97058|80.970605500300422|88|1
35.03469|094597a8bbb734a20a3e02f388e8e204bb802fe3|10.99|2014-11-24 17:39:00|1.4132775322775095|2|1834115102|82|0.6114706929155321|0|58|9937|-80.97058|885|35.03469|NFS POP SAUV/FUME BLANC|0.0|13|BAREFOOT SAUV BLANC 1.5L|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|0.61177642288969325|00018341151022|POPULAR (4-$7.99)|WINE|-80.97058|1.4132032182494703|82|1
35.03469|b6843cc2b14328c8b3cabf58b37ce7f7aa5ed8ee|9.99|2015-01-03 18:34:00|80.970593795509558|2|8769282102|82|35.068500514562629|0|4|463|-80.994596|84|35.061685|HARD CIDER|0.0|16|ANGRY ORCHARD CRISP APPLE 6PK|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00087692821021|SPECIALTY|BEER|-80.97058|80.970587132420093|475|1
35.03469|c5460479f06463854a1f3b2177230c377ca6e8e5|3.69|2014-10-21 19:24:00|80.970593795509558|2|7127926102|82|35.068500508622286|0|4|555|-80.992182|64|35.103409|PACKAGED SALADS|0.0|4|F.E. HEARTS OF ROMAINE|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00071279261027|FRESH PRODUCE|PRODUCE|-80.97058|80.970605500300422|88|1
35.03469|6d90b8656ee5116f9cb4b4da6508d014e312e255|19.99|2015-01-22 19:28:00|80.970593795509558|2|79500800100|82|35.068500514562629|0|4|8092|-80.994596|1705|35.061685|PROPANE EXCHANGE|0.0|18|BLUE RHINO CYLINDER EXCHANGE|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00795008001004|PROPANE|GM|-80.97058|80.970587132420093|475|1
35.03469|2e9630adfdc166949e4960b2c37eee8e96e40569|8.99|2015-02-14 15:44:00|1.4132775322775095|2|8380404721|82|0.6114706929155321|0|58|9983|-80.97058|889|35.03469|NFS-SPARKLING|0.0|13|CB-COOKS BRUT CHAMPAGNE|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|0.61177642288969325|00083804047211|SPARKLING|WINE|-80.97058|1.4132032182494703|82|1
35.03469|86e6232723bb9e291418d7c80708e3f30ed7a24e|6.99|2015-01-05 17:29:00|1.4132775322775095|2|8380404721|82|0.6114706929155321|0|58|9983|-80.97058|889|35.03469|NFS-SPARKLING|0.0|13|CB-COOKS BRUT CHAMPAGNE|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|0.61177642288969325|00083804047211|SPARKLING|WINE|-80.97058|1.4132032182494703|82|1
35.03469|5dc674fe04e8a946e50e25a1aba06da9e4425246|4.19|2014-12-21 16:35:00|1.4132775322775095|2|60308424372|82|0.6114706929155321|0|58|3592|-80.97058|1050|35.03469|HAIR STYLING HAIR SPRAY|1.69|17|S/T FRUCTI AERO HAIRSPRAY ULTR|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|0.61177642288969325|00603084260140|HAIR STYLING|HBC|-80.97058|1.4132032182494703|82|1
35.03469|ea2afa5edc03c0e1c7850882e4a998f602783914|6.95|2015-01-24 19:33:00|1.4132775322775095|2|4438606429|82|0.6114706929155321|0|58|3040|-80.97058|1000|35.03469|BRAND-PHYSICIAN FORMULA|0.0|17|PF ORGNICWR BB BTY CRM LGHTMED|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|0.61177642288969325|00044386064300|COSMETICS|HBC|-80.97058|1.4132032182494703|82|1
35.03469|09cd4a154d67adc63bdfca320a3219651d98e263|14.99|2015-01-10 19:12:00|80.970593795509558|2|3410057340|82|35.068500514562629|0|4|455|-80.994596|82|35.061685|DOMESTIC PREMIUM 12PK&>|0.0|16|MILLER LITE 18PK 12OZ CAN|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00034100573409|DOMESTIC BEER|BEER|-80.97058|80.970587132420093|475|1
35.03469|23a193679298cc91f218db4bb6b2f11eb6039a19|13.99|2014-11-29 18:00:00|80.970593795509558|2|1820015981|82|35.068500514562629|0|4|458|-80.994596|82|35.061685|CRAFT BEER|0.0|16|SHOCK TOP 12PK BOTTLES|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00018200159817|DOMESTIC BEER|BEER|-80.97058|80.970587132420093|475|1
35.03469|5a328bebc861a1e816fa023a39f93ae335dc2d02|13.99|2014-10-25 11:18:00|80.970593795509558|2|1820005990|82|35.068500508622286|0|4|456|-80.992182|82|35.103409|DOMESTIC SUPER PREM 12PK&>|0.0|16|MICHELOB ULTRA 12PK 12OZ BTL|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00018200059902|DOMESTIC BEER|BEER|-80.97058|80.970605500300422|88|1
35.03469|ad4ea29e1c66ac8459a0aa4c7180b09d8f6fce02|12.99|2014-09-13 17:06:00|80.970593795509558|2|1820005990|82|35.068500514562629|0|4|456|-80.994596|82|35.061685|DOMESTIC SUPER PREM 12PK&>|0.0|16|MICHELOB ULTRA 12PK 12OZ BTL|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00018200059902|DOMESTIC BEER|BEER|-80.97058|80.970587132420093|475|1
35.03469|ae5e483d64d9ea0d75c146d2b650980465bc52b1|27.98|2014-12-13 14:43:00|80.970593795509558|2|1820005990|82|35.068500514562629|0|4|456|-80.994596|82|35.061685|DOMESTIC SUPER PREM 12PK&>|0.0|16|MICHELOB ULTRA 12PK 12OZ BTL|c56b30d08e6dcaacba6fc70fa5623da4ff7b4169|2.33622494164417|35.073829668338668|00018200059902|DOMESTIC BEER|BEER|-80.97058|80.970587132420093|475|2
34.95459|30d2977e0e51331caab6bf67f8b27b9893c75f7f|1.59|2014-10-17 13:19:00|80.762257539052428|3|78616201000|182|34.985349287328077|0|54|31|-80.850065|4|35.030252|NON CARBONATED WATER|0.59|1|VIT WATER ZERO POWER- C|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00786162003737|BOTTLED WATER|G1 GROCERY|-80.758228|80.758242042658637|470|1
34.95459|0da5e978240b75b80e3a7844f7ea6712be8318c6|2.29|2014-10-27 12:22:00|80.762257539052428|3|78656001621|182|34.985349287328077|0|54|4778|-80.850065|1230|35.030252|BARS-PROTEIN|0.0|17|MET RX CHOC FUDGE 01641|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00786560016414|SPORTS NUTRITIONAL|HBC|-80.758228|80.758242042658637|470|1
34.95459|781a841808481965db613e1b87be543c9bb070d9|0.95|2014-09-19 12:13:00|80.762257539052428|3|61300871771|182|34.985349219985643|0|54|99|-80.80146|32|35.17739|LIQUID TEA|0.0|1|ARIZONA RASPBERRY TEA|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00613008735470|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.758228|80.758307791309576|208|1
34.95459|b5ccdc50cbc3e9730e0d0cc9a923b7303de64236|2.38|2014-11-06 13:14:00|80.762257539052428|3|7433686394|182|34.985349287328077|0|54|342|-80.850065|57|35.030252|FRESH MILK|0.4|3|HUNTER WHOLE MILK 14 OZ|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00074336863943|MILK|DAIRY|-80.758228|80.758242042658637|470|2
34.95459|275208880a820ab4ad272ad628610dbf348243d7|3.99|2014-09-22 12:23:00|80.762257539052428|3|87606300201|182|34.985349219985643|0|54|97|-80.80146|8|35.17739|ENERGY DRINKS|0.5|23|MUSCLE MILK BANANA CREME|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00876063002035|CARBONATED BEVERAGES|BEVERAGE|-80.758228|80.758307791309576|208|1
34.95459|80c6ec63037f535fac294bf3c16e6c6b9bd1c838|7.99|2015-02-01 15:02:00|1.4091206135396188|3|1820012989|182|0.6100726841846847|0|47|457|-80.758228|82|34.95459|DOMESTIC SINGLES/SIX PACKS|0.0|16|MICHELOB ULTRA LIME CACTUS 6PK|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|0.61242566243833529|00018200129896|DOMESTIC BEER|BEER|-80.758228|1.4094969766762753|182|1
34.95459|ac62272893965cbf50faae3b6df9dd6be2701bc1|4.38|2014-11-16 16:26:00|1.4091206135396188|3|7225003106|182|0.6100726841846847|0|47|1031|-80.758228|162|34.95459|ITALIAN|1.38|7|SPOLETTO ITALIAN BREAD|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|0.61242566243833529|00072250031066|SLICED BREAD|COMMERCIAL BAKERY|-80.758228|1.4094969766762753|182|2
34.95459|535f5d84a37c11c10243a946fd2db3ce1140f82a|3.49|2014-11-26 18:43:00|1.4091206135396188|3|4610000107|182|0.6100726841846847|0|47|331|-80.758228|52|34.95459|NATURAL SLICED|0.49|3|SARGENTO DS SHARP CHEDDAR SLIC|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|0.61242566243833529|00046100001134|CHEESE|DAIRY|-80.758228|1.4094969766762753|182|1
34.95459|8c1a4e5478ba2875225eacb82842269eb87b3817|1.69|2014-10-08 12:06:00|80.762257539052428|3|5200033875|182|34.985349287328077|0|54|171|-80.850065|20|35.030252|ISOTONIC DRINKS|0.31|1|GATORADE AM TROPICAL MANGO|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00052000322132|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.758228|80.758242042658637|470|1
34.95459|d83f7a7cd27b805de313f32d2ba592699ffc4639|1.79|2014-11-12 12:21:00|80.762257539052428|3|5200033875|182|34.985349287328077|0|54|171|-80.850065|20|35.030252|ISOTONIC DRINKS|0.9|1|GATORADE G2 GLACIER FREEZE|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00052000320152|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.758228|80.758242042658637|470|1
34.95459|9e54b0e2631bef40f77e44a15a489c548b4c73fc|3.65|2015-01-19 15:33:00|80.762257539052428|3|3800059663|182|34.985349287328077|0|54|61|-80.850065|9|35.030252|RTE CEREAL ADULT|0.0|1|KELLOGG RAISIN BRAN CRUNCH|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00038000870101|CEREAL|G1 GROCERY|-80.758228|80.758242042658637|470|1
34.95459|897f966777c465985b6c401bbd85f3c32658fa7a|0.77|2014-10-03 12:16:00|80.762257539052428|3|7203636010|182|34.985349219985643|0|54|30|-80.80146|4|35.17739|CARBONATED WATER|0.0|1|HT SIMPLY CLEAR PEACH|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00072036360137|BOTTLED WATER|G1 GROCERY|-80.758228|80.758307791309576|208|1
34.95459|7883eaef180741e992f021b762f827ba4a9e51ef|2.39|2014-09-29 12:39:00|80.762257539052428|3|7084781116|182|34.985349219985643|0|54|97|-80.80146|8|35.17739|ENERGY DRINKS|0.0|23|MONSTER KHAOS CAN|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00070847811749|CARBONATED BEVERAGES|BEVERAGE|-80.758228|80.758307791309576|208|1
34.95459|308696b275787075caa41f1a3d458fe01a55a19b|12.49|2014-11-17 10:06:00|1.4091206135396188|3|7185900016|182|0.6100726841846847|0|47|6921|-80.758228|1582|34.95459|BIRD SEED/FEED|0.0|18|KAYTEE GOURMET COCKATIEL DIET|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|0.61242566243833529|00071859000169|PET NEEDS|GM|-80.758228|1.4094969766762753|182|1
34.95459|d8b74b8e8a41cc709f8f36cc48d10495f042f18b|6.59|2014-10-09 16:53:00|80.762257539052428|3|7192196239|182|34.985349287328077|0|54|284|-80.850065|892|35.030252|SUPER PREMIUM PIZZA|0.0|5|DIGIORNO ORIGINAL PEPPERONI|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00071921962395|FROZEN PIZZA|FROZEN|-80.758228|80.758242042658637|470|1
34.95459|adc223342e3efaf819f262ee03538b946220e691|3.38|2014-09-30 12:21:00|80.762257539052428|3|5200033875|182|34.985349219985643|0|54|171|-80.80146|20|35.17739|ISOTONIC DRINKS|0.88|1|GATORADE G2 LEMON LIME|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00052000322514|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.758228|80.758307791309576|208|2
34.95459|7fd93b03720ac78e5d4c892ca74a9b573230433a|4.29|2014-10-21 13:05:00|80.762257539052428|3|2840015636|182|34.985349287328077|0|54|204|-80.850065|31|35.030252|TORTILLA CHIPS|0.0|1|DORITOS BOLD EXPERIMENT RED214|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00028400243346|SNACKS|G1 GROCERY|-80.758228|80.758242042658637|470|1
34.95459|450fe66d7fb3d973c2dbe28a78a0d75838c76563|4.89|2014-09-26 12:03:00|80.762257539052428|3|61126913344|182|34.985349219985643|0|54|97|-80.80146|8|35.17739|ENERGY DRINKS|0.0|23|RED BULL ENERGY 20 OZ|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00611269133448|CARBONATED BEVERAGES|BEVERAGE|-80.758228|80.758307791309576|208|1
34.95459|6f72ff531e982abeb37cb85f54c7c6395970d809|1.49|2014-12-17 11:47:00|80.762257539052428|3|7618316374|182|34.985349274862998|0|54|99|-81.027334|32|34.977331|LIQUID TEA|0.49|1|SNAPPLE ICE TEA|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00076183163740|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.758228|80.758264594589065|149|1
34.95459|27e66589667f65fa09d986b0379ce854b7d0b56b|1.69|2014-09-10 11:36:00|80.762257539052428|3|1200000129|182|34.985349219985643|0|54|55|-80.80146|8|35.17739|REGULAR|0.0|23|CB PEPSI COLA 20 0Z|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00012000001291|CARBONATED BEVERAGES|BEVERAGE|-80.758228|80.758307791309576|208|1
34.95459|2b599b109ba5f2689ceb84951786c71993142645|1.69|2014-09-12 11:37:00|80.762257539052428|3|1200000129|182|34.985349219985643|0|54|55|-80.80146|8|35.17739|REGULAR|0.0|23|CB PEPSI COLA 20 0Z|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00012000001291|CARBONATED BEVERAGES|BEVERAGE|-80.758228|80.758307791309576|208|1
34.95459|97e30160f9040a31b36ffe7948c787b88d630e44|1.0|2014-12-15 12:24:00|80.762257539052428|3|4000000435|182|34.985349274862998|0|54|47|-81.027334|7|34.977331|REGISTER BARS|0.2|1|(FE)SNICKERS CANDY BAR|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00040000424314|CANDY|G1 GROCERY|-80.758228|80.758264594589065|149|1
34.95459|0d7c4a320689658ecaaba70f35b20c1393ffe127|1.69|2015-02-24 13:22:00|80.762257539052428|3|1200000129|182|34.985349219985643|0|54|54|-80.80146|8|35.17739|DIET|0.0|23|CB DIET PEPSI 20 OZ NR|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00012000001307|CARBONATED BEVERAGES|BEVERAGE|-80.758228|80.758307791309576|208|1
34.95459|c3eb6b24631643a9983f5b81e9aea0a6dc8f53cf|3.19|2014-11-25 12:26:00|80.762257539052428|3|1200000180|182|34.985349287328077|0|54|854|-80.850065|32|35.030252|LIQUID ICED COFFEES|0.4|1|FRAPP COFFEE SINGLE|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00012000001802|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.758228|80.758242042658637|470|1
34.95459|09dd7861816e32e534b7ea15a963518852c73c80|1.69|2015-03-06 11:50:00|80.762257539052428|3|1200000129|182|34.985349219985643|0|54|54|-80.80146|8|35.17739|DIET|0.0|23|CB DIET PEPSI 20 OZ NR|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00012000001307|CARBONATED BEVERAGES|BEVERAGE|-80.758228|80.758307791309576|208|1
34.95459|10177315b75e74e1ea7086cc1b17e7501fdb02be|1.69|2015-02-23 12:27:00|80.762257539052428|3|1200000129|182|34.985349219985643|0|54|54|-80.80146|8|35.17739|DIET|0.0|23|CB DIET PEPSI 20 OZ NR|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00012000001307|CARBONATED BEVERAGES|BEVERAGE|-80.758228|80.758307791309576|208|1
34.95459|86ddcb1d8fad31b810f9031fb406bc43a2270012|0.77|2014-10-06 12:52:00|80.762257539052428|3|7203636010|182|34.985349219985643|0|54|30|-80.80146|4|35.17739|CARBONATED WATER|0.0|1|HT SIMPLY CLEAR TANGERINE LIME|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00072036030818|BOTTLED WATER|G1 GROCERY|-80.758228|80.758307791309576|208|1
34.95459|dc170ab3dda56ca6782ce3b15582b96ccbd939a6|1.69|2014-10-01 12:13:00|80.762257539052428|3|5200033875|182|34.985349219985643|0|54|171|-80.80146|20|35.17739|ISOTONIC DRINKS|0.44|1|GATORADE FRUIT PUNCH|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00052000338751|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.758228|80.758307791309576|208|1
34.95459|d9ff646854014bc7ce4f86e3372d7289e5de499a|2.49|2014-10-07 12:09:00|80.762257539052428|3|1200011046|182|34.985349287328077|0|54|97|-80.850065|8|35.030252|ENERGY DRINKS|0.8|23|MT DEW KICKSTART FRUIT PUNCH|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00012000110467|CARBONATED BEVERAGES|BEVERAGE|-80.758228|80.758242042658637|470|1
34.95459|c56f0fa48023bad5e7e63d017c881872f2901955|1.29|2014-11-24 12:15:00|80.762257539052428|3|1657191030|182|34.985349287328077|0|54|30|-80.850065|4|35.030252|CARBONATED WATER|0.29|1|SPARKLING ICE CRISP APPLE|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00016571940379|BOTTLED WATER|G1 GROCERY|-80.758228|80.758242042658637|470|1
34.95459|b69a2e7e0f4b9795fdd53da7430135cffefc0fa3|1.29|2014-12-18 12:20:00|80.762257539052428|3|1657191030|182|34.985349287328077|0|54|30|-80.850065|4|35.030252|CARBONATED WATER|0.29|1|SPARKLING ICE CRISP APPLE|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00016571940379|BOTTLED WATER|G1 GROCERY|-80.758228|80.758242042658637|470|1
34.95459|8abf22c0b368601909ee9491e41ca22c2c278431|1.19|2014-11-20 12:16:00|80.762257539052428|3|8265778540|182|34.985349287328077|0|54|30|-80.850065|4|35.030252|CARBONATED WATER|0.19|1|DEER PRK SPARKLIN LEMON 1L|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00082657710167|BOTTLED WATER|G1 GROCERY|-80.758228|80.758242042658637|470|1
34.95459|b0070a586c2020baf208cb8a5a72650085a2401e|1.19|2014-11-21 11:57:00|80.762257539052428|3|8265778540|182|34.985349287328077|0|54|30|-80.850065|4|35.030252|CARBONATED WATER|0.19|1|DEER PRK SPARKLIN LEMON 1L|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00082657710167|BOTTLED WATER|G1 GROCERY|-80.758228|80.758242042658637|470|1
34.95459|4f373c791426c1d745be65912e09e57c855c8fa8|0.77|2014-10-02 12:06:00|80.762257539052428|3|7203636010|182|34.985349219985643|0|54|30|-80.80146|4|35.17739|CARBONATED WATER|0.0|1|HT SIMPLY CLEAR GRAPE|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00072036360113|BOTTLED WATER|G1 GROCERY|-80.758228|80.758307791309576|208|1
34.95459|1c4cae431ad6502612da56922d6b9cfed44bd482|1.59|2014-11-22 11:42:00|80.762257539052428|3|1200011044|182|34.985349274862998|0|54|97|-81.027334|8|34.977331|ENERGY DRINKS|0.34|23|MT DEW KICKSTART ORANGE CAN|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00012000110443|CARBONATED BEVERAGES|BEVERAGE|-80.758228|80.758264594589065|149|1
34.95459|ac3fbc7f4fde32c2738d23f5b96f4d3bed21777f|4.98|2014-11-05 12:07:00|80.762257539052428|3|1200011044|182|34.985349287328077|0|54|97|-80.850065|8|35.030252|ENERGY DRINKS|1.6|23|MT DEW KICKSTART ORANGE CAN|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00012000110443|CARBONATED BEVERAGES|BEVERAGE|-80.758228|80.758242042658637|470|2
34.95459|fd2ec7f607a7f760adaa9d2b42361225dd21a940|0.77|2015-02-06 12:41:00|80.762257539052428|3|7203636010|182|34.985349219985643|0|54|30|-80.80146|4|35.17739|CARBONATED WATER|0.0|1|HT SPLY CLR RASP/BLACKBERRY|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00072036030801|BOTTLED WATER|G1 GROCERY|-80.758228|80.758307791309576|208|1
34.95459|857e7e539c5cd5bdcd23da90d581204a5eee8c4e|0.77|2015-02-13 12:32:00|80.762257539052428|3|7203636010|182|34.985349219985643|0|54|30|-80.80146|4|35.17739|CARBONATED WATER|0.0|1|HT SPLY CLR RASP/BLACKBERRY|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00072036030801|BOTTLED WATER|G1 GROCERY|-80.758228|80.758307791309576|208|1
34.95459|9c8451844ebfff678b764960e77a9a17809b7c5c|0.77|2015-02-26 12:11:00|80.762257539052428|3|7203636010|182|34.985349219985643|0|54|30|-80.80146|4|35.17739|CARBONATED WATER|0.17|1|HT SPLY CLR RASP/BLACKBERRY|c75edf8bd6ae37840c16b0d92e2e6a6fc8bea6b5|2.1253926220821144|34.983028186791387|00072036030801|BOTTLED WATER|G1 GROCERY|-80.758228|80.758307791309576|208|1
35.28326|e9ddde1049c3af0e5213145db5af92f4f1f6a94a|6.79|2014-12-24 10:39:00|80.66957994482128|4|7203000314|46|35.363825264857752|0|38|1685|-80.605588|385|35.43259|ENTENMANNS (SWEET GOODS)|0.0|14|ENT CHS DANISH TWIST PP|c963ad759c5603ddbfb001fd77bee9067acb8d49|5.56687471986298|35.385064306269825|00072030003146|SWEET GOODS|BAKERY|-80.66939|80.669572196964381|202|1
35.28326|ce838a8c0092a5911cd65e0bba086d081b082668|11.98|2015-01-28 14:31:00|80.66957994482128|4|4470001090|46|35.363825401262211|0|38|838|-80.780702|102|35.318911|PEGS|0.0|19|OSCAR MAYER HARD SALAMI|c963ad759c5603ddbfb001fd77bee9067acb8d49|5.56687471986298|35.385064306269825|00044700010907|LUNCHMEATS|CASE READY MEATS|-80.66939|80.669403382186573|167|2
35.28326|82690e075e14939b510b5c36c7d41781b3bb7d7a|23.38|2015-03-06 13:28:00|80.66957994482128|4|20140400000|46|35.363825264857752|0|38|296|-80.605588|49|35.43259|RANCHER BEEF|9.75|2|BEEF LOIN NY STRIP STEAK BNLS|c963ad759c5603ddbfb001fd77bee9067acb8d49|5.56687471986298|35.385064306269825|00201404000003|BEEF|MEAT|-80.66939|80.669572196964381|202|2
35.28326|914a4b1f0e583526bbfd701aecb8e63124d18866|15.78|2014-11-26 14:40:00|80.66957994482128|4|2770067902|46|35.363825264857752|0|38|265|-80.605588|307|35.43259|FROZEN PIES|3.95|5|M SMITHS ORIG FLAKY CRUST APPL|c963ad759c5603ddbfb001fd77bee9067acb8d49|5.56687471986298|35.385064306269825|00027700679022|DESSERTS FROZEN|FROZEN|-80.66939|80.669572196964381|202|2
34.95459|56b535db3b75fcf3963cf1c6ee998f5014c02050|3.29|2014-12-15 19:19:00|1.4091206135396188|4|1410008786|182|0.6100726841846847|0|47|1035|-80.758228|163|34.95459|SANDWICH ROLL|0.0|7|PEP 100%WHOLE WHEAT HOAGIE PP|ca5ee2c6274d77a0e02ad3b5a3db34f1321008df|1.0281271174619544|0.61242566243833529|00014100090861|BUNS/ROLLS|COMMERCIAL BAKERY|-80.758228|1.4094969766762753|182|1
34.95459|20987e96663735dd3e821e6ce6d7466411519ea6|4.19|2014-11-20 18:37:00|1.4091206135396188|4|2900007325|182|0.6100726841846847|0|47|1149|-80.758228|21|34.95459|PEANUTS|1.19|1|PLNTRS D/R HONEY ROSTD PNUTS|ca5ee2c6274d77a0e02ad3b5a3db34f1321008df|1.0281271174619544|0.61242566243833529|00029000073456|NUTS|G1 GROCERY|-80.758228|1.4094969766762753|182|1
34.95459|5a16f1a31f8808a4aee7b6c807ae47c022a3e8c7|2.19|2014-12-12 15:27:00|1.4091206135396188|4|4900005010|182|0.6100726841846847|0|47|55|-80.758228|8|34.95459|REGULAR|0.2|23|CLASSIC COKE 2 LT CONTOUR|ca5ee2c6274d77a0e02ad3b5a3db34f1321008df|1.0281271174619544|0.61242566243833529|00049000050103|CARBONATED BEVERAGES|BEVERAGE|-80.758228|1.4094969766762753|182|1
34.95459|cf2dc0d916952239815e1e0256d8b30d02e81ae0|4.29|2014-12-24 14:58:00|80.762257539052428|4|2840016014|182|34.969469346409014|0|54|201|-80.8062|31|35.037115|POTATO CHIPS|2.14|1|LAYS WAVY REGULAR|ca5ee2c6274d77a0e02ad3b5a3db34f1321008df|1.0281271174619544|34.983028186791387|00028400160209|SNACKS|G1 GROCERY|-80.758228|80.758239685093272|27|1
34.95459|9e03ace25212d495ebd5d6a14efbd65879747102|1.99|2014-11-17 12:42:00|1.4091206135396188|4|7127923100|182|0.6100726841846847|0|47|555|-80.758228|64|34.95459|PACKAGED SALADS|0.0|4|F.E. BABY SPRING SALAD MIX|ca5ee2c6274d77a0e02ad3b5a3db34f1321008df|1.0281271174619544|0.61242566243833529|00071279231006|FRESH PRODUCE|PRODUCE|-80.758228|1.4094969766762753|182|1
34.95459|500698b3921e38e8898f4e0f1870858c92a23bf7|3.99|2014-12-21 13:42:00|80.762257539052428|4|7022111559|182|34.969469346409014|0|54|727|-80.8062|7|35.037115|SEASONAL CANDY-SINGLE FAC|0.49|1|I/O(C14)TERRYS DRK ORANGE BALL|ca5ee2c6274d77a0e02ad3b5a3db34f1321008df|1.0281271174619544|34.983028186791387|00070221115593|CANDY|G1 GROCERY|-80.758228|80.758239685093272|27|1
35.23102|376616976476cc70b9e9d9a148d514286d216a92|8.97|2014-11-24 16:12:00|80.843809562956082|4|1380004717|205|35.278871196835311|0|37|1278|-80.945176|48|35.323246|SINGLE SERVE NUTRITIONAL|0.0|5|LC CAFE CLSSC PEPPERONI PIZZA|cb04cf0eafb43b4e849c35d8d917a7d5144fe35d|3.3064025562659136|35.255745041786184|00013800047175|FROZEN MEALS|FROZEN|-80.8438|80.8438292336741|166|3
35.23102|e09d66fe4411bd58c18fe7e25d5fbb4ec64e4d03|6.58|2015-01-10 15:58:00|80.843809562956082|4|1380004717|205|35.278871196835311|0|37|1278|-80.945176|48|35.323246|SINGLE SERVE NUTRITIONAL|2.58|5|LC CAFE CLSSC PEPPERONI PIZZA|cb04cf0eafb43b4e849c35d8d917a7d5144fe35d|3.3064025562659136|35.255745041786184|00013800047175|FROZEN MEALS|FROZEN|-80.8438|80.8438292336741|166|2
35.23102|bc7deb5d7869e1ab9619732a727e7fd83721ad3b|11.96|2015-02-08 15:25:00|80.843809562956082|4|1380004717|205|35.278871196835311|0|37|1278|-80.945176|48|35.323246|SINGLE SERVE NUTRITIONAL|0.0|5|LC CAFE CLSSC PEPPERONI PIZZA|cb04cf0eafb43b4e849c35d8d917a7d5144fe35d|3.3064025562659136|35.255745041786184|00013800047175|FROZEN MEALS|FROZEN|-80.8438|80.8438292336741|166|4
35.23102|b5ae4a1b04fa5fa0209cfb21abe80f1ff49f71d1|2.85|2014-10-12 16:12:00|80.843809562956082|4|1380010423|205|35.278871196835311|0|37|1279|-80.945176|48|35.323246|SINGLE SERVE FLAVOR|0.0|5|STOUFFER HARVEST APPLES|cb04cf0eafb43b4e849c35d8d917a7d5144fe35d|3.3064025562659136|35.255745041786184|00013800104236|FROZEN MEALS|FROZEN|-80.8438|80.8438292336741|166|1
35.04711|1e3035a1771bc8098f94fed0d82d0200892f000a|9.08|2014-10-26 13:37:00|80.648225123995502|2|20540500000|129|35.08525247146278|0|30|1832|-80.758228|415|34.95459|BH SLICING CHEESE|0.0|6|BR HD VERMONT CHEDDAR WHITE|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00205405000000|SLICING CHEESE|DELI|-80.64817|80.648238181271381|182|1
35.04711|2b931e1576018899eb7bae4df3908d2f6d093735|3.49|2015-02-22 13:57:00|80.648225123995502|2|7797509132|129|35.08525247146278|0|30|201|-80.758228|31|34.95459|POTATO CHIPS|0.49|1|SOH POPPERS 3  CHEESE|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00077975091432|SNACKS|G1 GROCERY|-80.64817|80.648238181271381|182|1
35.04711|6c435d7b33f52124ccba5b47939718bea56585a2|2.99|2015-02-15 13:03:00|80.648225123995502|2|88810915002|129|35.08525247146278|0|30|1045|-80.758228|173|34.95459|DONUTS|0.49|7|HOSTESS FROSTED MINI DONETTES|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00888109150020|SWEET BAKED GOODS|COMMERCIAL BAKERY|-80.64817|80.648238181271381|182|1
35.04711|f7fd74f656defd07031ee512d83a84a458380a71|3.39|2014-12-14 12:18:00|80.648225123995502|2|5000012734|129|35.08525247146278|0|30|341|-80.758228|57|34.95459|CREAMERS|0.89|3|COFFEEMATE SF FRENCH VANILLA|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00050000848119|MILK|DAIRY|-80.64817|80.648238181271381|182|1
35.04711|6432b6440d0b81eb970ca7d941c7aac7dba367ff|4.29|2015-01-03 12:26:00|80.648225123995502|2|2840006399|129|35.085252435645614|0|30|204|-80.837892|31|34.937113|TORTILLA CHIPS|0.29|1|TOSTITOS HINT OF LIME|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00028400064040|SNACKS|G1 GROCERY|-80.64817|80.648263419592254|372|1
35.04711|8a99a05d56d03bda40cbe50ba3c3d655f889026b|4.29|2014-12-23 16:42:00|80.648225123995502|2|2840006399|129|35.085252435645614|0|30|204|-80.837892|31|34.937113|TORTILLA CHIPS|1.29|1|TOSTITOS HINT OF LIME|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00028400064040|SNACKS|G1 GROCERY|-80.64817|80.648263419592254|372|1
35.04711|bad7920a15f8ed1bfea0aaabccea32ba6461215d|2.39|2014-09-13 11:45:00|80.648225123995502|2|2700038358|129|35.08525247146278|0|30|70|-80.758228|11|34.95459|KETCHUP|0.0|1|HUNTS KETCHUP 35|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00027000383582|CONDIMENTS|G1 GROCERY|-80.64817|80.648238181271381|182|1
35.04711|44d6e8bb3f6e3383c189377d8b849a374e919b66|3.99|2014-11-26 11:56:00|80.648225123995502|2|7203618377|129|35.085252435645614|0|30|887|-80.837892|152|34.937113|SALADS|1.02|12|CRAB QUESO DIP|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00072036183774|SALADS/DIPS|SEAFOOD|-80.64817|80.648263419592254|372|1
35.04711|128916ae178e42875e95b57cfc5a7edd0df5827b|1.69|2014-09-18 16:14:00|80.648225123995502|2|7203626064|129|35.08525247146278|0|30|719|-80.758228|10|34.95459|NFS-COFFEE FILTERS|0.0|1|HT UNBLCHD #4 CONE COFFEE FILT|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00072036260642|COFFEE|G1 GROCERY|-80.64817|80.648238181271381|182|1
35.04711|b941e3e12a4635bfe2ce94e8b5044c19a303ad4e|2.85|2014-11-16 15:46:00|80.648225123995502|2|7203604237|129|35.085252435645614|0|30|41|-80.837892|6|34.937113|BREAKFAST BARS|1.18|1|HT BAR CEREAL APPLE LF|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00072036042385|BREAKFAST FOODS|G1 GROCERY|-80.64817|80.648263419592254|372|1
35.04711|e871b7547039b5367de9c89468ef57a1484786ea|2.85|2014-09-22 17:21:00|80.648225123995502|2|7203604237|129|35.08525247146278|0|30|41|-80.758228|6|34.95459|BREAKFAST BARS|1.18|1|HT BAR CEREAL APPLE LF|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00072036042385|BREAKFAST FOODS|G1 GROCERY|-80.64817|80.648238181271381|182|1
35.04711|816159e0d72331a9241febbe723c89dc11710981|6.79|2014-11-13 16:53:00|80.648225123995502|2|4900002890|129|35.085252435645614|0|30|54|-80.837892|8|34.937113|DIET|6.79|23|DIET COKE W/LIME 12OZ 12PK CAN|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00049000036374|CARBONATED BEVERAGES|BEVERAGE|-80.64817|80.648263419592254|372|1
35.04711|171adfb61b4a24b4f804055770ed8f51a7fd60e4|4.99|2014-10-22 18:51:00|80.648225123995502|2|2301290130|129|35.08525247146278|0|30|1477|-80.758228|485|34.95459|SUSHI HYBRID|0.0|6|CALIFORNIA ROLL SP|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00023012901301|SUSHI|DELI|-80.64817|80.648238181271381|182|1
35.04711|9215024713b51dfd314475ed648c969f21343f1d|4.19|2014-09-14 19:22:00|80.648225123995502|2|4812127620|129|35.085252435645614|0|30|1037|-80.837892|164|34.937113|ENGLISH MUFFINS|2.1|7|THOMAS LITE MULTIGRAIN EM PP|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00048121276201|BREAKFAST|COMMERCIAL BAKERY|-80.64817|80.648263419592254|372|1
35.04711|a8f455dc9c5fcfd5ead2979e675c73e7dc6b3d5b|2.69|2014-11-30 17:43:00|80.648225123995502|2|4114312010|129|35.08525247146278|0|30|119|-80.758228|17|34.95459|RAISINS|0.0|1|SUN MAID 6PK RAISINS|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00041143120101|FRUIT-DRIED|G1 GROCERY|-80.64817|80.648238181271381|182|1
35.04711|28eed0b0c166c7a31ce95118375c3a3e291e7250|3.0|2015-02-01 16:18:00|80.648225123995502|2|4154875084|129|35.085252435645614|0|30|275|-80.837892|45|34.937113|SUPER PREMIUM ICE CREAM|0.0|5|EDY'S SLOW CHURN MINT CHOC CHP|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00041548750804|ICE CREAM|FROZEN|-80.64817|80.648263419592254|372|2
35.04711|e54d045357a1c689460948f6928ad1ea2eb3a281|19.99|2014-11-15 12:22:00|80.648225123995502|2|20496000000|129|35.085252507637279|0|30|755|-80.770346|87|35.052812|NFS-BALLOONS|0.0|9|*BALLOONS|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00204960000005|FLORAL|FLORAL|-80.64817|80.648193009927709|40|1
35.04711|6da5bd6ea727a6ae8b4e9194972716794349d725|1.13|2014-11-23 10:47:00|80.648225123995502|2||129|35.08525247146278|0|30|522|-80.758228|64|34.95459|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00204664000004|FRESH PRODUCE|PRODUCE|-80.64817|80.648238181271381|182|1
35.04711|121be33cb3340f54feb5ff8078e74c1492b9bbd6|4.39|2015-02-28 13:19:00|80.648225123995502|2|5215909004|129|35.085252435645614|0|30|682|-80.837892|61|34.937113|KIDS|0.0|3|YOKIDS  BLUEBERRY STRAW/VAN|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00052159090043|YOGURT|DAIRY|-80.64817|80.648263419592254|372|1
35.04711|adccf559617fe02ea3c5d606595ea5aaa4868885|4.19|2014-10-07 19:59:00|80.648225123995502|2|5215909004|129|35.085252435645614|0|30|682|-80.837892|61|34.937113|KIDS|0.0|3|YOKIDS  BLUEBERRY STRAW/VAN|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00052159090043|YOGURT|DAIRY|-80.64817|80.648263419592254|372|1
35.04711|0ba2246ad516974f3eb6ac3d388ffca01f530227|3.69|2015-01-09 19:26:00|80.648225123995502|2|7033063823|129|35.085252435645614|0|30|8727|-80.837892|1810|34.937113|LIGHTER|0.0|18|(FE)BIC SPECIAL EDITION LGHTER|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00070330638235|LIGHTERS|GM|-80.64817|80.648263419592254|372|1
35.04711|48c4a4ae91727c58ac3504706e90846cffa97c19|2.49|2015-01-20 16:57:00|80.648225123995502|2|7203688085|129|35.08525247146278|0|30|526|-80.758228|64|34.95459|FRESH MUSHROOMS|0.0|4|HT CREMINI MUSHROOMS|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00072036880857|FRESH PRODUCE|PRODUCE|-80.64817|80.648238181271381|182|1
35.04711|5e3fa756c563c06b1fd2be09ca96581d0c262916|13.99|2014-10-24 18:10:00|80.648225123995502|2|75452700024|129|35.08525247146278|0|30|458|-80.758228|82|34.95459|CRAFT BEER|0.0|16|NEW BELGIUM FAT TIRE 12PK|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00754527000240|DOMESTIC BEER|BEER|-80.64817|80.648238181271381|182|1
35.04711|44e9291f7152d40cfa70dfebc2b04a19b4af58de|4.19|2015-02-09 17:09:00|80.648225123995502|2|5215909003|129|35.08525247146278|0|30|690|-80.758228|61|34.95459|ORGANIC|0.0|3|SF YOKIDS CUPS 6PK-STWBRY/BAN|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00052159090036|YOGURT|DAIRY|-80.64817|80.648238181271381|182|1
35.04711|be79ce6d19c962be16cc5c117134aee43e311b12|4.19|2015-03-07 13:24:00|80.648225123995502|2|5215909003|129|35.08525247146278|0|30|690|-80.758228|61|34.95459|ORGANIC|0.0|3|SF YOKIDS CUPS 6PK-STWBRY/BAN|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00052159090036|YOGURT|DAIRY|-80.64817|80.648238181271381|182|1
35.04711|62d90e13839373a0aa2d92f41825959ac1eb8574|4.29|2014-10-22 16:50:00|80.648225123995502|2|4400002796|129|35.085252435645614|0|30|90|-80.837892|13|34.937113|SNACK CRACKERS|1.29|1|TRISCUIT ORIGINAL|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00044000027957|CRACKERS|G1 GROCERY|-80.64817|80.648263419592254|372|1
35.04711|d2605a26e9932668410aa7f63b9b71255b09aa67|7.58|2015-01-27 17:22:00|80.648225123995502|2|4850002013|129|35.085252464316127|0|30|335|-80.97058|56|35.03469|ORANGE JUICE-REGRIGERATED|1.29|3|TROPICANA PP W/CALCIUM|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00048500305690|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.64817|80.648243908613807|82|2
35.04711|bebc5a6cf169062be0cf48d125d27e973425b9a0|4.29|2014-10-18 18:30:00|80.648225123995502|2|5215970117|129|35.08525247146278|0|30|682|-80.758228|61|34.95459|KIDS|0.0|3|YOBABY BLUEBERRY/APPLE|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00052159701154|YOGURT|DAIRY|-80.64817|80.648238181271381|182|1
35.04711|75b2b2ecf46b4cd2259a60f65e27b7c3ef6781c1|2.19|2014-10-23 16:07:00|80.648225123995502|2|5100002549|129|35.08525247146278|0|30|1221|-80.758228|275|34.95459|PASTA SC VALUE|0.0|1|PREGO SC ALFREDO|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00051000197597|PASTA SAUCES|G1 GROCERY|-80.64817|80.648238181271381|182|1
35.04711|3d5e02225e5ac9e05980def21ff6c897d0cf3bdb|3.49|2014-12-30 18:01:00|80.648225123995502|2|7797508161|129|35.08525247146278|0|30|204|-80.758228|31|34.95459|TORTILLA CHIPS|1.74|1|SOH TWST OF LIME TORT CHIPS|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00077975034248|SNACKS|G1 GROCERY|-80.64817|80.648238181271381|182|1
35.04711|8efd65c28d021fa6aaf9941aa6362b5b3d3b68b9|1.0|2015-01-25 16:17:00|80.648225123995502|2|4000000435|129|35.085252435645614|0|30|47|-80.837892|7|34.937113|REGISTER BARS|0.5|1|(FE)M&M PEANUT CANDY|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00040000000327|CANDY|G1 GROCERY|-80.64817|80.648263419592254|372|1
35.04711|ee2c231278b90b5868a22d9254dc6182f2ab7bab|17.92|2014-11-08 17:22:00|80.648225123995502|2|20895500000|129|35.085252435645614|0|30|977|-80.837892|201|34.937113|FRESH HT CHICKEN|2.34|2|HT VALUE PK CHICKEN BNLS BRST|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00208955000001|POULTRY|MEAT|-80.64817|80.648263419592254|372|1
35.04711|19e74ebe3dbd22119abbc7940738883d49568c1b|0.87|2014-10-18 18:32:00|80.648225123995502|2|7203608080|129|35.08525247146278|0|30|120|-80.758228|15|34.95459|COATINGS & BREADERS|0.0|1|HT BREAD CRUMBS ITALIAN|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00072036080813|FLOUR|G1 GROCERY|-80.64817|80.648238181271381|182|1
35.04711|d7c25df10375c95b58be6fe8255cca0d9579cee7|7.58|2014-12-05 17:58:00|80.648225123995502|2|7127930104|129|35.08525247146278|0|30|555|-80.758228|64|34.95459|PACKAGED SALADS|0.0|4|F.E. CAESAR SUPREME COMPLETE|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00071279301044|FRESH PRODUCE|PRODUCE|-80.64817|80.648238181271381|182|2
35.04711|1dfd7b82820becb376346241bd1d24e1bba16c89|7.38|2014-12-04 16:42:00|80.648225123995502|2|1370071016|129|35.085252435645614|0|30|423|-80.837892|72|34.937113|NFS-DISPOSE PLATES/BOWLS|3.38|1|HEFTY PAPER DINER PLATE 10.125|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00013700710162|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.64817|80.648263419592254|372|2
35.04711|30bd60b99ff8f22dc95b62e75bbd7f8cb5d73e63|3.99|2014-12-21 12:55:00|80.648225123995502|2|7203663995|129|35.08525247146278|0|30|342|-80.758228|57|34.95459|FRESH MILK|0.0|3|HARRIS TEETER 2% MILK|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00072036639981|MILK|DAIRY|-80.64817|80.648238181271381|182|1
35.04711|74281b261cb3562f5149b6404df1183f69953de5|4.39|2014-11-29 13:57:00|80.648225123995502|2|7203670269|129|35.085252464316127|0|30|176|-80.97058|72|35.03469|NFS-DISPOSE CUPS|0.89|1|YH PLASTIC CUPS 18OZ|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00072036702692|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.64817|80.648243908613807|82|1
35.04711|34a400682dfb0d246621457514e48ccc246bf008|2.69|2014-12-31 14:26:00|80.648225123995502|2|7800000939|129|35.085252435645614|0|30|55|-80.837892|8|34.937113|REGULAR|0.0|23|VERNONS G ALE 6PK 12 OZ|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00078000009392|CARBONATED BEVERAGES|BEVERAGE|-80.64817|80.648263419592254|372|1
35.04711|7101dc05bcf409a8ff0ef7a791a73922e671eaa7|8.99|2015-01-31 17:35:00|80.648225123995502|2|72383000020|129|35.08525247146278|0|30|458|-80.758228|82|34.95459|CRAFT BEER|0.0|16|LAGUNITAS LIL SUMPIN SUMPIN|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00723830000209|DOMESTIC BEER|BEER|-80.64817|80.648238181271381|182|1
35.04711|65eb9ac020438f455a1435a4879802570b2a56d4|11.15|2015-02-19 20:31:00|80.648225123995502|2|2550000367|129|35.085252507637279|0|30|66|-80.770346|10|35.052812|GROUND CAN|2.16|1|FOLGERS COLOMBIAN CONTAINER|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00025500003856|COFFEE|G1 GROCERY|-80.64817|80.648193009927709|40|1
35.04711|04e672702850de8e86924dbb3f637c010860bb51|3.15|2014-12-11 17:51:00|80.648225123995502|2|7225003706|129|35.08525247146278|0|30|1026|-80.758228|162|34.95459|WHEAT|0.66|7|NATOWN HONEYWHEAT BRD|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00072250037068|SLICED BREAD|COMMERCIAL BAKERY|-80.64817|80.648238181271381|182|1
35.04711|4828470c9556f6c7426c14596f944869ac65fac6|2.27|2014-12-30 17:59:00|80.648225123995502|2|7203656065|129|35.085252507637279|0|30|315|-80.770346|52|35.052812|CHEESE-PROCESSED-SLICED|0.0|3|HT 2% SINGLE WRAP CHEESE|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00072036600844|CHEESE|DAIRY|-80.64817|80.648193009927709|40|1
35.04711|8e5dcf84a657d45f702c8b0416f4efbb9070ef9f|4.65|2015-02-01 16:20:00|80.648225123995502|2|97151|129|35.085252435645614|0|30|1589|-80.837892|369|34.937113|NFS BEVERAGE ESPRESSO|0.0|22|PUMPKIN SPICE LATTE GRANDE|d03d539772fc5944efc7b01f39abc9721bc31afb|2.6355554881544183|35.078006462436761|00000000971510|NFS STARBUCKS|COFFEE SHOP|-80.64817|80.648263419592254|372|1
35.116638|6e52712ef9797fdec2715489034525e94756e70b|1.99|2014-11-09 11:54:00|80.856688219393845|1|7203676376|204|35.138909913350226|0|15|104|-80.825175|16|35.152722|APPLESAUCE-CUPS|0.0|1|HTO 4PK APPLESC NAT|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036763761|FRUIT-CAN/JAR|G1 GROCERY|-80.85753|80.857544209964288|160|1
35.116638|bf71d50525f1da735daf3bc7399e53e72d2d8477|3.98|2015-01-27 15:05:00|80.856688219393845|1|7203676376|204|35.138909916134281|0|15|104|-80.824767|16|35.116751|APPLESAUCE-CUPS|0.0|1|HTO 4PK APPLESC NAT|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036763761|FRUIT-CAN/JAR|G1 GROCERY|-80.85753|80.857534065635704|294|2
35.116638|1a6b56173772b6ac423467857ca4f530a043f95a|1.99|2015-02-18 15:16:00|80.856688219393845|1|7203676376|204|35.138909913350226|0|15|104|-80.825175|16|35.152722|APPLESAUCE-CUPS|0.0|1|HTO 4PK APPLESC NAT|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036763761|FRUIT-CAN/JAR|G1 GROCERY|-80.85753|80.857544209964288|160|1
35.116638|23fde24a7fad163d3978213f8f92256e91b34cb3|3.98|2015-01-01 16:09:00|80.856688219393845|1|7203676415|204|35.138909913350226|0|15|1465|-80.825175|42|35.152722|ORGANIC FROZEN FRUIT|0.0|5|HTO ORGANIC STRAWBERRIES FROZE|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036764157|FROZEN FRUIT|FROZEN|-80.85753|80.857544209964288|160|2
35.116638|960261ae12e1d5c4cae1162f723a18dd88f54e7a|5.97|2014-10-06 13:22:00|80.856688219393845|1|7203676415|204|35.138909913350226|0|15|1465|-80.825175|42|35.152722|ORGANIC FROZEN FRUIT|0.0|5|HTO ORGANIC STRAWBERRIES FROZE|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036764157|FROZEN FRUIT|FROZEN|-80.85753|80.857544209964288|160|3
35.116638|3cc4061f8f5af034bf98e5522d0789690fa48f85|5.97|2014-12-28 09:16:00|80.856688219393845|1|7203676415|204|35.138909913350226|0|15|1465|-80.825175|42|35.152722|ORGANIC FROZEN FRUIT|0.0|5|HTO ORGANIC STRAWBERRIES FROZE|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036764157|FROZEN FRUIT|FROZEN|-80.85753|80.857544209964288|160|3
35.116638|bc7a39b33293c026b65d758b05b2ecd3246bfd5b|1.99|2014-10-17 12:45:00|80.856688219393845|1|7203676376|204|35.138909907643097|0|15|104|-80.80146|16|35.17739|APPLESAUCE-CUPS|0.0|1|HTO 4PK APPLESC NAT|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036763761|FRUIT-CAN/JAR|G1 GROCERY|-80.85753|80.857554124027018|208|1
35.116638|d60fd1609155faf89fb16b8955b8c1c9fc681efc|3.98|2014-10-19 12:47:00|80.856688219393845|1|7203676415|204|35.138909913350226|0|15|1465|-80.825175|42|35.152722|ORGANIC FROZEN FRUIT|0.0|5|HTO ORGANIC STRAWBERRIES FROZE|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036764157|FROZEN FRUIT|FROZEN|-80.85753|80.857544209964288|160|2
35.116638|452bc2de142a64e0b4969508ddf1a3804db79ecf|5.97|2014-11-14 12:02:00|80.856688219393845|1|7203676415|204|35.138909913350226|1|15|1465|-80.825175|42|35.152722|ORGANIC FROZEN FRUIT|0.0|5|HTO ORGANIC STRAWBERRIES FROZE|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036764157|FROZEN FRUIT|FROZEN|-80.85753|80.857544209964288|160|3
35.116638|baca5429a34bc609aa7572ffffea9051df085595|1.99|2014-12-21 11:19:00|80.856688219393845|1|7203676376|204|35.138909913350226|0|15|104|-80.825175|16|35.152722|APPLESAUCE-CUPS|0.0|1|HTO 4PK APPLESC NAT|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036763761|FRUIT-CAN/JAR|G1 GROCERY|-80.85753|80.857544209964288|160|1
35.116638|b585d6432a7256dcc560368ea20739848b3893d5|5.97|2014-09-22 12:37:00|80.856688219393845|1|7203676415|204|35.138909913350226|0|15|1465|-80.825175|42|35.152722|ORGANIC FROZEN FRUIT|0.0|5|HTO ORGANIC STRAWBERRIES FROZE|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036764157|FROZEN FRUIT|FROZEN|-80.85753|80.857544209964288|160|3
35.116638|81e2e3dc19453d944f830af31792489bae004b7b|3.98|2014-11-30 12:34:00|80.856688219393845|1|7203676415|204|35.138909913350226|0|15|1465|-80.825175|42|35.152722|ORGANIC FROZEN FRUIT|0.0|5|HTO ORGANIC STRAWBERRIES FROZE|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036764157|FROZEN FRUIT|FROZEN|-80.85753|80.857544209964288|160|2
35.116638|472409b9b042ff7575e15ee18faa9ad9f0d362af|2.49|2015-01-24 17:14:00|80.856688219393845|1|7203676415|204|35.138909916134281|0|15|1465|-80.824767|42|35.116751|ORGANIC FROZEN FRUIT|0.0|5|HTO ORGANIC STRAWBERRIES FROZE|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036764157|FROZEN FRUIT|FROZEN|-80.85753|80.857534065635704|294|1
35.116638|f0cd7334a01906d94586648d3c873650cf1476b3|5.97|2014-11-02 18:58:00|80.856688219393845|1|7203676376|204|35.138909913350226|0|15|104|-80.825175|16|35.152722|APPLESAUCE-CUPS|0.0|1|HTO 4PK APPLESC NAT|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036763761|FRUIT-CAN/JAR|G1 GROCERY|-80.85753|80.857544209964288|160|3
35.116638|4860482f83835d8d5c9837717814dd5fd1e269b5|4.98|2015-02-13 12:31:00|80.856688219393845|1|7203676415|204|35.138909913350226|0|15|1465|-80.825175|42|35.152722|ORGANIC FROZEN FRUIT|0.0|5|HTO ORGANIC STRAWBERRIES FROZE|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036764157|FROZEN FRUIT|FROZEN|-80.85753|80.857544209964288|160|2
35.116638|71f1ca0f55a371ab6cefbcd1466382f498aaf10c|3.98|2014-10-12 11:58:00|80.856688219393845|1|7203676415|204|35.138909913350226|0|15|1465|-80.825175|42|35.152722|ORGANIC FROZEN FRUIT|0.0|5|HTO ORGANIC STRAWBERRIES FROZE|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036764157|FROZEN FRUIT|FROZEN|-80.85753|80.857544209964288|160|2
35.116638|6538f20e55526c6834bb40d5977a542d9b722da1|1.99|2014-12-07 10:21:00|80.856688219393845|1|7203676376|204|35.138909913350226|0|15|104|-80.825175|16|35.152722|APPLESAUCE-CUPS|0.0|1|HTO 4PK APPLESC NAT|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036763761|FRUIT-CAN/JAR|G1 GROCERY|-80.85753|80.857544209964288|160|1
35.116638|73a1f04a77a1337226f01e601c64cb22b8041dc3|1.99|2015-01-11 18:03:00|80.856688219393845|1|7203676376|204|35.138909913350226|0|15|104|-80.825175|16|35.152722|APPLESAUCE-CUPS|0.0|1|HTO 4PK APPLESC NAT|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036763761|FRUIT-CAN/JAR|G1 GROCERY|-80.85753|80.857544209964288|160|1
35.116638|2b1e0422f66ebb27ad189394bacf21b06dc36f0f|3.98|2014-11-23 11:45:00|80.856688219393845|1|7203676376|204|35.138909913350226|0|15|104|-80.825175|16|35.152722|APPLESAUCE-CUPS|0.0|1|HTO 4PK APPLESC NAT|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036763761|FRUIT-CAN/JAR|G1 GROCERY|-80.85753|80.857544209964288|160|2
35.116638|a0687ac74eda55adb2b1ad8c7829a2487ab8923c|1.99|2014-10-24 14:19:00|80.856688219393845|1|7203676376|204|35.138909913350226|0|15|104|-80.825175|16|35.152722|APPLESAUCE-CUPS|0.0|1|HTO 4PK APPLESC NAT|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036763761|FRUIT-CAN/JAR|G1 GROCERY|-80.85753|80.857544209964288|160|1
35.116638|19da170166d817c19c04f4af43bb7f10e8a36717|5.97|2015-02-02 11:31:00|80.856688219393845|1|7203676376|204|35.138909916134281|0|15|104|-80.824767|16|35.116751|APPLESAUCE-CUPS|0.0|1|HTO 4PK APPLESC NAT|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036763761|FRUIT-CAN/JAR|G1 GROCERY|-80.85753|80.857534065635704|294|3
35.116638|06715d42c9ddc6c24e9b28cf526789631e4cba62|5.97|2014-12-12 16:50:00|80.856688219393845|1|7203676415|204|35.138909913350226|1|15|1465|-80.825175|42|35.152722|ORGANIC FROZEN FRUIT|0.0|5|HTO ORGANIC STRAWBERRIES FROZE|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036764157|FROZEN FRUIT|FROZEN|-80.85753|80.857544209964288|160|3
35.116638|533b3738f2ea376aaac94856eedfebc5e2a2c5d8|3.99|2014-09-19 15:16:00|80.856688219393845|1|75166677005|204|35.138909913350226|0|15|522|-80.825175|64|35.152722|FRESH TOMATOES|1.49|4|NATURESWEET CHERUBS 10.5 OZ|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00751666770058|FRESH PRODUCE|PRODUCE|-80.85753|80.857544209964288|160|1
35.116638|b3e96db735a235388cf85a196f835865606aa371|5.49|2015-02-04 14:59:00|80.856688219393845|1|29424000000|204|35.138909913350226|0|15|561|-80.825175|64|35.152722|FR PROD ORGANIC PRODUCE|0.5|4|ORG BLUEBERRIES 4.4 OZ|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00761635203951|FRESH PRODUCE|PRODUCE|-80.85753|80.857544209964288|160|1
35.116638|d5f82008c1b42b4560eac02f5731c93f07468041|1.39|2014-11-17 13:28:00|80.856688219393845|1|1500007607|204|35.138909916134281|0|15|6|-80.824767|1|35.116751|JARRED BABY FOOD|0.39|1|GERBER 2ND APPLE BLUEBRY|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00015000073473|BABY FOOD|G1 GROCERY|-80.85753|80.857534065635704|294|1
35.116638|cf3dc03ccadb0ad4f031a6da8181eebaa83e42f8|1.39|2014-12-06 08:53:00|80.856688219393845|1|1500007607|204|35.138909913350226|0|15|6|-80.825175|1|35.152722|JARRED BABY FOOD|0.39|1|GERBER 2ND GREEN BEANS 2PK|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00015000073121|BABY FOOD|G1 GROCERY|-80.85753|80.857544209964288|160|1
35.116638|0a575230e578f735519446e6857401e7c707b769|1.39|2015-01-04 14:05:00|80.856688219393845|1|1500007607|204|35.138909916134281|0|15|6|-80.824767|1|35.116751|JARRED BABY FOOD|0.28|1|GERBER 2ND GREEN BEANS 2PK|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00015000073121|BABY FOOD|G1 GROCERY|-80.85753|80.857534065635704|294|1
35.116638|928ccad893557ad27f229bac155b7bcd78a9d7b1|1.39|2015-01-31 15:12:00|80.856688219393845|1|1500007607|204|35.138909913350226|0|15|6|-80.825175|1|35.152722|JARRED BABY FOOD|0.27|1|GERBER 2ND GREEN BEANS 2PK|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00015000073121|BABY FOOD|G1 GROCERY|-80.85753|80.857544209964288|160|1
35.116638|60a7d1393c6e4aec598a510d4c16c1393a537bb2|4.9|2014-11-16 16:28:00|80.856688219393845|1|1450000253|204|35.138909913350226|1|15|1273|-80.825175|50|35.152722|BAG VEG NON STEAM|0.9|5|BE PEPPER STIR FRY|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00014500505637|VEGETABLES-FROZEN|FROZEN|-80.85753|80.857544209964288|160|2
35.116638|20a712b0ec378b79d79738333a2efc8af7418624|5.49|2015-01-06 12:24:00|80.856688219393845|1|29424000000|204|35.138909913350226|0|15|561|-80.825175|64|35.152722|FR PROD ORGANIC PRODUCE|0.0|4|ORG BLUEBERRIES|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00033383222325|FRESH PRODUCE|PRODUCE|-80.85753|80.857544209964288|160|1
35.116638|406fcec42bd4c57af9b4364a5ecfbd96234f1ebb|5.49|2015-02-09 13:54:00|80.856688219393845|1|29424000000|204|35.138909916134281|0|15|561|-80.824767|64|35.116751|FR PROD ORGANIC PRODUCE|0.5|4|ORG BLUEBERRIES|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00033383222325|FRESH PRODUCE|PRODUCE|-80.85753|80.857534065635704|294|1
35.116638|764e5646f95106243439d4428dabe9f08b4ac918|5.49|2015-01-15 11:56:00|80.856688219393845|1|29424000000|204|35.138909913350226|0|15|561|-80.825175|64|35.152722|FR PROD ORGANIC PRODUCE|1.0|4|ORG BLUEBERRIES|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00033383222325|FRESH PRODUCE|PRODUCE|-80.85753|80.857544209964288|160|1
35.116638|2b7d9ecb21a07d5ed55a479765776625f64401fa|5.49|2015-02-22 12:24:00|80.856688219393845|1|29424000000|204|35.138909913350226|0|15|561|-80.825175|64|35.152722|FR PROD ORGANIC PRODUCE|0.0|4|ORG BLUEBERRIES|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00033383222325|FRESH PRODUCE|PRODUCE|-80.85753|80.857544209964288|160|1
35.116638|35f2d69784d826d738f9868f3450b0ac8b65a70c|3.7|2015-03-08 18:13:00|80.856688219393845|1|5150060235|204|35.138909913350226|0|15|10|-80.825175|2|35.152722|LAYER CAKE MIX|1.36|1|PILLS MOIST SUPREME WHITE CAKE|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00051500605905|BAKING MIXES|G1 GROCERY|-80.85753|80.857544209964288|160|2
35.116638|f1ebf5577b661de9469d7ada234a3beb94ea2aa5|6.55|2014-09-28 11:52:00|80.856688219393845|1|5150072001|204|35.138909913350226|0|15|125|-80.825175|19|35.152722|PEANUT BUTTER|0.0|1|JIF NATURAL CREAMY PNUT BUTTER|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00051500243213|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.85753|80.857544209964288|160|1
35.116638|ce791e7a910668a3cabedb5725b4908ee2cddb21|5.99|2014-10-05 13:21:00|80.856688219393845|1|2484232111|204|35.138909913350226|0|15|1885|-80.825175|440|35.152722|PASTA SAUCE|0.0|6|BUITONI PESTO BASIL|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00024842321116|PASTA|DELI|-80.85753|80.857544209964288|160|1
35.116638|a82b90b40873e05b7c6e66d0563444694b0c2ae4|3.38|2015-03-07 17:54:00|80.856688219393845|1|7203698517|204|35.138909916134281|0|15|426|-80.824767|72|35.116751|NFS-PAPER TOWELS|0.71|1|YH ULT TOWEL 1 ROLL WHITE|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036010711|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.85753|80.857534065635704|294|2
35.116638|6a2e5202ab5e07b604e578241c0404b55adcf697|1.34|2014-12-09 14:51:00|80.856688219393845|1|7203653081|204|35.138909913350226|0|15|1275|-80.825175|50|35.152722|BOX VEG|0.0|5|HT CHOPPED SPINACH|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036530813|VEGETABLES-FROZEN|FROZEN|-80.85753|80.857544209964288|160|1
35.116638|c8feb1d95939fa952a1ce32809be7082eb62d803|4.99|2014-10-25 16:13:00|80.856688219393845|1|71575620002|204|35.138909916134281|0|15|504|-80.824767|64|35.116751|FRESH BERRIES|2.5|4|STRAWBERRIES 1LB CLAM|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00715756200023|FRESH PRODUCE|PRODUCE|-80.85753|80.857534065635704|294|1
35.116638|0d081808096515b7228a89e71148045e28e2d946|5.49|2014-12-27 15:14:00|80.856688219393845|1|82704802220|204|35.138909913350226|0|15|331|-80.825175|52|35.152722|NATURAL SLICED|1.5|3|ANDREW EVERERTT SWISS CHEESE|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00827048022203|CHEESE|DAIRY|-80.85753|80.857544209964288|160|1
35.116638|40edc3332d7b44cd8135c3a635cf358f47422736|0.67|2015-02-10 14:53:00|80.856688219393845|1|7203698078|204|35.138909913350226|0|15|242|-80.825175|39|35.152722|CANNED BEANS|0.17|1|HT BEANS BLACK|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036980786|VEGETABLES-CAN/JAR|G1 GROCERY|-80.85753|80.857544209964288|160|1
35.116638|45e6024af3eadbf473a53509f0dfbd9f8ff08d3e|2.01|2014-09-24 13:46:00|80.856688219393845|1|7203698078|204|35.138909913350226|0|15|242|-80.825175|39|35.152722|CANNED BEANS|0.0|1|HT BEANS BLACK|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036980786|VEGETABLES-CAN/JAR|G1 GROCERY|-80.85753|80.857544209964288|160|3
35.116638|546e5fa5a8b54a0b039a9230550af8cd4bf22473|9.99|2015-01-18 15:53:00|80.856688219393845|1|7203678030|204|35.138909913350226|0|15|458|-80.825175|82|35.152722|CRAFT BEER|0.0|16|HT CREATE YOUR OWN SAMPLER|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036780300|DOMESTIC BEER|BEER|-80.85753|80.857544209964288|160|1
35.116638|1e4ba44f1a13986be6d2a951c185eb4ca184efa1|1.69|2015-01-29 15:11:00|80.856688219393845|1|7203688040|204|35.138909916134281|0|15|561|-80.824767|64|35.116751|FR PROD ORGANIC PRODUCE|0.0|4|ORG HT BABY CARROTS 1LB BAG|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036880406|FRESH PRODUCE|PRODUCE|-80.85753|80.857534065635704|294|1
35.116638|4d2916b56fca7396ae6e456d392b387ae3016867|1.69|2015-03-02 13:30:00|80.856688219393845|1|7203688040|204|35.138909916134281|0|15|561|-80.824767|64|35.116751|FR PROD ORGANIC PRODUCE|0.0|4|ORG HT BABY CARROTS 1LB BAG|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036880406|FRESH PRODUCE|PRODUCE|-80.85753|80.857534065635704|294|1
35.116638|9085fffd16ea6c9036436ffc3f42ed11b9cd8a45|1.69|2014-09-15 12:28:00|80.856688219393845|1|7203688040|204|35.138909913350226|0|15|561|-80.825175|64|35.152722|FR PROD ORGANIC PRODUCE|0.19|4|ORG HT BABY CARROTS 1LB BAG|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036880406|FRESH PRODUCE|PRODUCE|-80.85753|80.857544209964288|160|1
35.116638|40e5f13edf769850f9bb79bf54732eba7ab68a28|1.69|2015-01-19 18:09:00|80.856688219393845|1|7203688040|204|35.138909913350226|0|15|561|-80.825175|64|35.152722|FR PROD ORGANIC PRODUCE|0.19|4|ORG HT BABY CARROTS 1LB BAG|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036880406|FRESH PRODUCE|PRODUCE|-80.85753|80.857544209964288|160|1
35.116638|e1a9ded860d240f14798a57693293a3fdc0fbfbb|2.99|2014-12-23 19:03:00|80.856688219393845|1|3338365583|204|35.138909913350226|0|15|522|-80.825175|64|35.152722|FRESH TOMATOES|0.2|4|SWEET GRAPE TOMATO (PINT)|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036880284|FRESH PRODUCE|PRODUCE|-80.85753|80.857544209964288|160|1
35.116638|46bcf7cf80a3e564dfb795b6e0316060f6722b64|4.98|2014-12-01 13:50:00|80.856688219393845|1|3080000920|204|35.138909907643097|0|15|727|-80.80146|7|35.17739|SEASONAL CANDY-SINGLE FAC|0.98|1|I/O(C15)SPNGLR MINI CANES|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00030800009200|CANDY|G1 GROCERY|-80.85753|80.857554124027018|208|2
35.116638|7b638347d5f83d39ebcfc316d262733fbf0d41e3|12.86|2014-12-14 11:32:00|80.856688219393845|1|20250700000|204|35.138909913350226|1|15|642|-80.825175|49|35.152722|NATURAL/ORGANIC BEEF|1.61|2|NATURAL 90% LEAN GRND BF CUSTM|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00202506000007|BEEF|MEAT|-80.85753|80.857544209964288|160|1
35.116638|bc00d1f3e3840fa9abf5f1a313caae3c1f41b31a|2.19|2014-12-17 18:30:00|80.856688219393845|1|7800008246|204|35.138909913350226|0|15|55|-80.825175|8|35.152722|REGULAR|0.33|23|DR PEPPER TEN 2 LITER|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00078000103465|CARBONATED BEVERAGES|BEVERAGE|-80.85753|80.857544209964288|160|1
35.116638|3f81541488fcd4db46ebb3b5b9ecb542b0571ae4|10.28|2014-11-23 11:50:00|80.856688219393845|1|20899300000|204|35.138909913350226|0|15|1419|-80.825175|201|35.152722|SMART CHICKEN ORGANIC|0.0|2|SMART ORGANIC BNLS CHICK BRST|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00208993000001|POULTRY|MEAT|-80.85753|80.857544209964288|160|1
35.116638|9a34d91ce0c68f24dcf067f1291dd6272a353b0b|1.22|2014-11-19 12:44:00|80.856688219393845|1||204|35.138909913350226|0|15|522|-80.825175|64|35.152722|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00204664000004|FRESH PRODUCE|PRODUCE|-80.85753|80.857544209964288|160|1
35.116638|b79ff36a6953b8543f64b9437748af0c7b8073c1|24.99|2015-03-08 16:49:00|80.856688219393845|1||204|35.138909913350226|0|15|565|-80.825175|64|35.152722|REDUCED PRODUCE|0.0|4|PRODUCE REWRAP BY CT|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00204845000007|FRESH PRODUCE|PRODUCE|-80.85753|80.857544209964288|160|1
35.116638|f1b4f2667ad2bb0536b740b81061fba911ac1110|3.85|2015-02-27 12:36:00|80.856688219393845|1|4812127620|204|35.138909916134281|0|15|1037|-80.824767|164|35.116751|ENGLISH MUFFINS|1.93|7|THOMAS 100% WHEAT ENG MUFN PP|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00048121184070|BREAKFAST|COMMERCIAL BAKERY|-80.85753|80.857534065635704|294|1
35.116638|3e7f5c6cf3d15c48801f3b6f3698026c6874bbce|11.99|2014-11-26 13:50:00|80.856688219393845|1|3700086209|204|35.138909913350226|0|15|1205|-80.825175|67|35.152722|NFS-JUMBO DIAPERS|3.0|1|PAMPERS BABY DRY JUMBO SIZE 4|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00037000862116|DISPOSABLE DIAPERS|G1 GROCERY|-80.85753|80.857544209964288|160|1
35.116638|944ce200a9edb7e820d8745e778d3c40d629e279|3.49|2015-01-31 10:48:00|80.856688219393845|1|4460000889|204|35.138909916134281|0|15|400|-80.824767|69|35.116751|NFS-LIQUID CLEANERS|0.0|1|FORMULA 409 A/P ANTI/BAC KITCN|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00044600008882|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.85753|80.857534065635704|294|1
35.116638|b99b3491879be1fd7d8afbfe905ccc67f2537bb8|7.59|2014-12-18 15:47:00|80.856688219393845|1|4850002073|204|35.138909913350226|0|15|335|-80.825175|56|35.152722|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA ORANGE JUICE|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00048500020739|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.85753|80.857544209964288|160|1
35.116638|942a648289f8e33ff24953c9a907965a09c7039f|8.99|2014-10-18 19:56:00|80.856688219393845|1|85375900076|204|35.138909913350226|0|15|458|-80.825175|82|35.152722|CRAFT BEER|0.0|16|SOUTHERN TIER SEASONAL 22OZ|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00853759000766|DOMESTIC BEER|BEER|-80.85753|80.857544209964288|160|1
35.116638|cf61e65284532bef37be31e0cfc3b6a517de653e|4.19|2015-02-08 17:21:00|80.856688219393845|1|30521500700|204|35.138909913350226|0|15|4834|-80.825175|1235|35.152722|COTTON/SWABS|0.0|17|Q-TIPS VALUE PACK-00700|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00305215007005|FIRST AID|HBC|-80.85753|80.857544209964288|160|1
35.116638|f30026bd0c6635fae31148f3c9db568d25c464fd|3.99|2014-09-10 12:32:00|80.856688219393845|1|67729499730|204|35.138909913350226|0|15|184|-80.825175|28|35.152722|SALAD DRESSINGS-LIQUID|0.0|1|CUCINA ANT DRS OG BALSAMICO|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00677294997301|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.85753|80.857544209964288|160|1
35.116638|86e207de028a1a716f1414e61c5492acb38883b3|9.99|2014-12-26 16:25:00|80.856688219393845|1|63848900061|204|35.138909916134281|0|15|458|-80.824767|82|35.116751|CRAFT BEER|0.0|16|DOGFISH HEAD 90 MINUTE IPA 4PK|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00638489000619|DOMESTIC BEER|BEER|-80.85753|80.857534065635704|294|1
35.116638|b0dbc3168da162cb62c5f53dc0916155c1df5058|3.99|2015-02-28 17:37:00|80.856688219393845|1|4610000094|204|35.138909913350226|0|15|333|-80.825175|52|35.152722|PARMESAN CHEESE|2.0|3|SARGENTO ARTISAN PARMESAN|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00046100000595|CHEESE|DAIRY|-80.85753|80.857544209964288|160|1
35.116638|ad1d429a13327f2c2f3368db7d645d9f8f9fe3f1|8.99|2015-02-13 17:35:00|80.856688219393845|1|72383000014|204|35.138909913350226|0|15|458|-80.825175|82|35.152722|CRAFT BEER|0.0|16|LAGUNITAS SEASONAL 6PK|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00723830000148|DOMESTIC BEER|BEER|-80.85753|80.857544209964288|160|1
35.116638|b0996f4e0fbbe1da7081077abce963482590853c|8.99|2015-01-09 18:05:00|80.856688219393845|1|72383000014|204|35.138909913350226|0|15|458|-80.825175|82|35.152722|CRAFT BEER|0.0|16|LAGUNITAS SEASONAL 6PK|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00723830000148|DOMESTIC BEER|BEER|-80.85753|80.857544209964288|160|1
35.116638|44590cc676b11410d88db423f0bf1236d0519582|3.49|2014-10-30 17:32:00|80.856688219393845|1|7797503697|204|35.138909916134281|0|15|199|-80.824767|31|35.116751|DIPS & SALSAS|0.49|1|SOH MILD CHUNKY SALSA|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00077975036976|SNACKS|G1 GROCERY|-80.85753|80.857534065635704|294|1
35.116638|cabfe0cbffaeab44c03b7fa8532e0b98a6b02ea2|9.99|2014-11-29 16:06:00|80.856688219393845|1|8858660384|204|35.138909916134281|0|15|9947|-80.824767|886|35.116751|NFS-PREM-CHARDONNAY|0.0|13|CB-CH ST MICH CHARDONNAY|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00088586603846|PREMIUM ($8-$10.99)|WINE|-80.85753|80.857534065635704|294|1
35.116638|a77eabf9eadfe440c3ec1e0ce6e2f560533ff6ac|1.75|2014-12-16 16:01:00|80.856688219393845|1||204|35.138909916134281|0|15|502|-80.824767|64|35.116751|FRESH BANANAS|0.0|4|BANANAS, YELLOW|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00204011000008|FRESH PRODUCE|PRODUCE|-80.85753|80.857534065635704|294|1
35.116638|54bc08548e44e08c64622a360af4a9fe3f27e2f7|26.99|2014-11-14 16:14:00|80.856688219393845|1|3700086223|204|35.138909916134281|0|15|1206|-80.824767|67|35.116751|NFS-BOX DIAPERS|1.0|1|PAMP BABYDRY SUPER PACK SIZE 4|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00037000862246|DISPOSABLE DIAPERS|G1 GROCERY|-80.85753|80.857534065635704|294|1
35.116638|73bc39b9979b101a003f3c17637627005cfe1498|4.99|2014-12-07 10:22:00|80.856688219393845|1|6827493471|204|35.138909913350226|0|15|31|-80.825175|4|35.152722|NON CARBONATED WATER|2.0|1|NESTLE PURE LIFE .5L 24PK|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00068274934711|BOTTLED WATER|G1 GROCERY|-80.85753|80.857544209964288|160|1
35.116638|aea36e1b05bca98b48af863a26a24ea82b9c6fe9|7.49|2015-02-01 18:06:00|80.856688219393845|1|8600300296|204|35.138909916134281|0|15|9938|-80.824767|885|35.116751|NFS POP PINOT GRS/GRIGIO|0.0|13|WOODBRIDGE PINOT GRIGIO 4PK|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00086003002968|POPULAR (4-$7.99)|WINE|-80.85753|80.857534065635704|294|1
35.116638|a42565f3f4f7738c7e6fce287561d4c8d813d328|1.99|2015-02-24 15:06:00|80.856688219393845|1|3338311008|204|35.138909916134281|0|15|507|-80.824767|64|35.116751|FRESH ORANGES|0.0|4|NAVEL ORANGE, CA 3LB BAG|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00033383119427|FRESH PRODUCE|PRODUCE|-80.85753|80.857534065635704|294|1
35.116638|4132c8c8415fc6d21a39345c1f938f05eddc6f79|15.64|2015-02-09 15:25:00|80.856688219393845|1|20898900000|204|35.138909916134281|0|15|1421|-80.824767|201|35.116751|SMART CHICKEN VEGETABLE FED|0.0|2|SMART CHICKEN BONELESS BREAST|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00208989000008|POULTRY|MEAT|-80.85753|80.857534065635704|294|2
35.116638|a78ea6f0e9a6489faf139d519effe383aed73b2d|7.99|2014-09-27 19:12:00|80.856688219393845|1|70277005801|204|35.138909916134281|0|15|458|-80.824767|82|35.116751|CRAFT BEER|0.0|16|WIDMER UPHEAVAL IPA 6PK|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00702770058013|DOMESTIC BEER|BEER|-80.85753|80.857534065635704|294|1
35.116638|82d1b1f9a4a4b29b32d94d658e7314eb3f461784|17.99|2014-11-11 18:13:00|80.856688219393845|1|4182700012|204|35.138909913350226|0|15|458|-80.825175|82|35.152722|CRAFT BEER|0.0|16|HARPOON MIX PACK 12PK|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00041827000125|DOMESTIC BEER|BEER|-80.85753|80.857544209964288|160|1
35.116638|e3ef94aaf900b94124d7a73018d4590b872a0e54|13.98|2015-01-21 14:06:00|80.856688219393845|1|2370001450|204|35.138909907643097|0|15|291|-80.80146|48|35.17739|FROZEN POUTLRY|0.0|5|TYSON CHICKEN NUGGETS 32OZ|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00023700028471|FROZEN MEALS|FROZEN|-80.85753|80.857554124027018|208|2
35.116638|cbbc77cfd1579e8c0d83aa1c1ee7fab99c85b0c9|11.19|2015-01-25 18:31:00|80.856688219393845|1|5400010060|204|35.138909916134281|0|15|427|-80.824767|72|35.116751|NFS-TOILET TISSUE|3.2|1|SCOTT 1000 WHITE 12 ROLL|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00054000100604|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.85753|80.857534065635704|294|1
35.116638|c57dd12c69408b2b7f6d7689c170c5ea44b0865b|4.49|2014-10-03 18:13:00|80.856688219393845|1|7203601053|204|35.138909913350226|0|15|364|-80.825175|55|35.152722|ORGANIC AND CF EGGS|0.0|3|HTN LG BROWN NEST EGGS|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00072036010537|EGGS FRESH|DAIRY|-80.85753|80.857544209964288|160|1
35.116638|1d5733ad5370d7e40e84cc14b5d8be6184c58d25|3.49|2014-10-05 09:15:00|80.856688219393845|1|664|204|35.138909913350226|0|15|1639|-80.825175|377|35.152722|BULK (DONUTS)|0.0|14|PICK 6  DONUTS|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00000000006640|DONUTS|BAKERY|-80.85753|80.857544209964288|160|1
35.116638|71f2193fde56c405c8d92073d1ccfa0bb24bbe6e|14.99|2015-02-21 16:36:00|80.856688219393845|1|8378316000|204|35.138909916134281|0|15|458|-80.824767|82|35.116751|CRAFT BEER|0.0|16|SIERRA NEVADA SEASONAL|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00083783160000|DOMESTIC BEER|BEER|-80.85753|80.857534065635704|294|1
35.116638|802f693007b72385524e82ebf83d7d931df5d830|9.99|2014-10-31 14:50:00|80.856688219393845|1|9425400015|204|35.138909913350226|0|15|458|-80.825175|82|35.152722|CRAFT BEER|0.0|16|BROOKLYN POST ROAD PUMPKIN 6PK|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00094254000152|DOMESTIC BEER|BEER|-80.85753|80.857544209964288|160|1
35.116638|f865cfdc5ae65c282e81cda2fe64adf997a68a62|7.69|2014-09-23 06:19:00|80.856688219393845|1|30045029604|204|35.138909913350226|0|15|4338|-80.825175|1205|35.152722|PAIN RELIEVER-CHILDREN|0.0|17|CHILD MOTR SUSP BERRY DYE FREE|d4ffaf4a76c42a2f56d1d207e1f8355c8a1df372|1.538935637278362|35.134355925261694|00300450184047|PAIN RELIEF|HBC|-80.85753|80.857544209964288|160|1
35.204336|dee307131534dc8d2947e5dd304de9b5ae96c2ac|3.91|2014-09-29 12:54:00|1.4094857484078087|4|20896500000|61|0.6144315741783704|0|26|977|-80.844274|201|35.204336|FRESH HT CHICKEN|0.0|2|HT FRESH CHICKEN DRUMMETTES|d683a4882eb556107ad43ec337e75f8996bcd18e|2.5089323459178745|0.61471665291522548|00208965000008|POULTRY|MEAT|-80.844274|1.4109987626844462|61|1
35.204336|5dc144e5e14d4e839c7fbbfccae1ddc236970d67|2.27|2014-11-22 15:53:00|80.843945456961976|4|7203605068|61|35.240645982298147|0|59|60|-80.825175|9|35.152722|HOT CEREAL|0.0|1|HT OATS 42 OLD FASHIONED|d683a4882eb556107ad43ec337e75f8996bcd18e|2.5089323459178745|35.232478750868765|00072036050687|CEREAL|G1 GROCERY|-80.844274|80.844294023164821|160|1
35.204336|1f5ed6ea3698b7bc43769b06b6b5df37b01d75c4|1.69|2014-10-06 16:26:00|80.843945456961976|4|4900000044|61|35.240645982298147|0|59|54|-80.825175|8|35.152722|DIET|0.0|23|CB DIET SPRITE ZERO20OZ|d683a4882eb556107ad43ec337e75f8996bcd18e|2.5089323459178745|35.232478750868765|00049000037197|CARBONATED BEVERAGES|BEVERAGE|-80.844274|80.844294023164821|160|1
35.096737|7da939ed5b8338704887250d186c0714dc62b00b|2.69|2014-12-05 20:21:00|80.782094729586973|4|70935100013|30|35.109125110105495|0|27|556|-80.816172|64|35.059823|PACKAGED VEGETABLES|0.0|4|APIO VEGETABLE STIR FRY|d7b277ee713b68fe22a77560f13b2552dcafb2f7|0.8559886108582246|35.102887530186244|00709351000157|FRESH PRODUCE|PRODUCE|-80.78468|80.784687977123795|66|1
35.175855|bc995e4c4f263c59b87a7f6f5a6d05b4eb78f384|1.99|2015-01-19 13:04:00|1.4094857484078087|4|7127915101|218|0.6139344869541099|0|26|555|-80.85013|64|35.175855|PACKAGED SALADS|0.0|4|F.E. SHREDS|d7dc253e6872cf5a30ab6f339087111b8ff7f50d|1.3424785122756886|0.61471665291522548|00071279151014|FRESH PRODUCE|PRODUCE|-80.85013|1.4111009691654428|218|1
35.175855|0799e118952ece687eeeed793a779afbf23a53f0|3.0|2014-09-29 18:32:00|1.4094857484078087|4|5000039758|218|0.6139344869541099|0|26|1147|-80.85013|229|35.175855|HOT COCOA MIX|0.0|1|NESTLE HOT COCOA RCH CHOCOLATE|d7dc253e6872cf5a30ab6f339087111b8ff7f50d|1.3424785122756886|0.61471665291522548|00050000397587|COCOAS CREAMERS SYRUPS|G1 GROCERY|-80.85013|1.4111009691654428|218|2
35.175855|238737a15e03309e16b9d7ee277cbeb729784bb6|3.59|2015-01-03 20:34:00|1.4094857484078087|4|7225002096|218|0.6139344869541099|0|26|1033|-80.85013|163|35.175855|HAMBURGER|0.6|7|CBC WHITE GRINDER SUB ROLL 6PK|d7dc253e6872cf5a30ab6f339087111b8ff7f50d|1.3424785122756886|0.61471665291522548|00072250020961|BUNS/ROLLS|COMMERCIAL BAKERY|-80.85013|1.4111009691654428|218|1
35.175855|c651ff8d49bfcad26719d0bf7d210ee668b920e9|3.59|2015-02-01 15:00:00|1.4094857484078087|4|7225002096|218|0.6139344869541099|0|26|1033|-80.85013|163|35.175855|HAMBURGER|0.6|7|CBC WHITE GRINDER SUB ROLL 6PK|d7dc253e6872cf5a30ab6f339087111b8ff7f50d|1.3424785122756886|0.61471665291522548|00072250020961|BUNS/ROLLS|COMMERCIAL BAKERY|-80.85013|1.4111009691654428|218|1
35.175855|8c044e31d747fe100a587aeb3d17fa4812eeedb7|3.59|2014-12-16 14:23:00|1.4094857484078087|4|7225002096|218|0.6139344869541099|0|26|1033|-80.85013|163|35.175855|HAMBURGER|0.6|7|CBC WHITE GRINDER SUB ROLL 6PK|d7dc253e6872cf5a30ab6f339087111b8ff7f50d|1.3424785122756886|0.61471665291522548|00072250020961|BUNS/ROLLS|COMMERCIAL BAKERY|-80.85013|1.4111009691654428|218|1
35.175855|2276727ab834c4d1d2e3ccf45443ee9a234a219c|3.59|2014-12-12 13:39:00|1.4094857484078087|4|7225002096|218|0.6139344869541099|0|26|1033|-80.85013|163|35.175855|HAMBURGER|0.6|7|CBC WHITE GRINDER SUB ROLL 6PK|d7dc253e6872cf5a30ab6f339087111b8ff7f50d|1.3424785122756886|0.61471665291522548|00072250020961|BUNS/ROLLS|COMMERCIAL BAKERY|-80.85013|1.4111009691654428|218|1
35.175855|9046a09df58e7b03824a4f01b579d90de46c2b2c|3.99|2015-01-27 14:17:00|1.4094857484078087|4|7464100992|218|0.6139344869541099|0|26|562|-80.85013|64|35.175855|FRESH CUT FRUIT|0.0|4|RED APPLE SLICES 14OZ|d7dc253e6872cf5a30ab6f339087111b8ff7f50d|1.3424785122756886|0.61471665291522548|00074641009920|FRESH PRODUCE|PRODUCE|-80.85013|1.4111009691654428|218|1
35.175855|afcc6746a4b3741f9c17cee67df8007a27da167a|3.99|2015-02-06 17:21:00|1.4094857484078087|4|7464100992|218|0.6139344869541099|0|26|562|-80.85013|64|35.175855|FRESH CUT FRUIT|0.0|4|RED APPLE SLICES 14OZ|d7dc253e6872cf5a30ab6f339087111b8ff7f50d|1.3424785122756886|0.61471665291522548|00074641009920|FRESH PRODUCE|PRODUCE|-80.85013|1.4111009691654428|218|1
35.175855|24bcc5ea3ce11f0ede4a6ebde540582f79e9fc5f|8.99|2015-01-05 14:19:00|1.4094857484078087|4|7203688113|218|0.6139344869541099|0|26|583|-80.85013|136|35.175855|NUTS|0.0|4|HT PECAN PIECES TRAY|d7dc253e6872cf5a30ab6f339087111b8ff7f50d|1.3424785122756886|0.61471665291522548|00072036881137|OTHER MERCHANDISE|PRODUCE|-80.85013|1.4111009691654428|218|1
35.175855|0d7fac135574be649c384b4a49f0e5fb319ea7f2|2.19|2015-01-23 12:59:00|1.4094857484078087|4|4900005010|218|0.6139344869541099|0|26|55|-80.85013|8|35.175855|REGULAR|0.2|23|CLASSIC COKE 2 LT CONTOUR|d7dc253e6872cf5a30ab6f339087111b8ff7f50d|1.3424785122756886|0.61471665291522548|00049000050103|CARBONATED BEVERAGES|BEVERAGE|-80.85013|1.4111009691654428|218|1
35.175855|9bfdc954e1973ebb31b60362e6d64f3ff175b9ca|8.58|2014-10-30 20:25:00|1.4094857484078087|4|4400003037|218|0.6139344869541099|0|26|90|-80.85013|13|35.175855|SNACK CRACKERS|2.14|1|WHEAT THINS ORIGINAL|d7dc253e6872cf5a30ab6f339087111b8ff7f50d|1.3424785122756886|0.61471665291522548|00044000030377|CRACKERS|G1 GROCERY|-80.85013|1.4111009691654428|218|2
35.175855|db1e1790becb173d3a9aa7422781a26a1e684bcd|1.69|2015-02-15 20:46:00|1.4094857484078087|4|4900000044|218|0.6139344869541099|0|26|55|-80.85013|8|35.175855|REGULAR|0.0|23|CB COKE SINGLE 20 OZ.|d7dc253e6872cf5a30ab6f339087111b8ff7f50d|1.3424785122756886|0.61471665291522548|00049000000443|CARBONATED BEVERAGES|BEVERAGE|-80.85013|1.4111009691654428|218|1
35.175855|564ca78107a8b12ec4f8fc8cf0b9a63b8f46f471|1.79|2014-12-22 13:23:00|1.4094857484078087|4|73801577742|218|0.6139344869541099|0|26|545|-80.85013|64|35.175855|FRESH SPROUTS|0.0|4|CLOVER SPROUTS, PKG|d7dc253e6872cf5a30ab6f339087111b8ff7f50d|1.3424785122756886|0.61471665291522548|00738015777425|FRESH PRODUCE|PRODUCE|-80.85013|1.4111009691654428|218|1
35.175855|8dbddb443787b3e185d7d1f03ca19994bbf8938f|1.79|2015-02-05 13:39:00|1.4094857484078087|4|73801577742|218|0.6139344869541099|0|26|545|-80.85013|64|35.175855|FRESH SPROUTS|0.0|4|CLOVER SPROUTS, PKG|d7dc253e6872cf5a30ab6f339087111b8ff7f50d|1.3424785122756886|0.61471665291522548|00738015777425|FRESH PRODUCE|PRODUCE|-80.85013|1.4111009691654428|218|1
35.175855|16fa348dc2ad2e10611cf7aed993d16af2a7ca1f|1.79|2014-12-05 13:53:00|1.4094857484078087|4|73801577742|218|0.6139344869541099|0|26|545|-80.85013|64|35.175855|FRESH SPROUTS|0.0|4|CLOVER SPROUTS, PKG|d7dc253e6872cf5a30ab6f339087111b8ff7f50d|1.3424785122756886|0.61471665291522548|00738015777425|FRESH PRODUCE|PRODUCE|-80.85013|1.4111009691654428|218|1
35.175855|8a62b7651935320967a2d984971507c27a1a332c|1.79|2014-12-10 13:27:00|1.4094857484078087|4|73801577742|218|0.6139344869541099|0|26|545|-80.85013|64|35.175855|FRESH SPROUTS|0.0|4|CLOVER SPROUTS, PKG|d7dc253e6872cf5a30ab6f339087111b8ff7f50d|1.3424785122756886|0.61471665291522548|00738015777425|FRESH PRODUCE|PRODUCE|-80.85013|1.4111009691654428|218|1
35.175855|e1f738fdedba92c7c2774cfb3ee8d8ef1c8c2218|1.79|2014-12-31 15:08:00|1.4094857484078087|4|73801577742|218|0.6139344869541099|0|26|545|-80.85013|64|35.175855|FRESH SPROUTS|0.0|4|CLOVER SPROUTS, PKG|d7dc253e6872cf5a30ab6f339087111b8ff7f50d|1.3424785122756886|0.61471665291522548|00738015777425|FRESH PRODUCE|PRODUCE|-80.85013|1.4111009691654428|218|1
35.175855|ea8a0a3b472ac352aa7d024f813ce663ea48f3a8|7.98|2015-01-02 06:28:00|1.4094857484078087|4|7127927100|218|0.6139344869541099|0|26|555|-80.85013|64|35.175855|PACKAGED SALADS|2.0|4|F.E. BABY SPINACH|d7dc253e6872cf5a30ab6f339087111b8ff7f50d|1.3424785122756886|0.61471665291522548|00071279271002|FRESH PRODUCE|PRODUCE|-80.85013|1.4111009691654428|218|2
35.175855|0d4dc774d7594dc3155ce78bf599c833e7eb2e79|3.99|2014-12-07 14:08:00|1.4094857484078087|4|7127927100|218|0.6139344869541099|0|26|555|-80.85013|64|35.175855|PACKAGED SALADS|0.99|4|F.E. BABY SPINACH|d7dc253e6872cf5a30ab6f339087111b8ff7f50d|1.3424785122756886|0.61471665291522548|00071279271002|FRESH PRODUCE|PRODUCE|-80.85013|1.4111009691654428|218|1
35.175855|afbb93210c9b535859bc0a24c76250e9a2bc6468|1.69|2014-09-20 13:18:00|1.4094857484078087|4|7203688003|218|0.6139344869541099|0|26|527|-80.85013|64|35.175855|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|d7dc253e6872cf5a30ab6f339087111b8ff7f50d|1.3424785122756886|0.61471665291522548|00072036880031|FRESH PRODUCE|PRODUCE|-80.85013|1.4111009691654428|218|1
35.175855|714f04a19d61bb08f6397688a0ccf6e544fe1a34|7.3500000000000005|2014-10-31 20:29:00|1.4094857484078087|4|1450000253|218|0.6139344869541099|0|26|1272|-80.85013|50|35.175855|BAG VEG STEAM|0.78|5|BE STEAMFRESH PREM BRUSS SPRTS|d7dc253e6872cf5a30ab6f339087111b8ff7f50d|1.3424785122756886|0.61471665291522548|00014500011589|VEGETABLES-FROZEN|FROZEN|-80.85013|1.4111009691654428|218|3
35.175855|0e88d0101c98ae2592c2b4d1005268251ad3c821|2.49|2014-12-19 11:31:00|1.4094857484078087|4|7203670298|218|0.6139344869541099|0|26|728|-80.85013|72|35.175855|NFS-PLASTIC FLATWARE|0.0|1|YH EVERYDAY HD SPOONS|d7dc253e6872cf5a30ab6f339087111b8ff7f50d|1.3424785122756886|0.61471665291522548|00072036702982|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.85013|1.4111009691654428|218|1
35.28326|f88d9ec6c9febda0e5e7fb8a6fdd830d5f5cc625|10.38|2014-09-15 12:34:00|1.4094857484078087|2|20895300000|46|0.6158090578372145|0|26|977|-80.66939|201|35.28326|FRESH HT CHICKEN|0.0|2|HT FRESH BNLS CHICKEN BREAST|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00208953000003|POULTRY|MEAT|-80.66939|1.4079464610753885|46|1
35.28326|399ee9566f0e1fb9fad3bf345acb1dd5d3fc89c4|58.779999999999994|2015-01-07 20:38:00|1.4094857484078087|2|20895300000|46|0.6158090578372145|0|26|977|-80.66939|201|35.28326|FRESH HT CHICKEN|6.15|2|HT FRESH BNLS CHICKEN BREAST|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00208953000003|POULTRY|MEAT|-80.66939|1.4079464610753885|46|6
35.28326|6624e5bac06393d7a9d9a8b00fd73e7376294b57|8.99|2014-11-16 16:19:00|80.669414401537693|2|63123430002|46|35.309074955099199|0|19|458|-80.662946|82|35.412407|CRAFT BEER|0.0|16|SWEETWATER 420 PALE ALE 6PK|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|35.305725790410776|00631234300026|DOMESTIC BEER|BEER|-80.66939|80.669433417044175|68|1
35.28326|2e6be6f8ae5e3d043a7ccb64f86e21302f3bba65|8.99|2014-11-24 13:38:00|80.669414401537693|2|71280823275|46|35.309074955099199|0|19|458|-80.662946|82|35.412407|CRAFT BEER|0.0|16|HIGHLANDS KASHMIR 6PK IPA|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|35.305725790410776|00712808232759|DOMESTIC BEER|BEER|-80.66939|80.669433417044175|68|1
35.28326|d34f8e33af45a1668ac10b238190ada270a6c882|2.99|2014-12-23 18:43:00|1.4094857484078087|2|88810915004|46|0.6158090578372145|0|26|1045|-80.66939|173|35.28326|DONUTS|1.5|7|HOSTESS POWERED MINI DONETTES|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00888109150044|SWEET BAKED GOODS|COMMERCIAL BAKERY|-80.66939|1.4079464610753885|46|1
35.28326|d9579d803b3d1c1c6530b350d61c91ced75a4e7c|12.19|2014-11-04 16:05:00|1.4094857484078087|2|1380023260|46|0.6158090578372145|0|26|1280|-80.66939|48|35.28326|MULTI SERVE MEALS|3.72|5|STOUFF FIESTA BAKE LRG FAMILY|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00013800312273|FROZEN MEALS|FROZEN|-80.66939|1.4079464610753885|46|1
35.28326|f38d9ab0549b1b39aabdf1bfc4487bac6b08704a|12.99|2014-11-29 16:28:00|80.669414401537693|2|2124212009|46|35.309074955099199|0|19|458|-80.662946|82|35.412407|CRAFT BEER|0.0|16|REDHOOK SAMPLER 12PK|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|35.305725790410776|00021242120097|DOMESTIC BEER|BEER|-80.66939|80.669433417044175|68|1
35.28326|81e762e26ab74a067b178b146d8fbdcf2fabcb75|2.89|2015-03-09 14:31:00|1.4094857484078087|2|7203655029|46|0.6158090578372145|0|26|331|-80.66939|52|35.28326|NATURAL SLICED|0.92|3|HT MEDIUM CHEDDAR SLICES|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00072036983930|CHEESE|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|e376648ddc6916ab40346a47d2b75038a7eaac8f|1.77|2015-02-01 14:07:00|1.4094857484078087|2|7203698067|46|0.6158090578372145|0|26|365|-80.66939|56|35.28326|REFRIGERATED TEAS|0.78|3|HARRIS TEETER UNSWEET TEA|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00072036982742|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|c442bd8b1e827ce684a9a75a45df716f7f48f8b6|1.77|2015-02-01 16:19:00|80.669414401537693|2|7203698067|46|35.309074955099199|0|19|365|-80.662946|56|35.412407|REFRIGERATED TEAS|0.78|3|HARRIS TEETER UNSWEET TEA|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|35.305725790410776|00072036982742|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.66939|80.669433417044175|68|1
35.28326|e79c93162771a8414eaebee79856500e7894146e|3.79|2015-02-04 17:22:00|1.4094857484078087|2|7203688014|46|0.6158090578372145|0|26|581|-80.66939|136|35.28326|FRESH SALSA|0.0|4|HT FRESH MEDIUM SALSA|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00072036880222|OTHER MERCHANDISE|PRODUCE|-80.66939|1.4079464610753885|46|1
35.28326|1f6bfc69f4b6e2cab4ef951fc17b22b0c78a7358|3.29|2014-10-17 14:06:00|1.4094857484078087|2|7203695076|46|0.6158090578372145|0|26|1609|-80.66939|371|35.28326|TAKE & BAKE BREAD|1.3|14|TAKE & BAKE SMALL WHEAT FRENCH|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00072036950765|BREAD|BAKERY|-80.66939|1.4079464610753885|46|1
35.28326|4ab697d2191d4a506e368bd7fe0901ff31130617|1.79|2015-01-22 19:49:00|1.4094857484078087|2|7203688032|46|0.6158090578372145|0|26|555|-80.66939|64|35.28326|PACKAGED SALADS|0.0|4|HT SHREDDED ICEBERG LETTUCE|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00072036880321|FRESH PRODUCE|PRODUCE|-80.66939|1.4079464610753885|46|1
35.28326|46625ac0c1def93fe7d2f81ab9e868433e43310b|3.39|2014-12-14 14:29:00|80.669414401537693|2|7550000011|46|35.309074955099199|0|19|76|-80.662946|11|35.412407|MEAT SAUCES|0.0|1|TEXAS PETE WING BUFFALO|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|35.305725790410776|00075500000119|CONDIMENTS|G1 GROCERY|-80.66939|80.669433417044175|68|1
35.28326|9a000512c06486cad9c2f275a57e32c5ede62057|3.89|2014-12-01 17:09:00|1.4094857484078087|2|7247000222|46|0.6158090578372145|0|26|1641|-80.66939|377|35.28326|PACKAGED DONUTS|0.0|14|K K 6 ORIG GLAZED DONUT  PP|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00072470002228|DONUTS|BAKERY|-80.66939|1.4079464610753885|46|1
35.28326|587ec4531a0ab964d5863a9f85d7b521c1d4881a|3.39|2015-01-03 16:07:00|80.669414401537693|2|7550000011|46|35.309074955099199|0|19|76|-80.662946|11|35.412407|MEAT SAUCES|0.0|1|TEXAS PETE WING BUFFALO|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|35.305725790410776|00075500000119|CONDIMENTS|G1 GROCERY|-80.66939|80.669433417044175|68|1
35.28326|46316d97723afbff38bec992f988b365de279f48|3.69|2014-11-07 11:59:00|1.4094857484078087|2|7797508822|46|0.6158090578372145|0|26|202|-80.66939|31|35.28326|PRETZELS|0.69|1|SOH BBQ PRETZEL PIECES|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00077975091364|SNACKS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|69ee2281ecbf8c69becc6cf78bf0f7bce47e8767|7.99|2015-01-30 22:20:00|1.4094857484078087|2|8382012360|46|0.6158090578372145|0|26|459|-80.66939|83|35.28326|IMPORT BEER|0.0|16|GUINNESS DRFT 4PK 14.9OZ CAN|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00083820123609|IMPORT BEER|BEER|-80.66939|1.4079464610753885|46|1
35.28326|2afa401ddc85c234d46fb169aba49358df364006|8.49|2014-10-02 13:42:00|1.4094857484078087|2|2301200013|46|0.6158090578372145|0|26|1477|-80.66939|485|35.28326|SUSHI HYBRID|0.0|6|PLUS ROLL|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00023012000134|SUSHI|DELI|-80.66939|1.4079464610753885|46|1
35.28326|52aeb73288fae152266c84cd8adeb02ed489d005|1.79|2015-02-17 17:10:00|1.4094857484078087|2|1799259110|46|0.6158090578372145|0|26|555|-80.66939|64|35.28326|PACKAGED SALADS|0.0|4|CHEF BUDDY DICED CAB/CARROT|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00017992591102|FRESH PRODUCE|PRODUCE|-80.66939|1.4079464610753885|46|1
35.28326|e711e6d4feebe60b062e03d0ba34dbcc521ff4f0|4.19|2014-10-14 12:24:00|1.4094857484078087|2|2100062503|46|0.6158090578372145|0|26|318|-80.66939|52|35.28326|SHREDDED/GRATED CHEESE|1.69|3|KRAFT FINELY SHREDDED SHARP C|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00021000638741|CHEESE|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|8362360f0ef69bc3a0f34958a5b60ef7432a8896|2.79|2015-02-19 17:24:00|1.4094857484078087|2|2740010307|46|0.6158090578372145|0|26|313|-80.66939|51|35.28326|MARGARINE|0.0|3|COUNTRY CROCK PLUS CALCIUM|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00027400800245|BUTTER & MARGARINE|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|fcd62711dc9c1968df7f2416b6800138caddca70|13.58|2014-10-31 11:23:00|1.4094857484078087|2|4900002890|46|0.6158090578372145|0|26|54|-80.66939|8|35.28326|DIET|3.4|23|VANILLA COKE ZERO 12PK CAN|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00049000048254|CARBONATED BEVERAGES|BEVERAGE|-80.66939|1.4079464610753885|46|2
35.28326|84219350cac60b0755e49af75d7af0923fb24261|4.69|2014-11-19 13:27:00|1.4094857484078087|2|4900002468|46|0.6158090578372145|0|26|54|-80.66939|8|35.28326|DIET|4.69|23|DIET COKE .5 LITER/6 PK.|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.66939|1.4079464610753885|46|1
35.28326|c2d4f6d6945669754db6946409914aef6e7d2308|2.65|2014-10-28 10:32:00|1.4094857484078087|2|4119601000|46|0.6158090578372145|0|26|1201|-80.66939|33|35.28326|RTS CANNED|0.0|1|PROG TRAD CHK CHEESE ENCHILADA|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00041196915136|SOUP|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|bcc7a8d33dff9f45948a7af905842ad0d1367145|5.97|2014-09-26 11:20:00|1.4094857484078087|2|3800084496|46|0.6158090578372145|0|26|201|-80.66939|31|35.28326|POTATO CHIPS|1.47|1|PRINGLES PIZZA|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00038000845024|SNACKS|G1 GROCERY|-80.66939|1.4079464610753885|46|3
35.28326|e726bba1b3d5b5c5127acf06c83807809d81ef90|4.69|2014-12-14 13:14:00|80.669414401537693|2|4900002468|46|35.309074955099199|0|19|55|-80.662946|8|35.412407|REGULAR|0.0|23|M. MAID LEMONADE .5L 6 PK|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|35.305725790410776|00025000058288|CARBONATED BEVERAGES|BEVERAGE|-80.66939|80.669433417044175|68|1
35.28326|d240b3f72fb4e52eb52c2d0fad06a1616006d9b8|5.98|2014-10-03 11:20:00|1.4094857484078087|2|2560000786|46|0.6158090578372145|0|26|1046|-80.66939|173|35.28326|CAKES|0.99|7|TSTYKAKE CHOC BAG DNTS|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00025600007877|SWEET BAKED GOODS|COMMERCIAL BAKERY|-80.66939|1.4079464610753885|46|2
35.28326|4b2978c08e025a01d500d3eabaa5c4523829bfdd|0.7|2015-01-06 17:55:00|1.4094857484078087|2||46|0.6158090578372145|0|26|522|-80.66939|64|35.28326|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00204664000004|FRESH PRODUCE|PRODUCE|-80.66939|1.4079464610753885|46|1
35.28326|8be1786155aa30e98fe5708ba7b3ea1e62d2242a|4.69|2014-10-11 11:00:00|80.669414401537693|2|4210000900|46|35.309074955099199|0|19|490|-80.662946|93|35.412407|NFS-INSECTICIDES, ETC|0.0|1|HOT SHOT WASP&HORNET|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|35.305725790410776|00042100009002|INSECTICIDES/PESTICIDES/RODENT|G1 GROCERY|-80.66939|80.669433417044175|68|1
35.28326|44a287eaae7b8ce64eb8b8e3429705407f527f6d|7.99|2015-03-01 20:05:00|1.4094857484078087|2|5200020805|46|0.6158090578372145|0|26|171|-80.66939|20|35.28326|ISOTONIC DRINKS|2.99|1|GATORADE FRUIT PUNCH 8PK|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00052000208061|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|ce9583f9ad4bcfd93ded4c4fcd240522f264e381|7.99|2014-10-07 14:22:00|1.4094857484078087|2|5200020805|46|0.6158090578372145|0|26|171|-80.66939|20|35.28326|ISOTONIC DRINKS|4.0|1|GATORADE FRUIT PUNCH 8PK|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00052000208061|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|d23bb165757ebb651a0b7d14419a03e569c2f039|15.98|2015-01-24 15:29:00|1.4094857484078087|2|5200020805|46|0.6158090578372145|0|26|171|-80.66939|20|35.28326|ISOTONIC DRINKS|5.98|1|GATORADE FRUIT PUNCH 8PK|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00052000208061|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.66939|1.4079464610753885|46|2
35.28326|d20d957ee7bc063791140ee24f47623f3001a03c|1.89|2014-11-24 09:30:00|80.669414401537693|2|5150020430|46|35.309074955099199|0|19|101|-80.662946|15|35.412407|FLOUR-ALL PURPOSE|0.0|1|PILLSBURY ALL PURPOSE FLOUR|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|35.305725790410776|00051500204306|FLOUR|G1 GROCERY|-80.66939|80.669433417044175|68|1
35.28326|9e4a883ec25f8112eaad43ee7b91804006bb5e16|2.99|2014-10-29 08:23:00|1.4094857484078087|2|7203695121|46|0.6158090578372145|0|26|1629|-80.66939|373|35.28326|TAKE & BAKE ROLLS|0.0|14|TAKE & BAKE WHEAT PETIT PN RL|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00072036951212|ROLLS|BAKERY|-80.66939|1.4079464610753885|46|1
35.28326|a0f7bddfd9857eadf41532d3b5ffa4b4251d49dc|10.98|2015-02-25 13:16:00|1.4094857484078087|2|7597140209|46|0.6158090578372145|0|26|1845|-80.66939|425|35.28326|FFM PRESLICED CHEESE|0.0|6|F.F.COLBY JACK CHEDDAR  CHEESE|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00072036010315|PRESLICED CHEESE|DELI|-80.66939|1.4079464610753885|46|2
35.28326|05790f25797553a7c754497f0b1b0eea352a2e91|0.75|2015-02-24 16:51:00|1.4094857484078087|2|7203641055|46|0.6158090578372145|0|26|257|-80.66939|39|35.28326|TOMATOES|0.25|1|HT TOMATOES PETITE DICED|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00072036410726|VEGETABLES-CAN/JAR|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|87478a502e7ece215a07ea6a5089814844da28ba|0.75|2015-02-15 21:09:00|1.4094857484078087|2|7203641055|46|0.6158090578372145|0|26|257|-80.66939|39|35.28326|TOMATOES|0.15|1|HT TOMATOES PETITE DICED|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00072036410726|VEGETABLES-CAN/JAR|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|0891ec89d6312f0a6f6543456df75677ab1819d0|7.99|2014-12-29 20:43:00|1.4094857484078087|2|7203676196|46|0.6158090578372145|0|26|36|-80.66939|10|35.28326|PREMIUM GROUND|2.42|1|HT TRADER COFFEE DEC G COLUMBN|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00072036761996|COFFEE|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|848fb787448605d511c68c72be43d82585f36935|23.97|2015-01-25 17:50:00|1.4094857484078087|2|7203676196|46|0.6158090578372145|0|26|36|-80.66939|10|35.28326|PREMIUM GROUND|0.0|1|HT TRADER COFFEE DEC G COLUMBN|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00072036761996|COFFEE|G1 GROCERY|-80.66939|1.4079464610753885|46|3
35.28326|abcc4e41f6d67a30f8910317a48a1c016e164e6c|23.97|2015-01-26 16:08:00|80.669414401537693|2|7203676196|46|35.309074979060284|0|19|36|-80.737839|10|35.297134|PREMIUM GROUND|0.0|1|HT TRADER COFFEE DEC G COLUMBN|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|35.305725790410776|00072036761996|COFFEE|G1 GROCERY|-80.66939|80.669395283861164|258|3
35.28326|7f4cd7c1fd643a68d00a2197095641d6c4ca82d3|5.98|2015-01-23 18:23:00|1.4094857484078087|2|7203695360|46|0.6158090578372145|0|26|1629|-80.66939|373|35.28326|TAKE & BAKE ROLLS|0.0|14|TAKE & BAKE PETITE PN RL 6 CT|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00072036953605|ROLLS|BAKERY|-80.66939|1.4079464610753885|46|2
35.28326|5db908b65d41d843eaa7e270f27c060a18e78936|1.99|2014-10-12 12:33:00|80.669414401537693|2|7203698370|46|35.309074955099199|0|19|205|-80.662946|31|35.412407|REMAINING SNACKS|0.49|1|HT SNACK MIX TRADITIONAL|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|35.305725790410776|00072036983701|SNACKS|G1 GROCERY|-80.66939|80.669433417044175|68|1
35.28326|d23fb3e17fd736c8deebe78754b927ea60d7d853|6.69|2015-02-01 16:19:00|80.669414401537693|2|4670462065|46|35.309074955099199|0|19|1277|-80.662946|279|35.412407|FROZEN SNACKS|0.0|5|TGIF MOZZARELLA STICKS|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|35.305725790410776|00046704620908|FROZEN SANDWICH AND SNACKS|FROZEN|-80.66939|80.669433417044175|68|1
35.28326|666ed830ac271e36e2ba9efc14f88394f9679d6c|11.99|2014-11-02 12:43:00|1.4094857484078087|2|7203663048|46|0.6158090578372145|0|26|297|-80.66939|49|35.28326|GROUND BEEF|1.0|2|93% LEAN GROUND BEEF 2 LB|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00072036630483|BEEF|MEAT|-80.66939|1.4079464610753885|46|1
35.28326|97ed71ca7cf504a8f35130115df45aa8c0a83e5f|113.88|2015-01-04 16:21:00|80.669414401537693|2|202108000000|46|35.309074979060284|0|19|299|-80.737839|49|35.297134|ANGUS BEEF|31.65|2|ANGUS TENDERLON WHOLE CUSTOM|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|35.305725790410776|02021080000009|BEEF|MEAT|-80.66939|80.669395283861164|258|1
35.28326|8921464adfd4736b5d9b707e5a2092a8539031fa|13.58|2014-12-17 16:00:00|1.4094857484078087|2|4900002890|46|0.6158090578372145|0|26|55|-80.66939|8|35.28326|REGULAR|0.0|23|MELLO YELLO 12OZ 12PK FP CN|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00049000028935|CARBONATED BEVERAGES|BEVERAGE|-80.66939|1.4079464610753885|46|2
35.28326|795cac533116171b23ab50cd1f0af928a5faf467|6.79|2014-09-20 19:25:00|1.4094857484078087|2|4900002890|46|0.6158090578372145|0|26|55|-80.66939|8|35.28326|REGULAR|3.4|23|MELLO YELLO 12OZ 12PK FP CN|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00049000028935|CARBONATED BEVERAGES|BEVERAGE|-80.66939|1.4079464610753885|46|1
35.28326|33ea1a16908740288abfd67d8a5b86f3df5f6fc9|3.69|2015-01-25 17:13:00|80.669414401537693|2|7518500003|46|35.309074979060284|0|19|1033|-80.737839|163|35.297134|HAMBURGER|0.0|7|MARTIN'S POTATO SANDWICH ROLLS|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|35.305725790410776|00075185000039|BUNS/ROLLS|COMMERCIAL BAKERY|-80.66939|80.669395283861164|258|1
35.28326|386a32a30c59c1d5e4d76a813f2007b3661cb331|4.29|2015-02-23 12:39:00|1.4094857484078087|2|2840016014|46|0.6158090578372145|0|26|201|-80.66939|31|35.28326|POTATO CHIPS|2.15|1|LAYS CLASSIC|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00028400160148|SNACKS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|9e96dd2e2f61fb146d98c0c862e19dc10998c3ed|4.29|2015-02-05 17:13:00|1.4094857484078087|2|2840016014|46|0.6158090578372145|0|26|201|-80.66939|31|35.28326|POTATO CHIPS|0.29|1|LAYS CLASSIC|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00028400160148|SNACKS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|fc7827699faab544a6f21c94e95e15b74fa43c56|6.87|2015-01-15 18:43:00|1.4094857484078087|2|7203601991|46|0.6158090578372145|0|26|1277|-80.66939|279|35.28326|FROZEN SNACKS|1.15|5|HT MINI PIZZA BAGELS PEPPERONI|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00072036019912|FROZEN SANDWICH AND SNACKS|FROZEN|-80.66939|1.4079464610753885|46|3
35.28326|0c62ae218f34f9369b2032b7cf9a09332311ae22|5.98|2014-12-13 16:33:00|1.4094857484078087|2|7203670465|46|0.6158090578372145|0|26|729|-80.66939|69|35.28326|NFS-SCOUR PAD/STEEL WOOL|1.98|1|YH X-STRENGTH CLEANING ERASERS|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00072036704658|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.66939|1.4079464610753885|46|2
35.28326|dbb672f6c58a4b2aa1a5cf364a736394900ba806|1.5|2015-02-01 15:55:00|1.4094857484078087|2|7203663107|46|0.6158090578372145|0|26|1262|-80.66939|57|35.28326|HALF N HALF WHIPPING CREAM|0.0|3|HT HALF & HALF|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00072036632036|MILK|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|405a865636897e23062f59d0498e290bfd37ad51|9.99|2015-01-16 17:46:00|1.4094857484078087|2|2370001118|46|0.6158090578372145|0|26|291|-80.66939|48|35.28326|FROZEN POUTLRY|2.0|5|TYSON ANTY GRILL WINGS ROTISS|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00023700037756|FROZEN MEALS|FROZEN|-80.66939|1.4079464610753885|46|1
35.28326|54b3abd45c596fbf3d64d60dbdba3a48d7db79e4|3.49|2014-12-02 16:22:00|80.669414401537693|2|2840008294|46|35.309074979060284|0|19|201|-80.737839|31|35.297134|POTATO CHIPS|0.99|1|LAYS KETTLE BBQ|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|35.305725790410776|00028400082938|SNACKS|G1 GROCERY|-80.66939|80.669395283861164|258|1
35.28326|0569c018e39c1f14f225220982b2adc8ef99f7e9|2.77|2014-10-11 21:01:00|80.669414401537693|2|3338353030|46|35.309074979060284|0|19|523|-80.737839|64|35.297134|FRESH POTATOES|0.0|4|RUSSET POTATO 8LB BAG|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|35.305725790410776|00033383530307|FRESH PRODUCE|PRODUCE|-80.66939|80.669395283861164|258|1
35.28326|2e72fa87af49333858d9e7585dc460c2130bfb12|12.99|2015-02-27 12:33:00|80.669414401537693|2|3125903266|46|35.309074979060284|0|19|9937|-80.737839|885|35.297134|NFS POP SAUV/FUME BLANC|0.0|13|YELLOW TAIL SAUV BLANC 1.5L|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|35.305725790410776|00031259032665|POPULAR (4-$7.99)|WINE|-80.66939|80.669395283861164|258|1
35.28326|684fa712264ced8812a390c45cce8762295d46f6|9.99|2014-09-28 12:02:00|80.669414401537693|2|8992427896|46|35.309074955099199|0|19|455|-80.662946|82|35.412407|DOMESTIC PREMIUM 12PK&>|0.0|16|YUENGLING LAGER 12PK 12OZ BTL|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|35.305725790410776|00089924278962|DOMESTIC BEER|BEER|-80.66939|80.669433417044175|68|1
35.28326|883accbbd50735e9fa2774732c3876368f83ee00|1.19|2015-02-22 15:45:00|80.669414401537693|2|7203653022|46|35.309074955099199|0|19|1273|-80.662946|50|35.412407|BAG VEG NON STEAM|0.0|5|HT CUT  GREEN BEANS|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|35.305725790410776|00072036530325|VEGETABLES-FROZEN|FROZEN|-80.66939|80.669433417044175|68|1
35.28326|b64e8568e788347675ab743e445fe2e181a185b2|5.83|2014-10-05 20:05:00|1.4094857484078087|2|20165500000|46|0.6158090578372145|0|26|297|-80.66939|49|35.28326|GROUND BEEF|0.0|2|HT PREMIUM GRND BEEF 80% LEAN|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00201655000005|BEEF|MEAT|-80.66939|1.4079464610753885|46|1
35.28326|f0915370c7b1b5bd740291e440aab3049b12c92a|13.98|2015-01-17 16:54:00|1.4094857484078087|2|7261345083|46|0.6158090578372145|0|26|389|-80.66939|66|35.28326|NFS-LAUNDRY DETERGENTS|2.0|1|WISK HE|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00072613450848|DETERGENTS|G1 GROCERY|-80.66939|1.4079464610753885|46|2
35.28326|ae7f6a61c90d88849ebaf013521c809dd86c5719|11.99|2015-01-03 17:11:00|80.669414401537693|2|8769200105|46|35.309074955099199|0|19|458|-80.662946|82|35.412407|CRAFT BEER|0.0|16|SAM ADAMS BOSTON LAGER 12PK|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|35.305725790410776|00087692001058|DOMESTIC BEER|BEER|-80.66939|80.669433417044175|68|1
35.28326|cd35bc25705b362f17e69d9c6117d36032659a16|1.0|2015-01-02 19:32:00|1.4094857484078087|2|3400000031|46|0.6158090578372145|0|26|47|-80.66939|7|35.28326|REGISTER BARS|0.0|1|HERSHEY KIT KAT BAR|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|0.61471665291522548|00034000002467|CANDY|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|89c2f795275dee10aa390239d410f2d0f695dd54|2.0|2015-02-27 12:38:00|80.669414401537693|2|2840000210|46|35.309074979060284|0|19|204|-80.737839|31|35.297134|TORTILLA CHIPS|0.0|1|SANTITAS WHITE CORN|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|35.305725790410776|00028400002103|SNACKS|G1 GROCERY|-80.66939|80.669395283861164|258|1
35.28326|f4f558c2a00af7782457416a503b5b36215cdbe7|9.75|2015-02-09 15:58:00|80.669414401537693|2|7203656080|46|35.309074979060284|0|19|318|-80.737839|52|35.297134|SHREDDED/GRATED CHEESE|0.0|3|HT FANCY SHRED SHARP CHED CHE|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|35.305725790410776|00072036550262|CHEESE|DAIRY|-80.66939|80.669395283861164|258|3
35.28326|9b58c43952127b3cc356be653e66500699fab1ee|7.99|2015-01-18 14:32:00|80.669414401537693|2|3410049805|46|35.309074955099199|0|19|458|-80.662946|82|35.412407|CRAFT BEER|0.0|16|LEINENKUGEL'S SUNSET WHEAT 6PK|de4b1fb5f316be64bd4aacd5f3dc1a1594bd7e6a|1.7837527370134665|35.305725790410776|00034100498054|DOMESTIC BEER|BEER|-80.66939|80.669433417044175|68|1
35.195689|877064a07d9052de005b4b0afe0aaaec402085aa|19.8|2015-03-03 16:12:00|1.4094857484078087|1|20165700000|412|0.6142806555579505|0|26|297|-80.826724|49|35.195689|GROUND BEEF|2.2|2|HT GROUND BEEF CHUCK 80% LEAN|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00201657000003|BEEF|MEAT|-80.826724|1.4106924574007214|412|3
35.195689|084b17df81bedc0dda6ab91f68d802f34e414772|26.86|2014-12-23 15:36:00|80.828402574597021|1|20228000000|412|35.211064415175038|0|8|299|-80.80146|49|35.17739|ANGUS BEEF|0.0|2|ANGUS BEEF BONELESS RUMP ROAST|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00202280000002|BEEF|MEAT|-80.826724|80.826725428806512|208|1
35.195689|01cf9008bf2a22a6a79f2c167c49ae01fb6980b6|10.64|2014-09-15 17:23:00|1.4094857484078087|1|20165700000|412|0.6142806555579505|0|26|297|-80.826724|49|35.195689|GROUND BEEF|1.18|2|HT GROUND BEEF CHUCK 80% LEAN|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00201657000003|BEEF|MEAT|-80.826724|1.4106924574007214|412|2
35.195689|e7f000af8f423c41dd0bc6410dbd6315be7b5dc6|22.96|2014-11-22 16:39:00|80.828402574597021|1|20003200000|412|35.211064413731144|0|8|974|-80.825175|201|35.152722|FRESH TURKEY|4.61|2|BUTTERBALL FRSH LT'L TURKEY|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00200032000003|POULTRY|MEAT|-80.826724|80.826732279057438|160|1
35.195689|e06e3d5003ceef093ba7eae40551aeb1b1e6ca02|13.510000000000002|2015-01-22 19:10:00|1.4094857484078087|1|20165700000|412|0.6142806555579505|0|26|297|-80.826724|49|35.195689|GROUND BEEF|1.5|2|HT GROUND BEEF CHUCK 80% LEAN|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00201657000003|BEEF|MEAT|-80.826724|1.4106924574007214|412|2
35.195689|fc913ad57ed0c56d33bcf7a59aed83d136627da4|13.07|2015-03-09 17:11:00|1.4094857484078087|1|20165700000|412|0.6142806555579505|0|26|297|-80.826724|49|35.195689|GROUND BEEF|0.98|2|HT GROUND BEEF CHUCK 80% LEAN|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00201657000003|BEEF|MEAT|-80.826724|1.4106924574007214|412|3
35.195689|b747830c67bc6462814821c9bf583795d7f3f92b|5.7|2014-12-19 16:04:00|1.4094857484078087|1|20165700000|412|0.6142806555579505|0|26|297|-80.826724|49|35.195689|GROUND BEEF|0.63|2|HT GROUND BEEF CHUCK 80% LEAN|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00201657000003|BEEF|MEAT|-80.826724|1.4106924574007214|412|1
35.195689|0988ae9140267d0474eac398addf345d1acad6e5|4.48|2014-09-20 15:38:00|80.828402574597021|1||412|35.211064413731144|0|8|501|-80.825175|64|35.152722|FRESH PEARS|0.45|4|BARTLETT PEARS|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00204409000009|FRESH PRODUCE|PRODUCE|-80.826724|80.826732279057438|160|1
35.195689|ee4fc1ef0521dacae4c522005043aa6c86a696b5|10.01|2014-10-18 15:56:00|80.828402574597021|1|20165700000|412|35.211064413731144|0|8|297|-80.825175|49|35.152722|GROUND BEEF|1.15|2|HT GROUND BEEF CHUCK 80% LEAN|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00201657000003|BEEF|MEAT|-80.826724|80.826732279057438|160|2
35.195689|b54477a64ee3c9e4c860b45878916f06beaaaec4|1.2|2015-03-03 16:53:00|1.4094857484078087|1|3663202717|412|0.6142806555579505|0|26|685|-80.826724|61|35.195689|GREEK|0.2|3|DANNON OIKOS TOASTED COCONUT|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00036632027276|YOGURT|DAIRY|-80.826724|1.4106924574007214|412|1
35.195689|55ab76c4ecb0cead65ad74a17424d700cb915db8|6.25|2014-09-25 16:13:00|1.4094857484078087|1|2400016286|412|0.6142806555579505|0|26|245|-80.826724|39|35.195689|VEGETABLES-CORE|0.0|1|DEL MONTE CRISP CORN|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00024000015444|VEGETABLES-CAN/JAR|G1 GROCERY|-80.826724|1.4106924574007214|412|5
35.195689|4f5526ed0fa83b586056ab2d0ffb3b63d40de1b3|3.79|2015-02-24 12:36:00|1.4094857484078087|1|2100062503|412|0.6142806555579505|0|26|318|-80.826724|52|35.195689|SHREDDED/GRATED CHEESE|1.29|3|KRAFT SHREDDED FIVE CHEESE|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00021000607082|CHEESE|DAIRY|-80.826724|1.4106924574007214|412|1
35.195689|92a58dd08d4db984cf53d2837d87dc7df1c176e8|4.99|2015-02-14 15:29:00|80.828402574597021|1|2410044068|412|35.211064413731144|0|8|87|-80.825175|13|35.152722|CHEESE CRACKERS|1.49|1|CHEEZ-IT PEPPERJACK|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00024100789252|CRACKERS|G1 GROCERY|-80.826724|80.826732279057438|160|1
35.195689|008f24dd9fb764ee3c6ea7afd4b85c79aa4e0ef9|4.29|2014-12-30 14:05:00|80.828402574597021|1|2840016014|412|35.211064415175038|0|8|201|-80.80146|31|35.17739|POTATO CHIPS|0.29|1|LAYS WAVY REGULAR|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00028400160209|SNACKS|G1 GROCERY|-80.826724|80.826725428806512|208|1
35.195689|e6467163d713ffab15210351830b5970148a294d|7.58|2015-01-13 12:02:00|80.828402574597021|1|2100062503|412|35.211064413731144|0|8|318|-80.825175|52|35.152722|SHREDDED/GRATED CHEESE|2.58|3|KRAFT SHREDDED FIVE CHEESE|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00021000607082|CHEESE|DAIRY|-80.826724|80.826732279057438|160|2
35.195689|8bd14e38c3252ed9f52aa65ff988cf5a84044ec0|3.49|2015-03-05 11:20:00|80.828402574597021|1|2840008294|412|35.211064413731144|0|8|201|-80.825175|31|35.152722|POTATO CHIPS|0.49|1|LAYS KETTLE REGULAR|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00028400082945|SNACKS|G1 GROCERY|-80.826724|80.826732279057438|160|1
35.195689|8d3ae419cab72942cb78616f15810de01d8998b6|3.49|2015-01-16 09:02:00|1.4094857484078087|1|2840008294|412|0.6142806555579505|0|26|201|-80.826724|31|35.195689|POTATO CHIPS|0.99|1|LAYS KETTLE REGULAR|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00028400082945|SNACKS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|38836361eec0a34426b3d2109997659fedaf4059|3.49|2014-12-12 12:53:00|1.4094857484078087|1|2840008294|412|0.6142806555579505|0|26|201|-80.826724|31|35.195689|POTATO CHIPS|0.99|1|LAYS KETTLE REGULAR|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00028400082945|SNACKS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|79bb732fef0ea589535517ea2cf3c1b606e2d2ae|3.69|2014-11-28 12:41:00|1.4094857484078087|1|2100062503|412|0.6142806555579505|0|26|318|-80.826724|52|35.195689|SHREDDED/GRATED CHEESE|0.69|3|KRAFT SHREDDED FIVE CHEESE|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00021000607082|CHEESE|DAIRY|-80.826724|1.4106924574007214|412|1
35.195689|45a7a2f7bf73f4ad2873f8ddb3abdf36bf75c6d2|6.25|2014-11-13 16:21:00|80.828402574597021|1|2400016286|412|35.211064413731144|0|8|245|-80.825175|39|35.152722|VEGETABLES-CORE|1.25|1|DEL MONTE CRISP CORN|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00024000015444|VEGETABLES-CAN/JAR|G1 GROCERY|-80.826724|80.826732279057438|160|5
35.195689|89e670bf4095605e569e8e821486edb6379b47b2|2.5|2014-10-07 12:48:00|80.828402574597021|1|2400016286|412|35.211064413731144|0|8|245|-80.825175|39|35.152722|VEGETABLES-CORE|0.0|1|DEL MONTE CRISP CORN|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00024000015444|VEGETABLES-CAN/JAR|G1 GROCERY|-80.826724|80.826732279057438|160|2
35.195689|f59005a8052737b9d3fe24dfd8a4ddee511f2788|5.0|2015-01-31 19:07:00|80.828402574597021|1|2400016286|412|35.211064413731144|0|8|245|-80.825175|39|35.152722|VEGETABLES-CORE|0.0|1|DEL MONTE CRISP CORN|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00024000015444|VEGETABLES-CAN/JAR|G1 GROCERY|-80.826724|80.826732279057438|160|4
35.195689|7bf2aa33e157cb5747eeb148d591d57db092ccf5|3.79|2015-02-19 17:06:00|1.4094857484078087|1|2100062503|412|0.6142806555579505|0|26|318|-80.826724|52|35.195689|SHREDDED/GRATED CHEESE|1.29|3|KRAFT SHREDDED FIVE CHEESE|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00021000607082|CHEESE|DAIRY|-80.826724|1.4106924574007214|412|1
35.195689|62badfaf2e09fd1a31c55b7580e74d12e216d65c|3.49|2015-01-24 14:18:00|1.4094857484078087|1|2840008294|412|0.6142806555579505|0|26|201|-80.826724|31|35.195689|POTATO CHIPS|0.99|1|LAYS KETTLE REGULAR|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00028400082945|SNACKS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|2a802a7c48b266b428f417648b7e193a735352a7|3.99|2014-11-15 13:25:00|80.828402574597021|1|79830413741|412|35.211064413731144|0|8|756|-80.825175|87|35.152722|NFS-FLORAL ACCESSORIES|0.0|9|GRETEA VOTIVE|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00798304137415|FLORAL|FLORAL|-80.826724|80.826732279057438|160|1
35.195689|1857cfc86c0f0dc5aca0f6b37c2defd3dcc87abb|6.19|2014-09-13 15:51:00|80.828402574597021|1|81075701030|412|35.211064413731144|0|8|26|-80.825175|271|35.152722|GLUTEN FREE|0.8|1|SCHAR GF CIABATTA PARBKD ROLLS|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00810757010210|GLUTEN FREE|G1 GROCERY|-80.826724|80.826732279057438|160|1
35.195689|8eee26ee9a1b88b96b152170d3b51ab8671b3ed6|39.96|2014-12-20 13:50:00|80.828402574597021|1|87293200629|412|35.211064413731144|0|8|6204|-80.825175|1548|35.152722|HIGH END|0.0|18|ARM&HAMMER AIR FILTER 12X12X1|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00872932006302|FURNACE FILTERS|GM|-80.826724|80.826732279057438|160|4
35.195689|78792056674dc8191355234d4391ea1de31d6dec|9.99|2014-11-01 13:29:00|80.828402574597021|1|81409101202|412|35.211064413731144|0|8|6911|-80.825175|1582|35.152722|DOG TOYS|0.0|18|R&W STUFFERZ|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00814091012022|PET NEEDS|GM|-80.826724|80.826732279057438|160|1
35.195689|feb5ad34a3775470d9c9945626945149b6b85c3b|4.19|2014-10-19 15:40:00|80.828402574597021|1|30521500700|412|35.211064413731144|0|8|4834|-80.825175|1235|35.152722|COTTON/SWABS|0.0|17|Q-TIPS VALUE PACK-00700|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00305215007005|FIRST AID|HBC|-80.826724|80.826732279057438|160|1
35.195689|458f2d066c295cd93350adf492c46e5a3df9983c|7.65|2015-01-13 12:59:00|1.4094857484078087|1|76211120604|412|0.6142806555579505|0|26|36|-80.826724|10|35.195689|PREMIUM GROUND|0.66|1|STARBUCKS BRKF BLND GRND COFFE|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00762111206251|COFFEE|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|74a23f05bdbb0f7f9cea5a8245404aa08b782a53|9.75|2014-12-16 16:26:00|80.828402574597021|1|36382427864|412|35.211064413731144|0|8|4236|-80.825175|1200|35.152722|DEX ADULT/CHILDREN|0.0|17|MUCINEX CHLD CLD,COUG,THRT BRY|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00363824278643|COUGH/COLD/SINUS|HBC|-80.826724|80.826732279057438|160|1
35.195689|457bd9fb23f9f68c62057ebd2b80e555da17a9b7|4.49|2014-09-18 16:03:00|80.828402574597021|1|74759930652|412|35.211064413731144|0|8|62|-80.825175|7|35.152722|SPECIALTY BAR/BOX CHOCOLATE|0.5|1|GHIR DRK CHOC CARAMEL SEASALT|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00747599303142|CANDY|G1 GROCERY|-80.826724|80.826732279057438|160|1
35.195689|ab78156624afe8a87db544827a0c175e9a846746|4.99|2014-10-12 14:47:00|80.828402574597021|1|30997611100|412|35.211064415175038|0|8|3097|-80.80146|1000|35.17739|IMPLEMENTS NAIL-REVLON|0.0|17|REV ADV DESIGN EYELASH CURLER|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00309976111001|COSMETICS|HBC|-80.826724|80.826725428806512|208|1
35.195689|1969506d68112e1b56a64f04100c3f90293f4a64|4.49|2015-02-16 15:58:00|1.4094857484078087|1|74759930652|412|0.6142806555579505|0|26|62|-80.826724|7|35.195689|SPECIALTY BAR/BOX CHOCOLATE|0.99|1|GHIR DRK CHOC CARAMEL SEASALT|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00747599303142|CANDY|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|473feccc4e4c59cd24cd1c0b153b8ca65a4eb179|2.35|2014-12-27 12:57:00|80.828402574597021|1|2150004209|412|35.211064413731144|0|8|71|-80.825175|11|35.152722|GROC CONDIMENTS MARINADE|0.0|1|LAWRYS MARINADE STEAK & CHOP|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00021500042178|CONDIMENTS|G1 GROCERY|-80.826724|80.826732279057438|160|1
35.195689|817020b5ce87dc8b317dc900b51c663bfeca06da|8.38|2014-10-14 13:17:00|1.4094857484078087|1|2100062503|412|0.6142806555579505|0|26|318|-80.826724|52|35.195689|SHREDDED/GRATED CHEESE|3.38|3|KRAFT FINELY SHREDDED SHARP C|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00021000638741|CHEESE|DAIRY|-80.826724|1.4106924574007214|412|2
35.195689|7847b0c293045bec5148b26db396e154e0b3c14d|3.79|2015-02-02 17:06:00|1.4094857484078087|1|2100062503|412|0.6142806555579505|0|26|318|-80.826724|52|35.195689|SHREDDED/GRATED CHEESE|1.9|3|KRAFT MEXICAN FOUR CHEESE SHR|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00021000638994|CHEESE|DAIRY|-80.826724|1.4106924574007214|412|1
35.195689|d765772da2fbb6965b106442da448d0583059933|2.4|2015-02-26 17:58:00|1.4094857484078087|1|3663202717|412|0.6142806555579505|0|26|685|-80.826724|61|35.195689|GREEK|0.4|3|DANNON OIKOS STRAWBERRY TRAD|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00036632032188|YOGURT|DAIRY|-80.826724|1.4106924574007214|412|2
35.195689|10f3215356e60187c9c3467bc4f8923b8131a70d|3.89|2014-10-06 17:21:00|1.4094857484078087|1|3800039118|412|0.6142806555579505|0|26|81|-80.826724|9|35.195689|RTE CEREAL KIDS|1.9|1|KELLOGG CORN POPS 12.5|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00038000391095|CEREAL|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|21cf523903ee9541718d418b9587b3d0c9617423|2.15|2015-02-08 17:20:00|1.4094857484078087|1|3800030110|412|0.6142806555579505|0|26|44|-80.826724|6|35.195689|TOASTER PASTRIES-SHELF STABLE|0.48|1|KELL POPTART UF BLUEBERRY|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00038000300103|BREAKFAST FOODS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|83e791a514a7c1f75a11e26c46997b6a8efc180e|3.49|2015-01-03 15:32:00|1.4094857484078087|1|3800039118|412|0.6142806555579505|0|26|81|-80.826724|9|35.195689|RTE CEREAL KIDS|0.0|1|KELLOGG CORN POPS 12.5|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00038000391095|CEREAL|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|e6ce33cb450f77074494a5f6eaa3d22127a432a8|4.49|2014-10-11 10:22:00|1.4094857484078087|1|2150000300|412|0.6142806555579505|0|26|221|-80.826724|34|35.195689|SALT SALT SUBSTITUTES|0.0|1|LAWRY'S SEASONED SALT|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00021500003001|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|9d445ddd67a79576635447daaccb803b8d2edf52|2.79|2015-01-19 15:27:00|1.4094857484078087|1|7225001130|412|0.6142806555579505|0|26|1033|-80.826724|163|35.195689|HAMBURGER|0.0|7|MERITA 8PK HAMBURGER BUNS|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00072250011303|BUNS/ROLLS|COMMERCIAL BAKERY|-80.826724|1.4106924574007214|412|1
35.195689|86ed19d4870b3e3d34b9750f132612f42cb6f12e|2.79|2015-02-08 14:32:00|1.4094857484078087|1|7225001130|412|0.6142806555579505|0|26|1033|-80.826724|163|35.195689|HAMBURGER|0.0|7|MERITA 8PK HAMBURGER BUNS|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00072250011303|BUNS/ROLLS|COMMERCIAL BAKERY|-80.826724|1.4106924574007214|412|1
35.195689|fc5cfefb5bcf3aa580bf1a5230b61d71d92de727|5.58|2015-01-09 10:42:00|1.4094857484078087|1|7225001130|412|0.6142806555579505|0|26|1033|-80.826724|163|35.195689|HAMBURGER|0.0|7|MERITA 8PK HAMBURGER BUNS|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00072250011303|BUNS/ROLLS|COMMERCIAL BAKERY|-80.826724|1.4106924574007214|412|2
35.195689|1e5bf6dde755a379c3e22494d885b448a84954b5|2.79|2015-01-15 17:55:00|80.828402574597021|1|7225001130|412|35.211064415175038|0|8|1033|-80.80146|163|35.17739|HAMBURGER|0.0|7|MERITA 8PK HAMBURGER BUNS|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00072250011303|BUNS/ROLLS|COMMERCIAL BAKERY|-80.826724|80.826725428806512|208|1
35.195689|a3f254d625b0987c4efe3043e2789b6e05374905|8.45|2014-10-23 10:59:00|80.828402574597021|1|7680828008|412|35.211064413731144|0|8|149|-80.825175|23|35.152722|WHSE PASTA CORE|0.0|1|BARILLA PASTA ANGEL HAIR|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00076808501063|PASTA|G1 GROCERY|-80.826724|80.826732279057438|160|5
35.195689|df00970637d46147e341215b24751f7408720164|4.99|2014-12-15 08:16:00|80.828402574597021|1|70210104593|412|35.211064415175038|0|8|29|-80.80146|3|35.17739|REMAINING BAKING SUPPLIES|0.7|1|I/O PENNANT RED CHERRIES|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00702101045132|BAKING SUPPLIES|G1 GROCERY|-80.826724|80.826725428806512|208|1
35.195689|7addc06dd815ea391c02fbbab513179c2559787f|19.99|2015-02-06 17:21:00|1.4094857484078087|1|72760006115|412|0.6142806555579505|0|26|1509|-80.826724|87|35.195689|FLOR-FLORAL-CANDY ARANGEMENT|0.0|9|SQUARE CHOCOLATE  SCV03GEN|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00727600061155|FLORAL|FLORAL|-80.826724|1.4106924574007214|412|1
35.195689|92ac3d3e6d3899e32c639eb45670f0f9cd0c1386|8.58|2014-12-06 13:48:00|1.4094857484078087|1|1090000015|412|0.6142806555579505|0|26|440|-80.826724|76|35.195689|NFS-ALUMINUM FOIL|2.58|1|REYNOLDS FOIL 75 FT|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00010900000154|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.826724|1.4106924574007214|412|2
35.195689|080a190aacef9f409b4cdf26ff6816e93a93eca1|4.69|2015-02-10 16:24:00|1.4094857484078087|1|81829001282|412|0.6142806555579505|0|26|685|-80.826724|61|35.195689|GREEK|1.19|3|CHOBANI COCONUT BLEND 2% 4PK|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00818290012777|YOGURT|DAIRY|-80.826724|1.4106924574007214|412|1
35.195689|9c1dc2da1f564d3ff841c5938c5c5e0de503ed9e|3.49|2014-10-01 16:50:00|80.828402574597021|1|7172000798|412|35.211064414469782|0|8|727|-80.85013|7|35.175855|SEASONAL CANDY-SINGLE FAC|0.5|1|I/O(H14)TOOTSIE CARML APPL POP|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00071720007983|CANDY|G1 GROCERY|-80.826724|80.826729875673564|218|1
35.195689|29cb1cf2ce1c7b551e9fa2acd004d3caf233053d|3.95|2015-02-22 15:33:00|1.4094857484078087|1||412|0.6142806555579505|0|26|507|-80.826724|64|35.195689|FRESH ORANGES|0.0|4|NAVEL ORANGE, LRG|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00233107000004|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|5
35.195689|aa24d980eb2fc8e8c0fcdfb2ebb495660627b29b|4.74|2015-03-01 12:55:00|1.4094857484078087|1||412|0.6142806555579505|0|26|507|-80.826724|64|35.195689|FRESH ORANGES|0.0|4|NAVEL ORANGE, LRG|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00233107000004|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|6
35.195689|153d9d0d7ef17974d9ca92ec8edd31d4ea62609c|3.49|2014-10-22 16:43:00|1.4094857484078087|1|65724334603|412|0.6142806555579505|0|26|273|-80.826724|43|35.195689|PREMIUM NOVELTIES|0.0|5|PHILLY SWIRL SORBET CUPS|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00657243046069|FROZEN NOVELTIES|FROZEN|-80.826724|1.4106924574007214|412|1
35.195689|a67346c618a628f714fbf2b5ee21ac591442fac2|4.45|2015-01-18 15:31:00|1.4094857484078087|1||412|0.6142806555579505|0|26|507|-80.826724|64|35.195689|FRESH ORANGES|0.29|4|NAVEL ORANGE, LRG|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00233107000004|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|5
35.195689|e75045a82bc04b45616d4a8b3149c9ff2795c0cd|3.95|2015-02-18 15:19:00|1.4094857484078087|1||412|0.6142806555579505|0|26|507|-80.826724|64|35.195689|FRESH ORANGES|0.0|4|NAVEL ORANGE, LRG|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00233107000004|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|5
35.195689|54bb53eacf456ef1171ad6a4e7ff1d8ba4b215d1|2.37|2015-03-08 12:20:00|80.828402574597021|1||412|35.211064413731144|0|8|507|-80.825175|64|35.152722|FRESH ORANGES|0.19|4|NAVEL ORANGE, LRG|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00233107000004|FRESH PRODUCE|PRODUCE|-80.826724|80.826732279057438|160|3
35.195689|99a6cccf5f35bec9f284fe591dd361f10ce9af0b|3.16|2015-02-27 16:17:00|1.4094857484078087|1||412|0.6142806555579505|0|26|507|-80.826724|64|35.195689|FRESH ORANGES|0.0|4|NAVEL ORANGE, LRG|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00233107000004|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|4
35.195689|e757caa0f469f96e53c8e6a9d7b208394ea3e067|3.16|2015-02-25 15:56:00|1.4094857484078087|1||412|0.6142806555579505|0|26|507|-80.826724|64|35.195689|FRESH ORANGES|0.0|4|NAVEL ORANGE, LRG|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00233107000004|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|4
35.195689|a8690535c18d09d0167a3203b22c68e3a4920ddf|5.53|2015-03-02 16:04:00|1.4094857484078087|1||412|0.6142806555579505|0|26|507|-80.826724|64|35.195689|FRESH ORANGES|0.0|4|NAVEL ORANGE, LRG|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00233107000004|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|7
35.195689|767408514222e21824ac83dc4a5ca8fba95a98cb|2.37|2015-03-07 17:14:00|1.4094857484078087|1||412|0.6142806555579505|0|26|507|-80.826724|64|35.195689|FRESH ORANGES|0.19|4|NAVEL ORANGE, LRG|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00233107000004|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|3
35.195689|b4a8fedf11bd2d3eec1ceed9a659acdcf7f7b966|4.74|2015-03-06 15:15:00|80.828402574597021|1||412|35.211064413731144|0|8|507|-80.825175|64|35.152722|FRESH ORANGES|0.19|4|NAVEL ORANGE, LRG|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00233107000004|FRESH PRODUCE|PRODUCE|-80.826724|80.826732279057438|160|6
35.195689|ff8014dd289c21849db62d4a0425a8bf0c3ea34c|3.49|2014-09-24 15:05:00|80.828402574597021|1|65724334603|412|35.211064415175038|0|8|273|-80.80146|43|35.17739|PREMIUM NOVELTIES|0.0|5|PHILLY SWIRL SORBET CUPS|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00657243046069|FROZEN NOVELTIES|FROZEN|-80.826724|80.826725428806512|208|1
35.195689|b0671c3a33d4ce0e1f114e9118774b6dee0bb28c|2.95|2014-11-06 11:32:00|80.828402574597021|1|76172005110|412|35.211064413731144|0|8|25|-80.825175|3|35.152722|BAKING SYRUPS|0.45|1|KARO DARK CORN SYRUP|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00761720050101|BAKING SUPPLIES|G1 GROCERY|-80.826724|80.826732279057438|160|1
35.195689|01ec3ceb917ff65cbec3b4d673980c06a42eebd2|3.38|2014-10-05 13:13:00|80.828402574597021|1|7203688003|412|35.211064413731144|0|8|527|-80.825175|64|35.152722|FRESH CARROTS|0.38|4|HT BABY CARROTS 1LB BAG|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00072036880031|FRESH PRODUCE|PRODUCE|-80.826724|80.826732279057438|160|2
35.195689|0e77b496d29b1372f33f787dab44cafdb9e523fc|3.38|2014-11-03 15:14:00|80.828402574597021|1|7203688003|412|35.211064413731144|0|8|527|-80.825175|64|35.152722|FRESH CARROTS|0.38|4|HT BABY CARROTS 1LB BAG|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00072036880031|FRESH PRODUCE|PRODUCE|-80.826724|80.826732279057438|160|2
35.195689|be0e3628592f6a43be63754ed00a3fb8d2c49f8b|3.38|2014-11-09 13:04:00|80.828402574597021|1|7203688003|412|35.211064413731144|0|8|527|-80.825175|64|35.152722|FRESH CARROTS|0.38|4|HT BABY CARROTS 1LB BAG|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00072036880031|FRESH PRODUCE|PRODUCE|-80.826724|80.826732279057438|160|2
35.195689|fa272b76c90f485756010613e806ab6bc0f184dc|3.38|2014-10-30 12:02:00|80.828402574597021|1|7203688003|412|35.211064413731144|0|8|527|-80.825175|64|35.152722|FRESH CARROTS|0.38|4|HT BABY CARROTS 1LB BAG|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00072036880031|FRESH PRODUCE|PRODUCE|-80.826724|80.826732279057438|160|2
35.195689|a648e06bd604ce5618bda217ee77a816ed244b52|3.38|2015-01-11 14:43:00|80.828402574597021|1|7203688003|412|35.211064413731144|0|8|527|-80.825175|64|35.152722|FRESH CARROTS|0.38|4|HT BABY CARROTS 1LB BAG|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00072036880031|FRESH PRODUCE|PRODUCE|-80.826724|80.826732279057438|160|2
35.195689|d07d08211ecd519f9c48ea31b088d765435df4d2|2.59|2014-11-06 19:23:00|1.4094857484078087|1|7203663996|412|0.6142806555579505|0|26|342|-80.826724|57|35.195689|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00072036631299|MILK|DAIRY|-80.826724|1.4106924574007214|412|1
35.195689|6f1a1bc31a0fc4500977d5b0fd3e4799f8b9d094|2.99|2015-01-04 11:36:00|1.4094857484078087|1|7203663104|412|0.6142806555579505|0|26|364|-80.826724|55|35.195689|ORGANIC AND CF EGGS|0.0|3|HTN NEST GRADE A LARGE EGG BRO|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00072036631046|EGGS FRESH|DAIRY|-80.826724|1.4106924574007214|412|1
35.195689|261306f2083d8af1a3dcfd9257113bf853a4447b|2.99|2014-09-27 13:25:00|80.828402574597021|1|7203663104|412|35.211064413731144|0|8|364|-80.825175|55|35.152722|ORGANIC AND CF EGGS|0.0|3|HTN NEST GRADE A LARGE EGG BRO|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00072036631046|EGGS FRESH|DAIRY|-80.826724|80.826732279057438|160|1
35.195689|8d873d6386e339a0d8033a58cf788aa540ae6c7a|2.99|2014-12-14 17:41:00|1.4094857484078087|1|7203663104|412|0.6142806555579505|0|26|364|-80.826724|55|35.195689|ORGANIC AND CF EGGS|0.0|3|HTN NEST GRADE A LARGE EGG BRO|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00072036631046|EGGS FRESH|DAIRY|-80.826724|1.4106924574007214|412|1
35.195689|24f90824d27e98182e3887b92fcf8ca41cd33497|2.99|2015-02-04 12:19:00|80.828402574597021|1|7203663104|412|35.211064413731144|0|8|364|-80.825175|55|35.152722|ORGANIC AND CF EGGS|0.0|3|HTN NEST GRADE A LARGE EGG BRO|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00072036631046|EGGS FRESH|DAIRY|-80.826724|80.826732279057438|160|1
35.195689|a201c6016f0ae48427b3d5138c698dc098dae271|2.99|2014-09-30 15:55:00|80.828402574597021|1|7203663104|412|35.211064413731144|0|8|364|-80.825175|55|35.152722|ORGANIC AND CF EGGS|0.0|3|HTN NEST GRADE A LARGE EGG BRO|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00072036631046|EGGS FRESH|DAIRY|-80.826724|80.826732279057438|160|1
35.195689|8bfcdbb8625aa1702c2f809593b032393f03b47f|2.99|2014-09-12 12:57:00|80.828402574597021|1|7203663104|412|35.211064414469782|0|8|364|-80.85013|55|35.175855|ORGANIC AND CF EGGS|0.0|3|HTN NEST GRADE A LARGE EGG BRO|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00072036631046|EGGS FRESH|DAIRY|-80.826724|80.826729875673564|218|1
35.195689|9acbda8b103d5088fba884ad97387f0c91148cac|11.83|2015-02-28 12:53:00|1.4094857484078087|1|20196000000|412|0.6142806555579505|0|26|299|-80.826724|49|35.195689|ANGUS BEEF|1.48|2|ANGUS BF FLAT IRON STK CUSTOM|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00201960000004|BEEF|MEAT|-80.826724|1.4106924574007214|412|1
35.195689|75f48f64eddaee77341c291502ba2f5b5b239398|6.98|2014-11-23 16:03:00|80.828402574597021|1|20455000000|412|35.211064413731144|0|8|542|-80.825175|64|35.152722|FRESH VEGETABLES REMAIN|0.98|4|BRUSSEL SPROUTS 1LB (RPC)|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00094922577160|FRESH PRODUCE|PRODUCE|-80.826724|80.826732279057438|160|2
35.195689|e96753de0540dc1d4219f20c1e25c8fffdcfb9b4|46.36|2014-12-05 13:12:00|1.4094857484078087|1|20324300000|412|0.6142806555579505|0|26|641|-80.826724|137|35.195689|PREMIUM PORK|11.39|2|PORK BABY BACK RIBS|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00203243000008|PORK|MEAT|-80.826724|1.4106924574007214|412|2
35.195689|92cdacaab2ab90bd6a780c22200f329135f5813d|3.09|2014-12-31 14:38:00|1.4094857484078087|1|20394300000|412|0.6142806555579505|0|26|643|-80.826724|137|35.195689|PORK OFFALS-FROZEN|0.25|2|MORTY PRIDE SMOKED HOCKS|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00203943000001|PORK|MEAT|-80.826724|1.4106924574007214|412|1
35.195689|ebd40d2d0a6314c60394b236c84b259f5e1b597f|10.47|2014-11-25 15:44:00|80.828402574597021|1|20455000000|412|35.211064413731144|0|8|542|-80.825175|64|35.152722|FRESH VEGETABLES REMAIN|1.47|4|BRUSSEL SPROUTS 1LB (RPC)|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00094922577160|FRESH PRODUCE|PRODUCE|-80.826724|80.826732279057438|160|3
35.195689|434a408427193282b338708f7dc1b1c002a70500|2.99|2014-11-13 18:52:00|1.4094857484078087|1|8201110007|412|0.6142806555579505|0|26|1250|-80.826724|12|35.195689|SPECIALTY COOKIES|0.99|1|MURRAY GINGER SNAPS|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00082011100078|COOKIES|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|31fb585d82e7c881c1dd90f0bc7cb4517117f6e1|3.19|2014-09-22 16:12:00|80.828402574597021|1|7641090137|412|35.211064415175038|0|8|1255|-80.80146|13|35.17739|LUNCH BOX CRACKERS|0.0|1|LANCE R/F TOASTCHEESE|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00076410523330|CRACKERS|G1 GROCERY|-80.826724|80.826725428806512|208|1
35.195689|f5ccd9eadfcd3e15c99d0f5eb9daa7fa92dfade9|2.29|2014-12-22 16:33:00|1.4094857484078087|1|7800023046|412|0.6142806555579505|0|26|55|-80.826724|8|35.195689|REGULAR|1.29|23|CHEERWINE 2 LTR NR|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00070925000300|CARBONATED BEVERAGES|BEVERAGE|-80.826724|1.4106924574007214|412|1
35.195689|dec3177b6c1173c392a90ac5a36b448ee35b7408|3.69|2014-09-14 16:38:00|80.828402574597021|1|7518500003|412|35.211064413731144|0|8|1033|-80.825175|163|35.152722|HAMBURGER|0.0|7|MARTIN'S POTATO SANDWICH ROLLS|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00075185000039|BUNS/ROLLS|COMMERCIAL BAKERY|-80.826724|80.826732279057438|160|1
35.195689|ea8328606dc90bdcd06ac6a006dff776cda6771f|6.5|2014-12-10 12:56:00|80.828402574597021|1|7203656080|412|35.211064413731144|0|8|318|-80.825175|52|35.152722|SHREDDED/GRATED CHEESE|3.25|3|HT SHRED WISC XTRA SHARP CHED|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00072036705181|CHEESE|DAIRY|-80.826724|80.826732279057438|160|2
35.195689|1f50d850e599db3a6583ae3474da01f720eb595e|7.99|2015-02-05 17:17:00|80.828402574597021|1|7940033944|412|35.211064413731144|0|8|3586|-80.825175|1050|35.152722|GELS|0.0|17|AXE SPIKED UP LOOK X HOLD GEL|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00079400339980|HAIR STYLING|HBC|-80.826724|80.826732279057438|160|1
35.195689|4936a2785cf4d9ea9a6ee8c890ddb0a72e703b69|2.99|2014-10-20 15:17:00|80.828402574597021|1|7482064552|412|35.211064415175038|0|8|6785|-80.80146|1568|35.17739|MAGAZINES WEEKLY|0.0|18|IN TOUCH WEEKLY|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00074820645529|MAGAZINES|GM|-80.826724|80.826725428806512|208|1
35.195689|d566ef901c7a7781d0c5bbb4ea19a0e6bdab2fba|8.36|2014-10-16 13:17:00|1.4094857484078087|1|20242200000|412|0.6142806555579505|0|26|299|-80.826724|49|35.195689|ANGUS BEEF|0.0|2|ANGUS BEEF SKIRT STEAK FAJITAS|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00202422000006|BEEF|MEAT|-80.826724|1.4106924574007214|412|1
35.195689|a5493436057643de7b22bb4c326dfaeb5937b906|19.02|2015-01-07 13:00:00|80.828402574597021|1|20250700000|412|35.211064413731144|0|8|642|-80.825175|49|35.152722|NATURAL/ORGANIC BEEF|2.38|2|NATURAL 90% LEAN GRND BF CUSTM|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00202506000007|BEEF|MEAT|-80.826724|80.826732279057438|160|1
35.195689|2a768580ab847209e2dcbb9eeb2612bf2cad45a5|32.52|2014-12-02 11:34:00|80.828402574597021|1|20250700000|412|35.211064413731144|0|8|642|-80.825175|49|35.152722|NATURAL/ORGANIC BEEF|4.07|2|NATURAL 90% LEAN GRND BF CUSTM|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00202506000007|BEEF|MEAT|-80.826724|80.826732279057438|160|1
35.195689|0da5aa4beadec32545324e1bbf8292cdde458fa4|3.49|2014-09-17 09:58:00|80.828402574597021|1|7080095048|412|35.211064415175038|0|8|357|-80.80146|104|35.17739|SMOKED SAUSAGE ROPES|1.02|19|SMITHFIELD SMOKED SAUSAGE LOOP|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00070800950485|DINNER SAUSAGE|CASE READY MEATS|-80.826724|80.826725428806512|208|1
35.195689|38e6bb9a768e352eab6fc5a1b989e4bff708a28c|1.3|2014-11-05 12:55:00|80.828402574597021|1|5000042264|412|35.211064413731144|0|8|154|-80.825175|24|35.152722|NFS-CAT FOOD WET|0.3|1|FRISKIES BUFFET SLICED CHICKEN|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00050000421947|PET FOOD/SUPPLIES|G1 GROCERY|-80.826724|80.826732279057438|160|2
35.195689|1adb9836c9702fcffd39917343b9ef9489573124|7.78|2015-01-27 13:00:00|80.828402574597021|1|4610000094|412|35.211064413731144|0|8|318|-80.825175|52|35.152722|SHREDDED/GRATED CHEESE|2.78|3|SARGENTO CB FOUR STATE CHEDDAR|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00046100011065|CHEESE|DAIRY|-80.826724|80.826732279057438|160|2
35.195689|ae00c4c4a53b740e12f652f8dfd46d6a87d281b2|2.39|2014-10-30 14:27:00|1.4094857484078087|1|5210004680|412|0.6142806555579505|0|26|734|-80.826724|3|35.195689|NFS-CANDLES/BIRTHDAY SUP|0.89|1|MC DECORATING TIPS|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00052100046808|BAKING SUPPLIES|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|367bf863f128bb0a12357b8af8f3842e886a663b|3.59|2014-12-03 16:50:00|80.828402574597021|1|4850002013|412|35.211064413731144|0|8|335|-80.825175|56|35.152722|ORANGE JUICE-REGRIGERATED|0.59|3|TROPICANA PP GROVESTAND|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00048500304143|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.826724|80.826732279057438|160|1
35.195689|77df25c52d065dbb9964e44b058e1f78880c4e84|5.34|2014-12-09 15:48:00|1.4094857484078087|1|7047045916|412|0.6142806555579505|0|26|685|-80.826724|61|35.195689|GREEK|1.34|3|YOPLAIT GREEK BLEND STWBRY RAS|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00070470459158|YOGURT|DAIRY|-80.826724|1.4106924574007214|412|4
35.195689|2cc8ac53602bdae8e577f1dd77a4269f4efaa1bd|4.99|2015-01-08 14:07:00|1.4094857484078087|1|7203688080|412|0.6142806555579505|0|26|523|-80.826724|64|35.195689|FRESH POTATOES|2.5|4|HT YUKON GOLD 5 LB BAG|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00072036880802|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|1
35.195689|4fb5544820062be80a5bc434c19807645f16081a|13.29|2015-01-08 17:48:00|1.4094857484078087|1|3700013882|412|0.6142806555579505|0|26|389|-80.826724|66|35.195689|NFS-LAUNDRY DETERGENTS|0.0|1|TIDE HE W/FEBREZE SPRING|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00037000875611|DETERGENTS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|0de9d625d7508e0260273cc1a3f61a64542e4049|8.3|2015-02-15 16:35:00|1.4094857484078087|1||412|0.6142806555579505|0|26|529|-80.826724|64|35.195689|FRESH ASPARAGUS|2.08|4|GREEN  ASPARAGUS|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00204080000008|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|1
35.195689|9989882f458f85a7ccc7e075dfa4dae17fbb0142|23.14|2014-12-28 14:45:00|1.4094857484078087|1||412|0.6142806555579505|0|26|500|-80.826724|64|35.195689|FRESH APPLES|3.87|4|HONEY CRISP APPLE|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00233283000003|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|1
35.195689|6aff9b2c5e5bb1dd8a118f222852c0c75351e953|13.93|2014-10-29 15:22:00|1.4094857484078087|1||412|0.6142806555579505|0|26|500|-80.826724|64|35.195689|FRESH APPLES|5.24|4|HONEY CRISP APPLE|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00233283000003|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|1
35.195689|1f800fb72432e7a876293f2ecb7a8270789cdd58|13.54|2015-01-26 17:02:00|1.4094857484078087|1||412|0.6142806555579505|0|26|500|-80.826724|64|35.195689|FRESH APPLES|0.0|4|HONEY CRISP APPLE|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00233283000003|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|1
35.195689|011e3b3f2b0fcb5479d4cf5c6aaa30c91e962517|11.98|2015-03-04 15:21:00|80.828402574597021|1||412|35.211064415175038|0|8|500|-80.80146|64|35.17739|FRESH APPLES|0.0|4|HONEY CRISP APPLE|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00233283000003|FRESH PRODUCE|PRODUCE|-80.826724|80.826725428806512|208|1
35.195689|8f4ef6ac342f62eddd85376f6270e1c06abe5601|14.06|2015-02-24 17:13:00|1.4094857484078087|1||412|0.6142806555579505|0|26|500|-80.826724|64|35.195689|FRESH APPLES|0.0|4|HONEY CRISP APPLE|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00233283000003|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|1
35.195689|7c44152658ace6b8931b45d5ee047fa2a7b7740b|2.99|2015-01-23 11:03:00|1.4094857484078087|1|7203695360|412|0.6142806555579505|0|26|1629|-80.826724|373|35.195689|TAKE & BAKE ROLLS|0.0|14|TAKE & BAKE PETITE PN RL 6 CT|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00072036953605|ROLLS|BAKERY|-80.826724|1.4106924574007214|412|1
35.195689|ed2a4e3962b03c4b2eec1f08e90210ceae6f9bed|8.99|2014-09-23 14:17:00|80.828402574597021|1|7203688113|412|35.211064413731144|0|8|583|-80.825175|136|35.152722|NUTS|0.0|4|HT PECAN PIECES TRAY|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00072036881137|OTHER MERCHANDISE|PRODUCE|-80.826724|80.826732279057438|160|1
35.195689|952dac487f9f460c0b0a440fb15d0e0e0e5371da|5.29|2014-10-02 13:00:00|80.828402574597021|1|5209220392|412|35.211064413731144|0|8|5827|-80.825175|1536|35.152722|FOILWARE CASSEROLE|0.0|18|CNC LASAGNA PAN W/LID|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00052092203920|FOILWARE|GM|-80.826724|80.826732279057438|160|1
35.195689|fc3f99edacac5bd764a2e79085aad44ca5a3f165|24.46|2014-11-29 16:04:00|80.828402574597021|1|20899100000|412|35.211064413731144|0|8|1421|-80.825175|201|35.152722|SMART CHICKEN VEGETABLE FED|0.0|2|SMART CHICKEN BREAST TENDERS|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00208991000003|POULTRY|MEAT|-80.826724|80.826732279057438|160|2
35.195689|c1e7fd1eb301ea455c02ed59c83b398ed34bf6e3|7.5|2015-01-01 12:49:00|80.828402574597021|1|4610000094|412|35.211064413731144|0|8|333|-80.825175|52|35.152722|PARMESAN CHEESE|2.5|3|SARGENTO ARTISAN PARMESAN|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00046100000595|CHEESE|DAIRY|-80.826724|80.826732279057438|160|2
35.195689|44eaaaa921e9f173966dcf220fc7353a16f60613|3.39|2014-12-07 15:16:00|1.4094857484078087|1|4450034122|412|0.6142806555579505|0|26|357|-80.826724|104|35.195689|SMOKED SAUSAGE ROPES|0.0|19|HILLSHIRE BEEF POLSKA KIELBASA|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00044500339048|DINNER SAUSAGE|CASE READY MEATS|-80.826724|1.4106924574007214|412|1
35.195689|7d0c84ce4c255978a6d0b8f846daadeb8aa895ff|2.78|2014-11-16 14:16:00|1.4094857484078087|1|4100002278|412|0.6142806555579505|0|26|238|-80.826724|38|35.195689|RICE FLAVORED|0.0|1|KNORR RICE CHEDDAR BROCCOLI|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00041000022784|RICE GRAINS AND BEANS|G1 GROCERY|-80.826724|1.4106924574007214|412|2
35.195689|261ce28aa2038fbba8049838db8139e4bcaca32c|2.78|2014-09-10 18:02:00|1.4094857484078087|1|4100002278|412|0.6142806555579505|0|26|238|-80.826724|38|35.195689|RICE FLAVORED|0.0|1|KNORR RICE CHEDDAR BROCCOLI|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00041000022784|RICE GRAINS AND BEANS|G1 GROCERY|-80.826724|1.4106924574007214|412|2
35.195689|5488babdb7a14e5d495aaae331c1c628be37bef9|2.75|2015-02-21 13:55:00|1.4094857484078087|1|5150002325|412|0.6142806555579505|0|26|126|-80.826724|19|35.195689|PRESERVES/MARMALADE|0.0|1|SMUKCER SIMPLY FRT SDL STRWBRY|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00051500025710|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|85f684d8c40e15bb478e8ac9939f3209ab2d7a3e|1.19|2015-02-02 17:09:00|1.4094857484078087|1|3940001747|412|0.6142806555579505|0|26|242|-80.826724|39|35.195689|CANNED BEANS|0.19|1|BUSH BEAN SND BLACK|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00039400018841|VEGETABLES-CAN/JAR|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|5f56d77faaa22752b863f0590c5d4bff8254c31c|2.29|2014-11-19 16:25:00|1.4094857484078087|1|7203695175|412|0.6142806555579505|0|26|1607|-80.826724|371|35.195689|FROZEN DOUGH (BREAD)|0.0|14|FRESH LRG FRENCH BREAD|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00072036951755|BREAD|BAKERY|-80.826724|1.4106924574007214|412|1
35.195689|fe7384cfad20f08da5c46160c54b05ffb1e62a78|1.69|2015-01-31 14:10:00|80.828402574597021|1|4900000044|412|35.211064414469782|0|8|55|-80.85013|8|35.175855|REGULAR|0.0|23|CB COKE SINGLE 20 OZ.|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00049000000443|CARBONATED BEVERAGES|BEVERAGE|-80.826724|80.826729875673564|218|1
35.195689|909214c01aa509603b1339bc3cf9b148c23cdcb9|1.67|2015-01-18 16:35:00|1.4094857484078087|1|1070002152|412|0.6142806555579505|0|26|53|-80.826724|7|35.195689|THEATER BOX|0.67|1|JOLLY RANCHR GUMMIES BOX|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00010700708601|CANDY|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|91b4e5479f3169a869c7566080105c06f850b7dc|6.98|2015-02-07 12:06:00|1.4094857484078087|1|75733955555|412|0.6142806555579505|0|26|68|-80.826724|11|35.195689|BARBECUE SAUCES|1.02|1|STICKY FNGR BBQ SC MEMPHIS.|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00757339222220|CONDIMENTS|G1 GROCERY|-80.826724|1.4106924574007214|412|2
35.195689|e568ee618dba4b9c5134e0c01a0bdbe941edb29a|55.769999999999996|2015-02-23 13:42:00|1.4094857484078087|1|2052518367|412|0.6142806555579505|0|26|4451|-80.826724|1210|35.195689|PROBIOTICS|19.799999999999997|17|DIGEST. ADV. PROBIOTIC GUMMIES|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00020525183675|STOMACH REMEDIES|HBC|-80.826724|1.4106924574007214|412|3
35.195689|5f3fa9e6af615123955a14ca83108fc4d8775df6|18.59|2014-12-20 16:47:00|1.4094857484078087|1|2052518367|412|0.6142806555579505|0|26|4451|-80.826724|1210|35.195689|PROBIOTICS|0.0|17|DIGEST. ADV. PROBIOTIC GUMMIES|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00020525183675|STOMACH REMEDIES|HBC|-80.826724|1.4106924574007214|412|1
35.195689|35d010afb836489cfa349af8da674ae8cc7701f0|2.59|2015-02-20 17:54:00|80.828402574597021|1|2073509418|412|35.211064413731144|0|8|365|-80.825175|56|35.152722|REFRIGERATED TEAS|0.0|3|TURKEY HILL P&C SWEET TEA|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00020735094181|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.826724|80.826732279057438|160|1
35.195689|58d28432cf22ee6852187716e7f93e9ec1973848|19.99|2015-01-21 18:06:00|1.4094857484078087|1|1780013476|412|0.6142806555579505|0|26|156|-80.826724|24|35.195689|NFS-DOG FOOD-DRY|5.0|1|BENEFUL HEALTHY FIESTA|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00017800141970|PET FOOD/SUPPLIES|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|4f4a6c6f9d453fb99ce1615c0ea62564bf40e4f8|4.29|2015-01-06 14:49:00|1.4094857484078087|1|2840016014|412|0.6142806555579505|0|26|201|-80.826724|31|35.195689|POTATO CHIPS|2.14|1|LAYS SOUR CREAM & ONION|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00028400160155|SNACKS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|395a5f8f0520dc95b876a3bf2bde23aea0052397|2.99|2014-10-02 15:19:00|80.828402574597021|1|9698667013|412|35.211064415175038|0|8|3179|-80.80146|1010|35.17739|POLISH RMVR-CUTEX|0.0|17|CUTEX POLISH RMV ADV REVIVE|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00096986670139|NAIL CARE|HBC|-80.826724|80.826725428806512|208|1
35.195689|58c77319e50b005e585da2682ea8c7b41a0292d8|39.98|2015-01-20 09:13:00|1.4094857484078087|1|79500800100|412|0.6142806555579505|0|26|8092|-80.826724|1705|35.195689|PROPANE EXCHANGE|0.0|18|BLUE RHINO CYLINDER EXCHANGE|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00795008001004|PROPANE|GM|-80.826724|1.4106924574007214|412|2
35.195689|8954e072015ff0d8e37ff46c4a1ed1adacbee58f|3.58|2015-01-20 18:30:00|1.4094857484078087|1|3940001614|412|0.6142806555579505|0|26|243|-80.826724|39|35.195689|BAKED BEANS|0.0|1|BUSH BKD BEAN W/ONION 28|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00039400016038|VEGETABLES-CAN/JAR|G1 GROCERY|-80.826724|1.4106924574007214|412|2
35.195689|63a1ec6ecd48c9f904b82fa1891fe6db615c402a|1.79|2015-01-13 17:21:00|1.4094857484078087|1|3940001614|412|0.6142806555579505|0|26|243|-80.826724|39|35.195689|BAKED BEANS|0.0|1|BUSH BKD BEAN W/ONION 28|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00039400016038|VEGETABLES-CAN/JAR|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|09838ec9a0f3f8edefa2660085b64332fef3a666|5.99|2015-02-18 17:34:00|1.4094857484078087|1|3700034036|412|0.6142806555579505|0|26|388|-80.826724|66|35.195689|NFS-DISHWASH PWDR/LIQUID|0.0|1|CASCADE CLOROX DISH PWD LEMON|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00037000340416|DETERGENTS|G1 GROCERY|-80.826724|1.4106924574007214|412|1
35.195689|8ef7502c053dc39b4bb55522f50d1fa477447815|4.58|2015-01-25 17:26:00|1.4094857484078087|1|20459300000|412|0.6142806555579505|0|26|532|-80.826724|64|35.195689|FRESH CUCUMBERS|0.58|4|HOT HOUSE CUCUMBERS|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00033383671017|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|2
35.195689|acd6678dff90ea312481bd55b926619cd8c5d152|4.58|2015-02-01 14:47:00|1.4094857484078087|1||412|0.6142806555579505|0|26|532|-80.826724|64|35.195689|FRESH CUCUMBERS|0.29|4|HOT HOUSE CUCUMBERS|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00204593000007|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|2
35.195689|938e597dc2121d9e64241929a978ce80f3d869fe|0.97|2015-02-06 12:58:00|1.4094857484078087|1|7203671102|412|0.6142806555579505|0|26|1025|-80.826724|162|35.195689|WHITE|0.0|7|HT OLD FASHIONED BREAD|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00072036711021|SLICED BREAD|COMMERCIAL BAKERY|-80.826724|1.4106924574007214|412|1
35.195689|153c9dff9ad63ec7ba3c61dc53a8d1ab24769a73|3.59|2014-09-30 15:56:00|80.828402574597021|1|8265750080|412|35.211064413731144|0|8|31|-80.825175|4|35.152722|NON CARBONATED WATER|0.3|1|DEER PARK 2.5 GAL SPRING WATER|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00082657500805|BOTTLED WATER|G1 GROCERY|-80.826724|80.826732279057438|160|1
35.195689|9937cf3cd310572ed364f57c1c9f690d2e5e041e|3.49|2015-03-03 17:18:00|1.4094857484078087|1|4154030376|412|0.6142806555579505|0|26|6680|-80.826724|1564|35.195689|MECHANICAL PENCIL|0.0|18|SHARPWRITER MP .7MM YEL 30376|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00041540303763|SCHOOL & OFFICE SUPPLY|GM|-80.826724|1.4106924574007214|412|1
35.195689|71f3a2d0f27ed67bc6b1e40aecb598491a32b21d|7.75|2015-01-07 15:51:00|80.828402574597021|1|1258760034|412|35.211064413731144|0|8|443|-80.825175|76|35.152722|NFS-GARBAGE BAGS|0.0|1|GLAD TALL KIT ODOR-LEMON 13 GL|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00012587783665|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.826724|80.826732279057438|160|1
35.195689|133774dda5ad07e100e8449b9102998662e96257|2.98|2014-12-13 13:53:00|80.828402574597021|1|519|412|35.211064413731144|0|8|1896|-80.825175|450|35.152722|SODA|0.0|6|24 OZ FOUNTAIN DRINK|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|35.209978091326001|00000000005190|BEVERAGES|DELI|-80.826724|80.826732279057438|160|2
35.195689|748c3481488c6f433db1f8f971a94a4adcf6d03c|11.58|2014-10-24 16:11:00|1.4094857484078087|1|1780015014|412|0.6142806555579505|0|26|152|-80.826724|24|35.195689|NFS-CAT FOOD DRY|2.89|1|PURINA CAT CHOW|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00017800150149|PET FOOD/SUPPLIES|G1 GROCERY|-80.826724|1.4106924574007214|412|2
35.195689|d82ef14df06bc2099d31c6e3d9e2adad4c2ea858|1.79|2014-12-05 17:53:00|1.4094857484078087|1||412|0.6142806555579505|0|26|525|-80.826724|64|35.195689|FRESH LETTUCE|0.0|4|ICEBERG LETTUCE|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00204061000003|FRESH PRODUCE|PRODUCE|-80.826724|1.4106924574007214|412|1
35.195689|6f7ca8072f70ff174ce2478723d16d9b4d2445f9|6.99|2015-02-13 11:13:00|1.4094857484078087|1|3680007384|412|0.6142806555579505|0|26|4439|-80.826724|1210|35.195689|DIARRHEA REMEDY-TABLET|0.0|17|TC ANTI DIARRHEAL CAPLET 07384|de98a8036bc53a3dc31d1e9cb8c1551ac2e724c6|1.062404061359639|0.61471665291522548|00036800073845|STOMACH REMEDIES|HBC|-80.826724|1.4106924574007214|412|1
35.17335|3a6c6212ef6ce5b010482c3352d0e763e64f8b0e|2.77|2015-01-08 14:11:00|1.4094857484078087|4|3338353030|174|0.6138907664563474|0|26|523|-80.70901|64|35.17335|FRESH POTATOES|0.0|4|RUSSET POTATO 8LB BAG|e04dc890b30fd1b61727728f0d17a3f73c9aef09|1.0688318552138325|0.61471665291522548|00033383530307|FRESH PRODUCE|PRODUCE|-80.70901|1.4086379605250285|174|1
35.17335|6a843a99231452f476c34a55752c9458bcf00649|2.85|2015-01-08 14:07:00|1.4094857484078087|4|4133500053|174|0.6138907664563474|0|26|184|-80.70901|28|35.17335|SALAD DRESSINGS-LIQUID|1.43|1|KENS DRS LT BLUE CHEESE|e04dc890b30fd1b61727728f0d17a3f73c9aef09|1.0688318552138325|0.61471665291522548|00041335001690|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.323246|b25142f8ba5437fb99025ceaa1f33f30c8b1a3e1|5.29|2014-11-11 20:20:00|1.4102725052409182|3|7365111710|166|0.6165069451919168|0|1|160|-80.945176|25|35.323246|OLIVES|0.0|1|MARIO OLIVE MANZ 21|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|0.61833652052202714|00073651117106|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|1c659398bc2fa3ac9cfcba298b70c1f2f5c9e5b2|4.99|2015-02-26 14:45:00|80.945255278477163|3|4900005235|166|35.363594674235387|0|13|55|-80.760919|8|35.024332|REGULAR|1.0|23|DR PEPPER 8PK  7.5 OZ|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|35.37387923947206|00078000009712|CARBONATED BEVERAGES|BEVERAGE|-80.945176|80.945288563660853|343|1
35.323246|35c84f48561750861a177ee4c3ba7d9a152b5222|1.6|2014-12-02 21:07:00|1.4102725052409182|3||166|0.6165069451919168|0|1|531|-80.945176|64|35.323246|FRESH CORN|0.0|4|COO YELLOW CORN|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|0.61833652052202714|00204078000003|FRESH PRODUCE|PRODUCE|-80.945176|1.4127598348062935|166|2
35.323246|8f8ebe050623bb2b165c46e2ae5c13cb88b721c7|7.99|2014-12-27 16:41:00|80.945255278477163|3|8143450009|166|35.363594774347874|0|13|9948|-80.810056|886|35.219587|NFS-PREM-CAB SAUVIGNON|0.0|13|BLACKSTONE CAB SAUV|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|35.37387923947206|00081434500090|PREMIUM ($8-$10.99)|WINE|-80.945176|80.945198992313095|401|1
35.323246|8da6614ecd7c5a504fe7b328df62dc95150cba74|4.99|2015-02-23 19:50:00|1.4102725052409182|3|7203660022|166|0.6165069451919168|0|1|355|-80.945176|104|35.323246|FRESH GRILLING SAUSAGE|1.99|19|HT HOT ITALIAN SAUSAGE|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|0.61833652052202714|00072036600233|DINNER SAUSAGE|CASE READY MEATS|-80.945176|1.4127598348062935|166|1
35.323246|9f4b29f1354e98fa5c58c66bfb38bda9dfb4a8e1|7.49|2015-02-09 17:57:00|80.945255278477163|3|73753919040|166|35.363594696273381|0|13|1435|-80.770346|19|35.052812|SHELF STABLE SPREADS|0.0|1|SUNBUTTER CREAMY|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|35.37387923947206|00737539191205|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.945176|80.945275988741727|40|1
35.323246|4cd4cd9624b6def2eb4e88fe1ba2a4fde4b60753|7.49|2015-01-28 19:34:00|1.4102725052409182|3|73753919040|166|0.6165069451919168|0|1|1435|-80.945176|19|35.323246|SHELF STABLE SPREADS|0.0|1|SUNBUTTER CREAMY|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|0.61833652052202714|00737539191205|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|b460facf1530c48cd2608c78be480d84bbabf8c2|3.69|2015-02-15 18:33:00|1.4102725052409182|3|2500005542|166|0.6165069451919168|0|1|338|-80.945176|56|35.323246|OTHER FRUIT JUICES|0.0|3|SIMPLY CRANBERRY|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|0.61833652052202714|00025000046285|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.945176|1.4127598348062935|166|1
35.323246|7ef5460f3137321e133cc9a8346e731fce6e8f3d|3.19|2015-01-30 10:41:00|80.945255278477163|3|5000062231|166|35.363594653001627|0|13|326|-80.992182|54|35.103409|COOKIES/BROWNIES-REFRIGERATED|0.69|3|NESTLE CHOC. CHIP BAR COOKIES|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|35.37387923947206|00050000622313|DOUGH PRODUCTS|DAIRY|-80.945176|80.94529947414749|88|1
35.323246|e45e78946db7a1d2fa4bd8377efa935d1efd9c57|9.57|2015-02-26 15:33:00|80.945255278477163|3|5000062231|166|35.363594696273381|0|13|326|-80.770346|54|35.052812|COOKIES/BROWNIES-REFRIGERATED|0.0|3|NESTLE CHOC. CHIP BAR COOKIES|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|35.37387923947206|00050000622313|DOUGH PRODUCTS|DAIRY|-80.945176|80.945275988741727|40|3
35.323246|ce82e24e2e0e755e4d4377a1fc5ec679ef21f97a|4.59|2014-10-02 20:33:00|1.4102725052409182|3|75379200201|166|0.6165069451919168|0|1|130|-80.945176|20|35.323246|CRANBERRY JUICE/DRINKS-SHELF|2.3|1|NORTHLAND CRNBRY POMEGRANATE|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|0.61833652052202714|00753792002317|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|3dd134278208903192d616a80d9566531c7a97d8|1.79|2015-03-08 13:13:00|1.4102725052409182|3||166|0.6165069451919168|0|1|540|-80.945176|64|35.323246|FRESH CELERY|0.0|4|COO CELERY (RPC) 24'S|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|0.61833652052202714|00204070000001|FRESH PRODUCE|PRODUCE|-80.945176|1.4127598348062935|166|1
35.323246|a6d8240a118f74ee1ddb40cb17e800089dfb761b|8.49|2014-11-30 16:20:00|1.4102725052409182|3|2301200013|166|0.6165069451919168|0|1|1477|-80.945176|485|35.323246|SUSHI HYBRID|0.0|6|PLUS ROLL|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|0.61833652052202714|00023012000134|SUSHI|DELI|-80.945176|1.4127598348062935|166|1
35.323246|04ccc05a47741b5024ec09c617ddb94ccd39efe7|3.39|2015-03-07 11:19:00|80.945255278477163|3|61126917452|166|35.363594769659279|0|13|97|-80.737839|8|35.297134|ENERGY DRINKS|0.39|23|RED BULL RED EDITION|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|35.37387923947206|00611269174526|CARBONATED BEVERAGES|BEVERAGE|-80.945176|80.945209125424157|258|1
35.323246|16922de52ba5052179dd6800bc774af0f3cf5e49|1.9|2014-11-04 19:22:00|1.4102725052409182|3|4600028869|166|0.6165069451919168|0|1|77|-80.945176|272|35.323246|HISP SAUCES/SEASONINGS|0.4|1|OEP SEASONING TACO HOT & SPICY|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|0.61833652052202714|00046000288758|HISPANIC PREP. FOODS|G1 GROCERY|-80.945176|1.4127598348062935|166|2
35.323246|dc3c1eb2c7c49e20c0c7a2bb890f444ef0512693|1.39|2014-12-18 10:39:00|80.945255278477163|3|2200000488|166|35.363594653001627|0|13|48|-80.992182|7|35.103409|REGISTER GUM|0.0|1|(FE)ORBIT SPEARMINT GUM 14 PC|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|35.37387923947206|00022000004840|CANDY|G1 GROCERY|-80.945176|80.94529947414749|88|1
35.323246|2f803952f7196399d4e122862c51e537d9e17fcd|3.99|2015-02-01 10:18:00|1.4102725052409182|3|85420800508|166|0.6165069451919168|0|1|577|-80.945176|136|35.323246|OTHER MERCH FR MSC JUICE|1.49|4|ORG. SUJA CARROT CRUSH|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|0.61833652052202714|00854208005066|OTHER MERCHANDISE|PRODUCE|-80.945176|1.4127598348062935|166|1
35.323246|dfb9d0fa71ac0a6adba3512a01eecd023d32e697|2.99|2014-12-28 16:54:00|1.4102725052409182|3|8201110007|166|0.6165069451919168|0|1|1250|-80.945176|12|35.323246|SPECIALTY COOKIES|0.49|1|MURRAY GINGER SNAPS|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|0.61833652052202714|00082011100078|COOKIES|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|bdcb0c10a6e401fdc1c057d6c261c880bffc8413|3.99|2015-02-11 15:32:00|80.945255278477163|3|4157005982|166|35.363594674235387|0|13|1148|-80.760919|21|35.024332|ALMONDS|0.0|1|BLUE DIAMOND ALM SALT/VINEGAR|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|35.37387923947206|00041570053386|NUTS|G1 GROCERY|-80.945176|80.945288563660853|343|1
35.323246|4dc3413982cbc948af8dc62a02b272b72ba76542|4.29|2014-11-22 17:20:00|1.4102725052409182|3|4400002796|166|0.6165069451919168|0|1|90|-80.945176|13|35.323246|SNACK CRACKERS|2.15|1|TRISCUIT ORIGINAL|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|0.61833652052202714|00044000027957|CRACKERS|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|4d952a4689a49f4dc36ee8c911b0d69116ee2104|5.99|2014-12-02 08:13:00|80.945255278477163|3|85598300259|166|35.363594674235387|0|13|583|-80.760919|136|35.024332|NUTS|0.0|4|CREATIVE SNACK GRN BEAN CHIPS|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|35.37387923947206|00855983002592|OTHER MERCHANDISE|PRODUCE|-80.945176|80.945288563660853|343|1
35.323246|522fbf9c60f927c2e4b34a186767b2c8d3e31f10|2.19|2015-01-30 19:28:00|1.4102725052409182|3|4900005010|166|0.6165069451919168|0|1|55|-80.945176|8|35.323246|REGULAR|0.2|23|CLASSIC COKE 2 LT CONTOUR|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|0.61833652052202714|00049000050103|CARBONATED BEVERAGES|BEVERAGE|-80.945176|1.4127598348062935|166|1
35.323246|1bf53fe23a860267cb774e6a608e40423af15906|7.99|2015-02-05 09:28:00|80.945255278477163|3|64786510001|166|35.363594674235387|0|13|4195|-80.760919|1200|35.024332|COUGH & COLD REMEDY-ADULT|1.0|17|(FE)(JHK)AIRBORNE REG  ORANGE|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|35.37387923947206|00647865100010|COUGH/COLD/SINUS|HBC|-80.945176|80.945288563660853|343|1
35.323246|9a87b40557afc881c8edd6c047fc245f12fbcaff|2.99|2014-11-23 15:14:00|1.4102725052409182|3|7203670407|166|0.6165069451919168|0|1|5607|-80.945176|1512|35.323246|BRUSH-LINT|0.0|18|YH LINT ROLLER|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|0.61833652052202714|00072036704078|BROOMS/MOPS & BRUSHES|GM|-80.945176|1.4127598348062935|166|1
35.323246|f14daecb4124709f5c9807a58b3d7a5722b8df9c|5.99|2014-12-06 16:58:00|1.4102725052409182|3|88552321821|166|0.6165069451919168|0|1|1403|-80.945176|389|35.323246|THAW AND SELL PIES|0.0|14|"8"" NO SGR ADD PUMPKIN PIE"|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|0.61833652052202714|00885523218213|PIES|BAKERY|-80.945176|1.4127598348062935|166|1
35.323246|b0d1cdc897716f56eab7b2df632dc552b150f484|10.99|2014-09-21 18:15:00|1.4102725052409182|3|8273434124|166|0.6165069451919168|0|1|9955|-80.945176|886|35.323246|NFS-PREM-MALBEC|0.0|13|TRIVENTO MALBEC|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|0.61833652052202714|00082734341246|PREMIUM ($8-$10.99)|WINE|-80.945176|1.4127598348062935|166|1
35.323246|2239034cfd3b5c07bacd54fbbc18333665136f03|10.99|2014-12-31 21:10:00|1.4102725052409182|3|8500001773|166|0.6165069451919168|0|1|9983|-80.945176|889|35.323246|NFS-SPARKLING|0.0|13|CB-LA MARCA PROSECCO|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|0.61833652052202714|00085000017739|SPARKLING|WINE|-80.945176|1.4127598348062935|166|1
35.323246|8eb2b2330aff2fa819b5426738a8b3eaa7ea1d98|1.79|2014-12-29 14:49:00|1.4102725052409182|3|5100005977|166|0.6165069451919168|0|1|212|-80.945176|33|35.323246|CONDENSED SOUP|0.54|1|CAMP HLTHY REQ HOME CHICK NOOD|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|0.61833652052202714|00051000167217|SOUP|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|d0c14766716ada8a825f19f6347d1d38f4f9562d|3.99|2015-01-05 13:16:00|80.945255278477163|3|72243011016|166|35.363594674235387|0|13|577|-80.760919|136|35.024332|OTHER MERCH FR MSC JUICE|0.0|4|ORG. GT KOMBUCHA CRANBERRY|e4245e980d62003bc90fdaa9e3692bef8fbe3552|2.788003169817851|35.37387923947206|00722430300160|OTHER MERCHANDISE|PRODUCE|-80.945176|80.945288563660853|343|1
35.412407|6e5070a743d429899bacf047b586ce3095eefaca|5.54|2015-01-04 09:39:00|1.4102725052409182|4|7433610202|68|0.6180630982062877|0|1|318|-80.662946|52|35.412407|SHREDDED/GRATED CHEESE|0.0|3|HC SHREDDED MOZZARELLA|e48a051bd3d597842fef40a1115d932d57d81bba|2.319680121896889|0.61833652052202714|00074336102028|CHEESE|DAIRY|-80.662946|1.40783399205839|68|2
35.412407|4423264f67895198cf3ae5c6d32791a22805ba78|8.58|2014-10-25 15:04:00|1.4102725052409182|4|2840016014|68|0.6180630982062877|0|1|201|-80.662946|31|35.412407|POTATO CHIPS|2.14|1|LAYS WAVY REGULAR|e48a051bd3d597842fef40a1115d932d57d81bba|2.319680121896889|0.61833652052202714|00028400160209|SNACKS|G1 GROCERY|-80.662946|1.40783399205839|68|2
35.412407|7bac2605202f572470dfde70f795720ce69d9045|2.99|2015-02-01 13:32:00|1.4102725052409182|4|7433610102|68|0.6180630982062877|0|1|342|-80.662946|57|35.412407|FRESH MILK|0.0|3|HIGHLAND CREST WHOLE MILK|e48a051bd3d597842fef40a1115d932d57d81bba|2.319680121896889|0.61833652052202714|00074336879203|MILK|DAIRY|-80.662946|1.40783399205839|68|1
35.412407|5730937e7cbd001845972396af5abfda6eb16f13|2.69|2014-10-11 12:17:00|1.4102725052409182|4|7203630050|68|0.6180630982062877|0|1|184|-80.662946|28|35.412407|SALAD DRESSINGS-LIQUID|0.81|1|HT DRS VIN FF ITALIAN|e48a051bd3d597842fef40a1115d932d57d81bba|2.319680121896889|0.61833652052202714|00072036300522|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.662946|1.40783399205839|68|1
35.412407|b11a01129fd506b96a04729ffab84d3ee48a3a7f|3.79|2015-01-11 13:06:00|1.4102725052409182|4|4850002013|68|0.6180630982062877|0|1|335|-80.662946|56|35.412407|ORANGE JUICE-REGRIGERATED|0.79|3|TROP  50 NO PULP|e48a051bd3d597842fef40a1115d932d57d81bba|2.319680121896889|0.61833652052202714|00048500020135|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.662946|1.40783399205839|68|1
35.412407|c03d9b21ff64cc54eb273a10f5724d276801ca66|6.02|2014-11-23 12:17:00|1.4102725052409182|4|20165700000|68|0.6180630982062877|0|1|297|-80.662946|49|35.412407|GROUND BEEF|0.67|2|HT GROUND BEEF CHUCK 80% LEAN|e48a051bd3d597842fef40a1115d932d57d81bba|2.319680121896889|0.61833652052202714|00201657000003|BEEF|MEAT|-80.662946|1.40783399205839|68|1
35.04711|eb8fef8013d624d2b3ebd857b7241df5a5ae0f50|9.99|2014-11-22 15:31:00|80.648225123995502|3|7203678030|129|35.062250797108646|0|30|458|-80.699909|82|35.002628|CRAFT BEER|0.0|16|HT CREATE YOUR OWN SAMPLER|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|35.078006462436761|00072036780300|DOMESTIC BEER|BEER|-80.64817|80.648182915224893|477|1
35.04711|e91de5bae06134842c5f441bac136d0c582e9509|9.99|2015-02-06 14:25:00|80.648225123995502|3|7203678030|129|35.062250797108646|0|30|458|-80.699909|82|35.002628|CRAFT BEER|0.0|16|HT CREATE YOUR OWN SAMPLER|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|35.078006462436761|00072036780300|DOMESTIC BEER|BEER|-80.64817|80.648182915224893|477|1
35.04711|c03ea8e2c866dd2b75b6aa83dc922555a6ca2e47|9.99|2014-09-26 11:50:00|80.648225123995502|3|7203678030|129|35.062250797108646|0|30|458|-80.699909|82|35.002628|CRAFT BEER|0.0|16|HT CREATE YOUR OWN SAMPLER|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|35.078006462436761|00072036780300|DOMESTIC BEER|BEER|-80.64817|80.648182915224893|477|1
35.04711|5fa0ef9715c1cf968d2290612c80ee71d07afd06|3.99|2014-12-17 12:37:00|80.648225123995502|3|7203676382|129|35.062250796829829|0|30|122|-80.699686|19|35.000049|HONEY|0.99|1|HTO HONEY WILDFLOWER|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|35.078006462436761|00072036763822|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.64817|80.648183394113659|249|1
35.04711|2eb96f2f062ca413eacab9adc371d53cd6301ee6|9.99|2014-09-29 13:25:00|80.648225123995502|3|7203678030|129|35.062250800798374|0|30|458|-80.7007|82|35.06858|CRAFT BEER|0.0|16|HT CREATE YOUR OWN SAMPLER|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|35.078006462436761|00072036780300|DOMESTIC BEER|BEER|-80.64817|80.648170261798327|273|1
35.04711|3ff9b5c2933379c266e20c91c45f475ecd3ad996|3.59|2015-02-14 13:25:00|80.648225123995502|3|7203695890|129|35.062250796829829|0|30|1654|-80.699686|381|35.000049|DESSERT CAKES|0.0|14|GRANDE FINALE CAKE SLICE|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|35.078006462436761|00072036958907|CAKES|BAKERY|-80.64817|80.648183394113659|249|1
35.04711|cf3b7578aa5a7ac020e0974aaf1885ccdcc5f8a2|19.98|2014-10-20 13:53:00|80.648225123995502|3|7203678030|129|35.062250797108646|0|30|458|-80.699909|82|35.002628|CRAFT BEER|0.0|16|HT CREATE YOUR OWN SAMPLER|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|35.078006462436761|00072036780300|DOMESTIC BEER|BEER|-80.64817|80.648182915224893|477|2
35.04711|5e95c7f5b3482cf174e68e8654ea325bdba8f015|1.29|2015-02-20 19:14:00|1.4091206135396188|3|4146039883|129|0.6116874628086298|0|47|75|-80.64817|34|35.04711|GRAVY MIXES|0.29|1|PIONEER CNTRY SAUSAGE GRAVY MX|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00041460398832|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|524bb9c494a8bde0674ec88554e097678e1d4582|2.49|2014-11-23 10:04:00|1.4091206135396188|3|4410010755|129|0.6116874628086298|0|47|341|-80.64817|57|35.04711|CREAMERS|1.24|3|BAILEYS MUDSLIDE CREAMER|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00044100107665|MILK|DAIRY|-80.64817|1.407576102208115|129|1
35.04711|16856f7aed50c8871b603b34ff76dfd2cb4ef1f6|0.65|2014-12-11 08:23:00|1.4091206135396188|3|5000042264|129|0.6116874628086298|0|47|154|-80.64817|24|35.04711|NFS-CAT FOOD WET|0.1|1|FRISKIES SPECIAL DIET CHICKEN|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00050000425242|PET FOOD/SUPPLIES|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|2165f18835161301ee49867f239d4021193bbce3|0.65|2014-11-09 18:43:00|1.4091206135396188|3|5000042264|129|0.6116874628086298|0|47|154|-80.64817|24|35.04711|NFS-CAT FOOD WET|0.15|1|FRISKIES MARINERS CATCH|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00050000425044|PET FOOD/SUPPLIES|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|7e2cc3b1419bc4332e807a0b13a7ef7be52c954f|0.65|2014-11-01 15:28:00|1.4091206135396188|3|5000042264|129|0.6116874628086298|0|47|154|-80.64817|24|35.04711|NFS-CAT FOOD WET|0.15|1|FRISKIES SPECIAL DIET CHICKEN|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00050000425242|PET FOOD/SUPPLIES|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|df373bb8c8c371339e711114cc6f75d551b05dcb|0.65|2014-11-23 12:13:00|1.4091206135396188|3|5000042264|129|0.6116874628086298|0|47|154|-80.64817|24|35.04711|NFS-CAT FOOD WET|0.1|1|FRISKIES CANNED SHRED CHX/SALM|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00050000445691|PET FOOD/SUPPLIES|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|50411a4c0f047916f9faa6d5e657103bd5e017ab|1.99|2014-12-28 10:32:00|1.4091206135396188|3|78616233800|129|0.6116874628086298|0|47|31|-80.64817|4|35.04711|NON CARBONATED WATER|0.99|1|CB SMARTWATER 1 LTR PET SINGLE|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00786162338006|BOTTLED WATER|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|aeba19a2013dcac5dd9326d58731d0e2d9d50f76|3.99|2015-02-12 17:29:00|1.4091206135396188|3|78843411430|129|0.6116874628086298|0|47|4784|-80.64817|1230|35.04711|DRINKS-PROTEIN|1.99|17|(FE) OH YEAH RTD VANILLA|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00788434114356|SPORTS NUTRITIONAL|HBC|-80.64817|1.407576102208115|129|1
35.04711|b6984d98a926d29afbb88abb13f524f8bbfe26d9|1.89|2014-11-13 13:34:00|1.4091206135396188|3|2700038249|129|0.6116874628086298|0|47|70|-80.64817|11|35.04711|KETCHUP|0.89|1|HUNTS KETCHUP 24|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00027000382493|CONDIMENTS|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|ee0f30be6b68d33416a0ddd12ce8392acb0f5902|2.89|2014-12-31 15:49:00|1.4091206135396188|3|5150028064|129|0.6116874628086298|0|47|12|-80.64817|2|35.04711|PANCAKE MIXES|0.92|1|H JACK WHEAT BLND BLUBRY PNCKE|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00051500101476|BAKING MIXES|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|dd98dd156fe9f11cb707837bddd3fb489225e00c|1.39|2015-02-22 11:34:00|1.4091206135396188|3|5210094269|129|0.6116874628086298|0|47|80|-80.64817|34|35.04711|SEASONING PACKETS|0.42|1|E  MC CHILI SEASONING MIX|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00052100091501|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|ef1b79ee03263077d6c07120800f6a5cc04f03d1|2.66|2014-09-22 12:54:00|1.4091206135396188|3|7047043332|129|0.6116874628086298|0|47|685|-80.64817|61|35.04711|GREEK|0.66|3|YOPLAIT GREEK 100 BLK CHERRY|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00070470435794|YOGURT|DAIRY|-80.64817|1.407576102208115|129|2
35.04711|d604b038d9bb59d05a2e8ea19414e5f58f67313c|0.65|2015-01-18 16:22:00|1.4091206135396188|3|5000042264|129|0.6116874628086298|0|47|154|-80.64817|24|35.04711|NFS-CAT FOOD WET|0.15|1|FRISKIES SHREDDED SALMON&SAUCE|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00050000572014|PET FOOD/SUPPLIES|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|bfca7a1794df7f217038f6fda9636f21a94752b1|3.79|2015-01-30 12:22:00|1.4091206135396188|3|7203688014|129|0.6116874628086298|0|47|581|-80.64817|136|35.04711|FRESH SALSA|1.66|4|HT FRESH MEDIUM SALSA|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00072036880222|OTHER MERCHANDISE|PRODUCE|-80.64817|1.407576102208115|129|1
35.04711|77ce4c035c4443a0731551560a6bd957d71086db|3.98|2015-02-08 11:35:00|1.4091206135396188|3|81162002002|129|0.6116874628086298|0|47|1263|-80.64817|57|35.04711|GOOD FOR YOU MILK|1.98|3|FAIRLIFE 2% CHOC MILK SINGLE|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00811620020039|MILK|DAIRY|-80.64817|1.407576102208115|129|2
35.04711|3f61f1fabbd858f661956a532c671036621b85de|2.19|2014-10-07 09:18:00|1.4091206135396188|3|1200004139|129|0.6116874628086298|0|47|854|-80.64817|32|35.04711|LIQUID ICED COFFEES|0.2|1|STARBUCKS ICED COF CHOC MLK LC|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00012000041419|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|34ea292d357d0ca5a6fd3e11973cd2e5028f3f61|0.69|2014-10-13 14:13:00|1.4091206135396188|3|82927400616|129|0.6116874628086298|0|47|154|-80.64817|24|35.04711|NFS-CAT FOOD WET|0.04|1|MEOW MIX MRKT SEL SAL & CRAB|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00829274006163|PET FOOD/SUPPLIES|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|16c9b8ee0c4a2fa4b4e4c3eaf4f535eeb598c0f2|1.55|2014-11-30 13:06:00|1.4091206135396188|3|78616201000|129|0.6116874628086298|0|47|31|-80.64817|4|35.04711|NON CARBONATED WATER|0.55|1|VIT WATER REVIVE 20 OZ|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00786162110008|BOTTLED WATER|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|5be9fc8ccc49f041450910545ac20c183cca133b|18.76|2014-12-13 13:47:00|1.4091206135396188|3|4900002468|129|0.6116874628086298|0|47|54|-80.64817|8|35.04711|DIET|9.38|23|COKE ZERO .5L 6PK PET|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00049000045840|CARBONATED BEVERAGES|BEVERAGE|-80.64817|1.407576102208115|129|4
35.04711|a858814c08d3135a4a3e746bf5580981bce021bb|3.99|2014-09-28 09:41:00|80.648225123995502|3|7203663995|129|35.062250796284211|0|30|342|-80.654118|57|35.123768|FRESH MILK|1.02|3|HARRIS TEETER 2% MILK|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|35.078006462436761|00072036639981|MILK|DAIRY|-80.64817|80.648184284889595|473|1
35.04711|34a23349d1c9c9aad16d9c49a324ad7c98e0bc7c|3.99|2014-10-28 12:09:00|1.4091206135396188|3|4470003050|129|0.6116874628086298|0|47|840|-80.64817|102|35.04711|TUBS|0.99|19|OM DELI FRESH HAM/TURK COMBO|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00044700034071|LUNCHMEATS|CASE READY MEATS|-80.64817|1.407576102208115|129|1
35.04711|fef30aba9ebaaeffdbc65a7db0479bf9abc770b5|1.55|2015-01-24 13:27:00|1.4091206135396188|3|78616201000|129|0.6116874628086298|0|47|31|-80.64817|4|35.04711|NON CARBONATED WATER|0.55|1|VIT WATER ZERO XXX|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00786162002969|BOTTLED WATER|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|57ff9ab7332053fc0a6e883a4ce623e642084fbb|3.49|2015-01-17 17:08:00|1.4091206135396188|3|2840024053|129|0.6116874628086298|0|47|198|-80.64817|31|35.04711|CORN CHIPS|1.74|1|FRITOS REGULAR|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00028400240536|SNACKS|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|dd00efc2a751898ac8b0ead6a7648cb7ca7bde28|3.35|2015-02-13 12:03:00|1.4091206135396188|3|2529300098|129|0.6116874628086298|0|47|1263|-80.64817|57|35.04711|GOOD FOR YOU MILK|0.0|3|SILK PURE CASHEW MILK|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00025293002746|MILK|DAIRY|-80.64817|1.407576102208115|129|1
35.04711|605812aab4ebf2e3483795f6e92491106cfab6f0|3.89|2015-01-15 21:29:00|1.4091206135396188|3|7457000400|129|0.6116874628086298|0|47|275|-80.64817|45|35.04711|SUPER PREMIUM ICE CREAM|0.55|5|H DAZS BUTTER PECAN-|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00074570114009|ICE CREAM|FROZEN|-80.64817|1.407576102208115|129|1
35.04711|653ed379bc069e0f77692e94cb5f79cc7c45d027|3.99|2014-10-20 13:53:00|80.648225123995502|3|4157005982|129|35.062250797108646|0|30|1148|-80.699909|21|35.002628|ALMONDS|0.99|1|B D ALMONDS B JALAPENO SMK HSE|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|35.078006462436761|00041570052327|NUTS|G1 GROCERY|-80.64817|80.648182915224893|477|1
35.04711|fe452d798cb5aef3cd3a76a5bd79f73643a2d5b6|5.39|2015-03-06 13:41:00|1.4091206135396188|3|5000001547|129|0.6116874628086298|0|47|152|-80.64817|24|35.04711|NFS-CAT FOOD DRY|1.89|1|FRISKIES RISE&SHINE DRY CATFD|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00050000585045|PET FOOD/SUPPLIES|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|e8e1ce9232c24a0ee18b6e5f6897d74265c18aa3|3.69|2014-11-02 08:54:00|1.4091206135396188|3|2340099821|129|0.6116874628086298|0|47|393|-80.64817|68|35.04711|NFS-AIR FRESHENERS|0.7|1|RENUZIT PEARLS AFTER THE RAIN|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00023400998210|FRESHENERS/DEODORIZERS|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|9c1b64686db19aeaacf9447926c57c3475ba1e34|2.0|2014-09-11 09:47:00|1.4091206135396188|3||129|0.6116874628086298|0|47|565|-80.64817|64|35.04711|REDUCED PRODUCE|0.0|4|PRODUCE REWRAP BY CT|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00204845000007|FRESH PRODUCE|PRODUCE|-80.64817|1.407576102208115|129|2
35.04711|13eb8fc27a234bbbd1fbe07af54f2baf73404d38|4.79|2014-11-22 15:32:00|80.648225123995502|3|18685200031|129|35.062250797108646|0|30|275|-80.699909|45|35.002628|SUPER PREMIUM ICE CREAM|2.39|5|TALENTI CARAMEL COOKIE GELATO|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|35.078006462436761|00186852000334|ICE CREAM|FROZEN|-80.64817|80.648182915224893|477|1
35.04711|a150fad46ea06dc7b8db74527feb521094c31355|1.69|2014-11-11 14:12:00|1.4091206135396188|3|4900000044|129|0.6116874628086298|0|47|54|-80.64817|8|35.04711|DIET|0.0|23|CB DIET DR PEPPER 20OZ NR|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00078000083408|CARBONATED BEVERAGES|BEVERAGE|-80.64817|1.407576102208115|129|1
35.04711|11c1533f36e0f858029fd9e735c7b5a28b47c950|9.99|2014-09-14 13:08:00|1.4091206135396188|3|2301286482|129|0.6116874628086298|0|47|1477|-80.64817|485|35.04711|SUSHI HYBRID|0.0|6|"CHEF SAMPLER ""B"""|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00023012864828|SUSHI|DELI|-80.64817|1.407576102208115|129|1
35.04711|d53124851d5eafcd55e21498995724e458f55d4b|3.99|2015-02-07 11:19:00|80.648225123995502|3|7166261216|129|35.062250796565678|0|30|6570|-80.760919|1564|35.024332|CHALK|0.0|18|CRAYOLA SIDEWALK CHALK|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|35.078006462436761|00071662612160|SCHOOL & OFFICE SUPPLY|GM|-80.64817|80.648183832537129|343|1
35.04711|2eec2a5ace1941d31637c3e8c591b8d26f9b7031|4.29|2015-01-06 15:44:00|1.4091206135396188|3|2840006399|129|0.6116874628086298|0|47|204|-80.64817|31|35.04711|TORTILLA CHIPS|0.29|1|TOSTITOS ROLLS|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|0.61242566243833529|00028400288651|SNACKS|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|193bfae9e03adc512499a9da3afb40aacca0aadd|6.98|2015-02-09 13:58:00|80.648225123995502|3|7203604187|129|35.062250796829829|0|30|335|-80.699686|56|35.000049|ORANGE JUICE-REGRIGERATED|1.02|3|HT PREM GROVES BEST ORANGE JCE|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|35.078006462436761|00072036041845|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.64817|80.648183394113659|249|2
35.04711|e5c7aa96a9c48778ce83f41ffe87b83a00a15ad5|3.38|2014-10-04 13:29:00|80.648225123995502|3|79386630001|129|35.062250797108646|0|30|458|-80.699909|82|35.002628|CRAFT BEER|0.0|16|LEFT HAND SAWTOOTH ALE 12OZ|e7e42907edada453cd0cfd5d6e9b1a05e775819b|1.0461927715475534|35.078006462436761|00793866300017|DOMESTIC BEER|BEER|-80.64817|80.648182915224893|477|2
35.053394|e48ce4dbd901a819f2cd9118a1e08690984c1264|2.99|2014-12-24 06:50:00|80.848351720559364|4|86322300000|11|35.073487954212595|0|25|312|-80.78468|51|35.096737|BUTTER|0.0|3|SHANNONGOLD SALT BUTTER 8OZ|e871b88da1717e8ed1c7f0ce916fae4fa94f6d1d|1.3884440910102207|35.082633588753836|00863223000000|BUTTER & MARGARINE|DAIRY|-80.848528|80.848546164672939|30|1
35.053394|20cf5890539103766792fe824f85eac45bb1cc05|11.99|2014-09-10 13:23:00|80.848351720559364|4|20595400000|11|35.073487958832274|0|25|1823|-80.847383|410|35.024464|BH HAM|2.0|6|BOARS HEAD TRIO|e871b88da1717e8ed1c7f0ce916fae4fa94f6d1d|1.3884440910102207|35.082633588753836|00205954000001|BH MEAT|DELI|-80.848528|80.848535269471213|317|1
35.053394|791be367a7a6131496e12eebb4409499932d92dc|1.49|2015-01-26 12:49:00|80.848351720559364|4|4900005537|11|35.073487856512628|0|25|55|-80.66939|8|35.28326|REGULAR|0.49|23|CLASSIC 1.25 LITER BOTTLE|e871b88da1717e8ed1c7f0ce916fae4fa94f6d1d|1.3884440910102207|35.082633588753836|00049000055375|CARBONATED BEVERAGES|BEVERAGE|-80.848528|80.848606679386165|46|1
35.053394|7abfd8cafce4c0a6abc3a1986362ca19f41466ea|5.99|2014-10-17 19:37:00|80.848351720559364|4|7203695643|11|35.073487959257051|0|25|1663|-80.816172|381|35.059823|CREME CAKE|0.0|14|44 OZ CHOC CREME CAKE|e871b88da1717e8ed1c7f0ce916fae4fa94f6d1d|1.3884440910102207|35.082633588753836|00072036956644|CAKES|BAKERY|-80.848528|80.848533231147655|66|1
35.444064|d2abedcc615cbd21cd9b45be5595743142e63db7|2.99|2014-09-28 12:15:00|1.4102725052409182|3|7203698553|121|0.6186156170875914|0|1|427|-80.995484|72|35.444064|NFS-TOILET TISSUE|0.49|1|HT BATH PLUSH 4RL|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00072036985538|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|6ac51530328856e12d1e913de544ffb4838a1e52|3.0|2015-01-17 10:26:00|1.4102725052409182|3|7203697890|121|0.6186156170875914|0|1|61|-80.995484|9|35.444064|RTE CEREAL ADULT|0.0|1|HT CER SPECIAL IT'S BERRY|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00072036978905|CEREAL|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|7aaeeb699ae86655ee43d4acc854cd9e1cb7e753|2.39|2014-10-02 08:58:00|1.4102725052409182|3|7203698241|121|0.6186156170875914|0|1|442|-80.995484|76|35.444064|NFS-COOKING-STORAGE BAGS|0.72|1|YH RESEALABLE SANDWICH BAGS|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00072036982414|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|0cf69f4bc5be0d0e49d68f9cc9541fd9b7ae8664|3.0|2015-01-31 09:35:00|1.4102725052409182|3|7203697890|121|0.6186156170875914|0|1|61|-80.995484|9|35.444064|RTE CEREAL ADULT|0.0|1|HT CER SPECIAL IT'S BERRY|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00072036978905|CEREAL|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|95f040600880a61f2b82eaa3c7853835efefddb8|4.65|2014-10-30 09:41:00|1.4102725052409182|3|7218063473|121|0.6186156170875914|0|1|284|-80.995484|892|35.444064|SUPER PREMIUM PIZZA|0.66|5|RED BARON RISING SAU&PEPP PZZA|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00072180567345|FROZEN PIZZA|FROZEN|-80.995484|1.413637875046387|121|1
35.444064|2dfd735108d92a6f9ea6f552512cb4a5526f7750|3.0|2015-01-22 09:22:00|1.4102725052409182|3|7203697890|121|0.6186156170875914|0|1|61|-80.995484|9|35.444064|RTE CEREAL ADULT|0.0|1|HT CER SPECIAL IT'S BERRY|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00072036978905|CEREAL|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|fea7bc1f3306420c837c6efca8a2e7857f188847|3.99|2015-03-05 09:10:00|1.4102725052409182|3|7203688049|121|0.6186156170875914|0|1|562|-80.995484|64|35.444064|FRESH CUT FRUIT|0.5|4|HT MIXED FRUIT CHUNKS 16OZ|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00072036880499|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|72f716b9eae14c86a831714670d237859c5d0b41|1.34|2015-02-10 16:22:00|80.995508130988839|3|7203641111|121|35.450744791874904|0|40|242|-80.861571|39|35.444615|CANNED BEANS|0.0|1|HT PEAS BLACKEYE|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|35.466476270328783|00072036411143|VEGETABLES-CAN/JAR|G1 GROCERY|-80.995484|80.995489033769758|340|2
35.444064|3ffe08858676830fcb70ed78b6f3c9bc553b97ee|1.17|2014-12-29 08:49:00|1.4102725052409182|3|7203628014|121|0.6186156170875914|0|1|162|-80.995484|25|35.444064|PICKLES|0.0|1|HT CHIPS BREAD & BUTTER 16|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00072036280145|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|b611ced76a5c95383c0172c2f65c7e62f04c0e71|2.85|2014-11-13 09:20:00|1.4102725052409182|3|3040077852|121|0.6186156170875914|0|1|427|-80.995484|72|35.444064|NFS-TOILET TISSUE|0.0|1|ANGEL SOFT SOFT/STRONG 4DR|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00030400778520|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|62f579343f4c0f80949ef039dbd2e56951429758|3.69|2014-09-25 09:42:00|1.4102725052409182|3|4178000159|121|0.6186156170875914|0|1|201|-80.995484|31|35.444064|POTATO CHIPS|0.9|1|UTZ CLASSIC REGULAR|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00041780001597|SNACKS|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|1aef93503949430fe3652a3d830ef668f34ca43b|4.49|2014-12-18 09:21:00|1.4102725052409182|3|4470003050|121|0.6186156170875914|0|1|840|-80.995484|102|35.444064|TUBS|2.25|19|OM DELI FRESH SMOKED HAM|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00044700030486|LUNCHMEATS|CASE READY MEATS|-80.995484|1.413637875046387|121|1
35.444064|0b6174f0cdbde712e165ce65c3a2b14e6e56f3ee|3.79|2015-02-05 14:02:00|1.4102725052409182|3|4850002013|121|0.6186156170875914|0|1|335|-80.995484|56|35.444064|ORANGE JUICE-REGRIGERATED|0.79|3|TROPICANA PP HOMESTYLE|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00048500301395|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|f8d892c700162d4dcc5e1007da6f2c40df211ffd|8.99|2014-12-26 13:21:00|80.995508130988839|3|8066095605|121|35.450744792711497|0|40|459|-80.737839|83|35.297134|IMPORT BEER|0.0|16|CORONA EXTRA 6PK 12OZ BTL|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|35.466476270328783|00080660956053|IMPORT BEER|BEER|-80.995484|80.995486914639599|258|1
35.444064|8859313858339f1b7b1f2fe68ffc4aa2581e5884|4.89|2015-02-25 08:01:00|1.4102725052409182|3|3700084609|121|0.6186156170875914|0|1|3592|-80.995484|1050|35.444064|HAIR STYLING HAIR SPRAY|0.9|17|VS FLEXIBLE HOLD HAIR SPRAY|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00037000846925|HAIR STYLING|HBC|-80.995484|1.413637875046387|121|1
35.444064|9cd38c11c8b88c3631da80018542c01b5473ad36|2.85|2014-11-06 09:06:00|1.4102725052409182|3|4400000055|121|0.6186156170875914|0|1|88|-80.995484|13|35.444064|FLAKED SODA CRACKERS|0.35|1|NABISCO PREMIUMS|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00044000000578|CRACKERS|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|4f930480a326da999d0989230bc62857522a511c|3.34|2014-10-23 09:25:00|1.4102725052409182|3|7203643010|121|0.6186156170875914|0|1|252|-80.995484|45|35.444064|PREMIUM ICE CREAM|0.0|5|HT SMTH & CRMY CARAMEL DEL IC|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00072036981752|ICE CREAM|FROZEN|-80.995484|1.413637875046387|121|1
35.444064|6a924edaaef4ee0852d7496e179deaf9bbe21009|2.89|2015-02-15 15:32:00|1.4102725052409182|3|7203655029|121|0.6186156170875914|0|1|331|-80.995484|52|35.444064|NATURAL SLICED|1.22|3|HT MEDIUM CHEDDAR SLICES|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00072036983930|CHEESE|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|3ff038a659c1f576c36409943980f77bc14d07ec|1.69|2015-02-02 18:42:00|1.4102725052409182|3|7203688003|121|0.6186156170875914|0|1|527|-80.995484|64|35.444064|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00072036880031|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|d462183f6e5a789d056d1063f21a50688ddc8535|1.57|2014-10-13 13:18:00|1.4102725052409182|3|7203697658|121|0.6186156170875914|0|1|44|-80.995484|6|35.444064|TOASTER PASTRIES-SHELF STABLE|0.79|1|HT TSTR PASTRY UF STRAWBERRY|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00072036976567|BREAKFAST FOODS|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|f819cac578e86aabffb2b803788161cc25d30365|3.99|2014-09-17 15:58:00|80.995508130988839|3|7203695676|121|35.450744792456739|0|40|1656|-80.8955|381|35.4437|CUP CAKES|0.5|14|FFM MINI VANILLA CUPCAKES|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|35.466476270328783|00072036956767|CAKES|BAKERY|-80.995484|80.995487691114619|272|1
35.444064|411bb4e45d840309a6933612f01527bab83a9330|2.5|2014-11-29 10:52:00|1.4102725052409182|3|7203697755|121|0.6186156170875914|0|1|81|-80.995484|9|35.444064|RTE CEREAL KIDS|0.83|1|HT CER FROSTED FLAKES|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00072036977557|CEREAL|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|10358cbd880f18648c217574722a844836e21e51|2.5|2014-11-20 08:37:00|1.4102725052409182|3|7203697755|121|0.6186156170875914|0|1|81|-80.995484|9|35.444064|RTE CEREAL KIDS|0.53|1|HT CER FROSTED FLAKES|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00072036977557|CEREAL|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|8a2b8549829c4a2adc758227ab9914998deb9675|3.29|2014-09-13 10:26:00|1.4102725052409182|3|5250005002|121|0.6186156170875914|0|1|182|-80.995484|28|35.444064|MAYO|0.0|1|DUKES MAYONNAISE 16|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00052500050023|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|4cb22fc26a27dd6c32d1aa08c1114ce4a52bea56|3.29|2015-02-10 18:00:00|1.4102725052409182|3|5210002570|121|0.6186156170875914|0|1|220|-80.995484|34|35.444064|PEPPER|0.0|1|MC LEMON PEPPER CA. STYLE|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00052100025704|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|b195de2ca1d465e359f6c86ae1fe384a7f06a1b2|2.77|2015-02-25 16:22:00|1.4102725052409182|3|3338353030|121|0.6186156170875914|0|1|523|-80.995484|64|35.444064|FRESH POTATOES|0.0|4|RUSSET POTATO 8LB BAG|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00033383530307|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|42ee49326dfc5157fde5c27e46c685a2aa9efd65|3.39|2014-12-11 09:03:00|1.4102725052409182|3|2113150605|121|0.6186156170875914|0|1|1279|-80.995484|48|35.444064|SINGLE SERVE FLAVOR|0.89|5|M CALLENDER FETTUCINI CHK/BROC|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00021131504755|FROZEN MEALS|FROZEN|-80.995484|1.413637875046387|121|1
35.444064|bad0b1a020ea431fe6c2087598c2f2c746e58202|1.34|2015-01-05 09:39:00|1.4102725052409182|3|2100001087|121|0.6186156170875914|0|1|714|-80.995484|274|35.444064|MICROWAVE MEALS|0.0|1|KRAFT MAC CUP ORIGINAL|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00021000010875|PREP FOODS DINNERS|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|89180ccf112f7b984f86f2143184bc03fa9ccfb3|3.59|2014-10-16 09:07:00|1.4102725052409182|3|7641090137|121|0.6186156170875914|0|1|1255|-80.995484|13|35.444064|LUNCH BOX CRACKERS|0.59|1|LANCE R/F TOASTCHEESE|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00076410523330|CRACKERS|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|b7dbdede1e979b5adc1ca9f4794d21d9f9dfe696|1.79|2014-12-08 13:16:00|1.4102725052409182|3|5100001047|121|0.6186156170875914|0|1|212|-80.995484|33|35.444064|CONDENSED SOUP|0.12|1|CAMP COND BEEF VEGETABL BARLEY|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00051000011114|SOUP|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|8a6afa26eb889b279c787e42eca23b08f2a2ad9e|12.99|2015-01-04 14:38:00|80.995508130988839|3|1338585182|121|35.450744792711497|0|40|9951|-80.737839|886|35.297134|NFS-PREM-PINOT GRIS/GRIG|0.0|13|BILTMORE PINOT GRIGIO|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|35.466476270328783|00013385851822|PREMIUM ($8-$10.99)|WINE|-80.995484|80.995486914639599|258|1
35.444064|bc18ebe0c4f864b954eecfb1abb442bf5d19ac68|3.19|2014-11-18 19:06:00|1.4102725052409182|3|7294561221|121|0.6186156170875914|0|1|1039|-80.995484|166|35.444064|DINNER ROLLS|0.0|7|SARA LEE HAWAIIAN ROLLS PP|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00072945612211|MEAL ACCOMPANIMENT|COMMERCIAL BAKERY|-80.995484|1.413637875046387|121|1
35.444064|19f4d27d40e12a70e0ff7047005c89ac79af0877|2.97|2014-11-25 13:38:00|1.4102725052409182|3|7203658035|121|0.6186156170875914|0|1|358|-80.995484|100|35.444064|REGULAR BACON|0.0|19|HT LOW SALT SLICED BACON|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00072036590237|BACON|CASE READY MEATS|-80.995484|1.413637875046387|121|1
35.444064|903802df30bc58ed2a9198e727f10fa18611cb79|2.49|2014-12-07 13:07:00|1.4102725052409182|3|61611206143|121|0.6186156170875914|0|1|581|-80.995484|136|35.444064|FRESH SALSA|0.0|4|WHOLLY SALSA AVO VERDE|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00616112061435|OTHER MERCHANDISE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|b9efa90f9cfd2d5960431af0dff35d6f2203be04|0.66|2015-01-13 09:46:00|1.4102725052409182|3||121|0.6186156170875914|0|1|502|-80.995484|64|35.444064|FRESH BANANAS|0.0|4|BANANAS, YELLOW|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|2493b6c701b65e919e3e66e20ca4f4921bd5b431|3.39|2014-12-20 11:40:00|1.4102725052409182|3|7203656059|121|0.6186156170875914|0|1|333|-80.995484|52|35.444064|PARMESAN CHEESE|0.0|3|HT GRATED PARMESAN CHEESE|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00072036560599|CHEESE|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|9e63f2171d309a9ccc892ff06b91232229e3a13d|6.99|2014-11-03 13:09:00|1.4102725052409182|3|7203695440|121|0.6186156170875914|0|1|1403|-80.995484|389|35.444064|THAW AND SELL PIES|3.0|14|"8"" SWEET POTATO PIE"|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00072036959362|PIES|BAKERY|-80.995484|1.413637875046387|121|1
35.444064|c9ffe8440c659ccabcfd9f174601e2e5d301ab84|21.45|2014-11-23 10:47:00|1.4102725052409182|3|7343500004|121|0.6186156170875914|0|1|1631|-80.995484|373|35.444064|THAW & SELL (ROLLS)|6.45|14|KING'S HAWAIIAN 12CT ROLLS|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00073435000044|ROLLS|BAKERY|-80.995484|1.413637875046387|121|5
35.444064|6d87e140ef29182189756703822aa92ab0ee3e37|3.99|2014-11-09 08:54:00|1.4102725052409182|3|7203663995|121|0.6186156170875914|0|1|342|-80.995484|57|35.444064|FRESH MILK|1.02|3|HARRIS TEETER 2% MILK|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00072036639981|MILK|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|ee36b3effdaee9b0477b1e88881f5e53657eaeed|5.99|2014-10-07 15:49:00|1.4102725052409182|3|7203695440|121|0.6186156170875914|0|1|1403|-80.995484|389|35.444064|THAW AND SELL PIES|3.0|14|"8"" PUMPKIN PIE"|ead207a0f22b78f0932b76bc180d6ffb6ab10503|0.4616266719835398|0.61833652052202714|00072036954404|PIES|BAKERY|-80.995484|1.413637875046387|121|1
35.444064|d9aadc07d04d32a46cc5f0a06fc10441fc9609a2|8.3|2015-01-31 10:47:00|80.995508130988839|3|4400000488|121|35.44925829308513|0|40|89|-80.8955|12|35.4437|GRAHAM CRACKERS|1.3|1|HONEYMAID GRAHAMFULS S'MORES|ec5d0948adecc063d17f94029ab51776acf1ebf0|0.3589131447681155|35.466476270328783|00044000033972|COOKIES|G1 GROCERY|-80.995484|80.995486869775874|272|2
35.444064|5892c3806da9a303f7f4887f6a1919b6ee91586c|3.79|2015-02-15 10:13:00|1.4102725052409182|3|3890003098|121|0.6186156170875914|0|1|115|-80.995484|16|35.444064|REMAINING FRUIT|1.0|1|DOLE JAR MANDARINS LS|ec5d0948adecc063d17f94029ab51776acf1ebf0|0.3589131447681155|0.61833652052202714|00038900030995|FRUIT-CAN/JAR|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|db65527b02b28485119d734bb21cf48f5cc4f410|2.65|2014-10-12 12:18:00|80.995508130988839|3|4119640471|121|35.44925829308513|0|40|1201|-80.8955|33|35.4437|RTS CANNED|0.65|1|PROG LIGHT BEEF POT ROAST|ec5d0948adecc063d17f94029ab51776acf1ebf0|0.3589131447681155|35.466476270328783|00041196404814|SOUP|G1 GROCERY|-80.995484|80.995486869775874|272|1
35.444064|a52c1aefcb29bb3a906a200ba55d587e062a46a1|3.79|2014-10-20 12:27:00|1.4102725052409182|3|3890003098|121|0.6186156170875914|0|1|115|-80.995484|16|35.444064|REMAINING FRUIT|0.0|1|DOLE JAR MANDARINS LS|ec5d0948adecc063d17f94029ab51776acf1ebf0|0.3589131447681155|0.61833652052202714|00038900030995|FRUIT-CAN/JAR|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|35e163430a8035f3dca347b7b7c4139c72fdf7b4|7.49|2014-12-22 11:10:00|80.995508130988839|3|88133400051|121|35.449258292632756|0|40|36|-80.861571|10|35.444615|PREMIUM GROUND|1.5|1|DUNKIN'D FRENCH VANILLA GROUND|ec5d0948adecc063d17f94029ab51776acf1ebf0|0.3589131447681155|35.466476270328783|00881334000474|COFFEE|G1 GROCERY|-80.995484|80.995487913666338|340|1
35.444064|52d8ab6862c3e41f6a0f6605a17f4a1c91116079|5.05|2015-01-02 10:16:00|1.4102725052409182|3||121|0.6186156170875914|0|1|561|-80.995484|64|35.444064|FR PROD ORGANIC PRODUCE|0.84|4|ORG FUJI APPLES|ec5d0948adecc063d17f94029ab51776acf1ebf0|0.3589131447681155|0.61833652052202714|00294131000002|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|ad1ba0837fac7ff326278346559c6491bc4923f7|1.98|2014-11-30 09:32:00|80.995508130988839|3|7339000780|121|35.449258292632756|0|40|48|-80.861571|7|35.444615|REGISTER GUM|0.2|1|MENTOS MINT ROLL 15CT|ec5d0948adecc063d17f94029ab51776acf1ebf0|0.3589131447681155|35.466476270328783|00073390000110|CANDY|G1 GROCERY|-80.995484|80.995487913666338|340|2
35.444064|397e5705ea9b7bc42da17d5ace4c6232362ec789|3.99|2014-09-15 09:25:00|1.4102725052409182|3|4812121657|121|0.6186156170875914|0|1|1036|-80.995484|164|35.444064|BREAKFAST BAGELS|2.0|7|THOMAS B/S CINN MINI BAGELS PP|ec5d0948adecc063d17f94029ab51776acf1ebf0|0.3589131447681155|0.61833652052202714|00048121216757|BREAKFAST|COMMERCIAL BAKERY|-80.995484|1.413637875046387|121|1
35.444064|f6b6e3c1e93f20a2aef765cb9eab06815ef8cc88|9.99|2014-12-05 18:42:00|80.995508130988839|3|73692011392|121|35.44925829308513|0|40|458|-80.8955|82|35.4437|CRAFT BEER|0.0|16|GOOSE ISLAND SIXTH DAY 6PK|ec5d0948adecc063d17f94029ab51776acf1ebf0|0.3589131447681155|35.466476270328783|00736920113925|DOMESTIC BEER|BEER|-80.995484|80.995486869775874|272|1
35.444064|b7cd2513f0c8cd3c5d4b5bb11514f75472fd045e|4.99|2014-10-28 09:17:00|1.4102725052409182|3|71575620002|121|0.6186156170875914|0|1|504|-80.995484|64|35.444064|FRESH BERRIES|2.5|4|STRAWBERRIES 1LB CLAM|ec5d0948adecc063d17f94029ab51776acf1ebf0|0.3589131447681155|0.61833652052202714|00071430007525|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|e7f437f668a2f6a22003865aac1daa9965739d43|14.99|2014-10-04 18:10:00|1.4102725052409182|3|1820019991|121|0.6186156170875914|0|1|458|-80.995484|82|35.444064|CRAFT BEER|0.0|16|SHOCK TOP SEASONAL 12PK BTL|ec5d0948adecc063d17f94029ab51776acf1ebf0|0.3589131447681155|0.61833652052202714|00018200199912|DOMESTIC BEER|BEER|-80.995484|1.413637875046387|121|1
35.444064|826a9c05a61ba102b7ea90d69756d3aff09cb0e4|2.79|2014-12-16 09:45:00|80.995508130988839|3|1600030140|121|35.449258292632756|0|40|15|-80.861571|2|35.444615|REMAINING BAKING MIXES|0.0|1|BC SUGAR COOKIE MIX|ec5d0948adecc063d17f94029ab51776acf1ebf0|0.3589131447681155|35.466476270328783|00016000306301|BAKING MIXES|G1 GROCERY|-80.995484|80.995487913666338|340|1
35.17335|bbe2559716ffc4ad50feab656109e8e26677a717|11.99|2014-12-07 13:17:00|80.709059419360486|1|20595400000|174|35.192448872290427|0|31|1823|-80.66939|410|35.28326|BH HAM|2.0|6|BOARS HEAD TRIO|ec878eeefb0cc1364593c2ad99a232646c5a7f63|1.3196871103156553|35.187384292804154|00205954000001|BH MEAT|DELI|-80.70901|80.709040945402933|46|1
35.17335|ca6cb023081b22568df244aa558e3df4e833c43a|12.94|2014-11-16 15:23:00|80.709059419360486|1|20254300000|174|35.192448886594086|0|31|299|-80.709466|49|35.124987|ANGUS BEEF|2.2|2|VALUE PK ANGUS STEW MEAT|ec878eeefb0cc1364593c2ad99a232646c5a7f63|1.3196871103156553|35.187384292804154|00202543000008|BEEF|MEAT|-80.70901|80.70902181990985|157|1
35.17335|5a247868e581216c8dcc3b91dc31c6c4adb1203c|4.38|2014-10-05 17:20:00|80.709059419360486|1||174|35.192448872290427|0|31|501|-80.66939|64|35.28326|FRESH PEARS|0.44|4|BARTLETT PEARS|ec878eeefb0cc1364593c2ad99a232646c5a7f63|1.3196871103156553|35.187384292804154|00204409000009|FRESH PRODUCE|PRODUCE|-80.70901|80.709040945402933|46|1
35.17335|c4208daaa4b8f16a4c78be40b398ea2c9014f9f9|5.53|2014-09-28 15:44:00|80.709059419360486|1||174|35.192448872290427|0|31|501|-80.66939|64|35.28326|FRESH PEARS|0.83|4|BARTLETT PEARS|ec878eeefb0cc1364593c2ad99a232646c5a7f63|1.3196871103156553|35.187384292804154|00204409000009|FRESH PRODUCE|PRODUCE|-80.70901|80.709040945402933|46|1
35.17335|4718b80ddf68ce5760c7fd185bdbcf933ff22b0f|8.79|2015-01-03 14:20:00|80.709059419360486|1|9955508520|174|35.192448886594086|0|31|37|-80.709466|10|35.124987|PODS/CUPS/SINGLES|1.8|1|GREEN MTN K-CUPS HALF CAFF|ec878eeefb0cc1364593c2ad99a232646c5a7f63|1.3196871103156553|35.187384292804154|00099555089998|COFFEE|G1 GROCERY|-80.70901|80.70902181990985|157|1
35.17335|fed9c43b2d722c759a131b828e7ab045a387588a|3.99|2015-03-07 15:39:00|80.709059419360486|1|7203602701|174|35.192448886594086|0|31|1878|-80.709466|435|35.124987|HUMMUS|0.3|6|FFM ARTISAN RED PEPPER HUMMUS|ec878eeefb0cc1364593c2ad99a232646c5a7f63|1.3196871103156553|35.187384292804154|00072036027030|SALADS|DELI|-80.70901|80.70902181990985|157|1
35.17335|de7d4d03a7656682e60d46c39cdb4804c34a8f56|39.4|2014-11-08 13:32:00|80.709059419360486|1|20129900000|174|35.192448886594086|0|31|296|-80.709466|49|35.124987|RANCHER BEEF|0.0|2|VALUE PK BEEF LOIN STRIP STEAK|ec878eeefb0cc1364593c2ad99a232646c5a7f63|1.3196871103156553|35.187384292804154|00201299000003|BEEF|MEAT|-80.70901|80.70902181990985|157|2
35.17335|e0376540485bfc8c58103c7bb678b9e0390bbd67|2.99|2014-09-20 12:05:00|80.709059419360486|1|1600081341|174|35.192448886594086|0|31|8|-80.709466|2|35.124987|BROWNIE MIXES|0.99|1|BC SUP/HERSHEY ULTIMATE FUDGE|ec878eeefb0cc1364593c2ad99a232646c5a7f63|1.3196871103156553|35.187384292804154|00016000813397|BAKING MIXES|G1 GROCERY|-80.70901|80.70902181990985|157|1
35.17335|f472df42c65f1a1018650c62508b91400b581983|4.29|2014-10-25 13:42:00|80.709059419360486|1|2840016014|174|35.192448886594086|0|31|201|-80.709466|31|35.124987|POTATO CHIPS|2.15|1|LAYS WAVY REGULAR|ec878eeefb0cc1364593c2ad99a232646c5a7f63|1.3196871103156553|35.187384292804154|00028400160209|SNACKS|G1 GROCERY|-80.70901|80.70902181990985|157|1
35.17335|f45bc6c86803241388032e458cc5db3b583fc1c3|4.29|2014-10-11 16:58:00|80.709059419360486|1|2840016014|174|35.192448886594086|0|31|201|-80.709466|31|35.124987|POTATO CHIPS|0.29|1|LAYS WAVY REGULAR|ec878eeefb0cc1364593c2ad99a232646c5a7f63|1.3196871103156553|35.187384292804154|00028400160209|SNACKS|G1 GROCERY|-80.70901|80.70902181990985|157|1
35.17335|d2f9120657f240fd9ec7d1835899f55635986ed1|2.99|2014-11-08 13:37:00|80.709059419360486|1|3338365583|174|35.192448886594086|0|31|522|-80.709466|64|35.124987|FRESH TOMATOES|0.2|4|SWEET GRAPE TOMATO (PINT)|ec878eeefb0cc1364593c2ad99a232646c5a7f63|1.3196871103156553|35.187384292804154|00072036880284|FRESH PRODUCE|PRODUCE|-80.70901|80.70902181990985|157|1
35.17335|3a2b79b05a696c2172cce8dc3c7f0f3e58985b7a|13.99|2014-09-24 14:20:00|80.709059419360486|1|7203695696|174|35.192448888613562|0|31|1653|-80.661096|381|35.172688|CELEBRATION CAKES|0.0|14|1/8 SHEET DL MBL W/WHT BUTCRM|ec878eeefb0cc1364593c2ad99a232646c5a7f63|1.3196871103156553|35.187384292804154|00072036956965|CAKES|BAKERY|-80.70901|80.709014922746533|474|1
35.17335|d486a45d77c0e76995c0535256f325e8116920c4|5.29|2014-11-03 13:33:00|80.709059419360486|1|5150024177|174|35.192448888171036|0|31|125|-80.826724|19|35.195689|PEANUT BUTTER|1.3|1|JIF CREAMY PEANUT BUTTER|ec878eeefb0cc1364593c2ad99a232646c5a7f63|1.3196871103156553|35.187384292804154|00051500241776|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.70901|80.70901703831629|412|1
35.17335|b8567419444ecf5cadf5ab560cd0ddf10a096613|4.99|2015-02-24 15:40:00|80.709059419360486|1|5000034934|174|35.192448876610591|0|31|144|-80.78468|229|35.096737|CEAMERS-POWDERED|0.0|1|COFFEE MATE HAZELNUT SUGAR FRE|ec878eeefb0cc1364593c2ad99a232646c5a7f63|1.3196871103156553|35.187384292804154|00050000349340|COCOAS CREAMERS SYRUPS|G1 GROCERY|-80.70901|80.709036656775623|30|1
35.17335|39cdd23cad7020b0e42cadd941b74aef11296d05|7.99|2015-02-14 12:32:00|80.709059419360486|1|8500001845|174|35.192448886594086|0|31|9939|-80.709466|885|35.124987|NFS POP PINOT NOIR|0.0|13|THE NAKED GRAPE PINOT NOIR|ec878eeefb0cc1364593c2ad99a232646c5a7f63|1.3196871103156553|35.187384292804154|00085000018453|POPULAR (4-$7.99)|WINE|-80.70901|80.70902181990985|157|1
35.17335|4b9a13471a3065d366677e8c67459453ca372018|8.49|2015-02-22 13:12:00|80.709059419360486|1|78260516150|174|35.192448888613562|0|31|37|-80.661096|10|35.172688|PODS/CUPS/SINGLES|2.5|1|KAUAI K-CUP ISLAND SUNRSE MILD|ec878eeefb0cc1364593c2ad99a232646c5a7f63|1.3196871103156553|35.187384292804154|00782605161514|COFFEE|G1 GROCERY|-80.70901|80.709014922746533|474|1
35.140781|0c6d3a091331081615c3af8c93cb19d682739f00|40.98|2014-11-14 14:34:00|80.632521683083056|4|7023666338|39|35.170088500729086|0|39|751|-80.661096|87|35.172688|NFS-BOUQUETS|0.0|9|$19.99 EN VOUGUE|f21e95851758cb8f74a95d0c0c0442303d8c9afd|2.0250775514967287|35.177497916598789|00070236663386|FLORAL|FLORAL|-80.62331|80.62331576583513|474|2
35.140781|13a0742e57b482bcf0a70ab15ee40d92a485d600|2.99|2015-01-15 18:44:00|1.4091206135396188|4|3120020007|39|0.6133223301722653|0|47|130|-80.62331|20|35.140781|CRANBERRY JUICE/DRINKS-SHELF|0.0|1|OSPRAY CRAN LEMONADE|f21e95851758cb8f74a95d0c0c0442303d8c9afd|2.0250775514967287|0.61242566243833529|00031200201676|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.62331|1.4071422133560694|39|1
35.140781|632b78f0a2dbe27de4d93179f77d25fe6408a330|18.99|2015-02-14 09:06:00|1.4091206135396188|4|20496100000|39|0.6133223301722653|0|47|754|-80.62331|87|35.140781|NFS-SGLE STEM CUT FLOWER|0.0|9|*SINGLE STEM CUT FLOWERS|f21e95851758cb8f74a95d0c0c0442303d8c9afd|2.0250775514967287|0.61242566243833529|00204961000004|FLORAL|FLORAL|-80.62331|1.4071422133560694|39|1
35.140781|f213ad85110b2d33e7c966e14f5262a5b2afecab|2.0|2015-02-06 18:09:00|1.4091206135396188|4|7203663159|39|0.6133223301722653|0|47|1134|-80.62331|57|35.140781|CARTON MILK|0.0|3|HARRIS TEETER CHOCOLATE MILK|f21e95851758cb8f74a95d0c0c0442303d8c9afd|2.0250775514967287|0.61242566243833529|00072036631596|MILK|DAIRY|-80.62331|1.4071422133560694|39|1
35.140781|00e0f82844f6e7c6d26b7f8e6b2cb0f41b3b671d|4.15|2014-09-14 19:55:00|1.4091206135396188|4|7203670344|39|0.6133223301722653|0|47|443|-80.62331|76|35.140781|NFS-GARBAGE BAGS|0.0|1|YH CLR LAWN N LEAF BAGS|f21e95851758cb8f74a95d0c0c0442303d8c9afd|2.0250775514967287|0.61242566243833529|00072036703514|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.62331|1.4071422133560694|39|1
35.152722|38d3e23d387274e81cb8694980ec4812d9714cca|28.49|2014-09-28 03:23:00|80.825044058860698|4|3700086268|160|35.154107980622896|0|29|1206|-80.737839|67|35.297134|NFS-BOX DIAPERS|2.5|1|PAMP CRUISER SUPER PACK SIZE 6|f29a1bfdae0ca2588dd93160ad423aaa4208a94b|0.09576808655544278|35.157881615307893|00037000862710|DISPOSABLE DIAPERS|G1 GROCERY|-80.825175|80.825178217761746|258|1
35.152722|63ed044a00b31c6a91a40f3d02557c3df75fa771|53.98|2014-12-09 14:53:00|80.825044058860698|4|3700086268|160|35.154107980622896|0|29|1206|-80.737839|67|35.297134|NFS-BOX DIAPERS|4.0|1|PAMP CRUISER SUPER PACK SIZE 6|f29a1bfdae0ca2588dd93160ad423aaa4208a94b|0.09576808655544278|35.157881615307893|00037000862710|DISPOSABLE DIAPERS|G1 GROCERY|-80.825175|80.825178217761746|258|2
35.152722|ec43a581eff0e715f3470efd256ba671a910b41c|2.39|2014-10-28 18:22:00|80.825044058860698|4|3760048669|160|35.154107980622896|0|29|362|-80.737839|102|35.297134|PEPPERONIS|0.0|19|HORMEL SLICED PEPPERONI|f29a1bfdae0ca2588dd93160ad423aaa4208a94b|0.09576808655544278|35.157881615307893|00037600486699|LUNCHMEATS|CASE READY MEATS|-80.825175|80.825178217761746|258|1
35.152722|85ebdfdefe34a15febad6362bddc4da5e6dffa08|10.99|2014-10-20 20:06:00|80.825044058860698|4|3700086258|160|35.154107980622896|0|29|1205|-80.737839|67|35.297134|NFS-JUMBO DIAPERS|1.0|1|PAMPERS CRUISERS JUMBO SIZE 6|f29a1bfdae0ca2588dd93160ad423aaa4208a94b|0.09576808655544278|35.157881615307893|00037000862611|DISPOSABLE DIAPERS|G1 GROCERY|-80.825175|80.825178217761746|258|1
35.152722|25d11bb8d19dc8c1ab87d8337092bfcfed9203d9|3.39|2015-02-25 21:01:00|80.825044058860698|4|3800031829|160|35.154107980622896|0|29|74|-80.737839|9|35.297134|RTE CEREAL ALL FAMILY|0.89|1|KELL MIN WH LIL BITES ORIG|f29a1bfdae0ca2588dd93160ad423aaa4208a94b|0.09576808655544278|35.157881615307893|00038000596827|CEREAL|G1 GROCERY|-80.825175|80.825178217761746|258|1
35.152722|39e2a33be907b05e76b0341490a987410e6f1e75|19.95|2015-02-04 18:05:00|80.825044058860698|4|20931900000|160|35.154107980622896|0|29|676|-80.737839|148|35.297134|TAILS|0.0|12|WC LOBSTER TAILS 2/3 OZ  (CA)|f29a1bfdae0ca2588dd93160ad423aaa4208a94b|0.09576808655544278|35.157881615307893|00209319000002|LOBSTERS|SEAFOOD|-80.825175|80.825178217761746|258|1
35.152722|3d7e3a42ab4bee147b5122f543b1e08fdc763c7a|4.29|2015-01-11 21:15:00|80.825044058860698|4|2840015938|160|35.154107980622896|0|29|201|-80.737839|31|35.297134|POTATO CHIPS|2.15|1|RUFFLES REGULAR|f29a1bfdae0ca2588dd93160ad423aaa4208a94b|0.09576808655544278|35.157881615307893|00028400159388|SNACKS|G1 GROCERY|-80.825175|80.825178217761746|258|1
35.152722|2ee141b2fbb1fe59042c976e26434115fbf0eaf8|6.99|2015-02-20 15:42:00|80.825044058860698|4|4900002890|160|35.154107980622896|0|29|55|-80.737839|8|35.297134|REGULAR|3.5|23|SPRITE 12OZ 12PK FRIDGE CAN|f29a1bfdae0ca2588dd93160ad423aaa4208a94b|0.09576808655544278|35.157881615307893|00049000028928|CARBONATED BEVERAGES|BEVERAGE|-80.825175|80.825178217761746|258|1
35.152722|209b4b273fcb1fc0150a18e37dd84f972bfd73b9|3.99|2015-03-03 21:01:00|80.825044058860698|4|7660660269|160|35.154107980622896|0|29|208|-80.737839|32|35.297134|NFS-COCKTAIL ACCESSORIES|0.0|1|HH MARASCHINO CHERRY|f29a1bfdae0ca2588dd93160ad423aaa4208a94b|0.09576808655544278|35.157881615307893|00076606602696|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.825175|80.825178217761746|258|1
35.152722|b45be9c4c3e38e36cefa9b97b531c9811e740731|3.69|2015-02-24 17:14:00|80.825044058860698|4|2500005542|160|35.154107980622896|0|29|335|-80.737839|56|35.297134|ORANGE JUICE-REGRIGERATED|0.0|3|SIMPLY ORANGE ORIGINAL|f29a1bfdae0ca2588dd93160ad423aaa4208a94b|0.09576808655544278|35.157881615307893|00025000055423|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.825175|80.825178217761746|258|1
35.152722|faa39e85fc13ed5a65d38013b3ce99c106bd7afb|0.92|2014-11-13 19:56:00|80.825044058860698|4||160|35.154107980622896|0|29|524|-80.737839|64|35.297134|FRESH PROD FRESH ONIONS|0.0|4|COO YELLOW ONIONS, LRG|f29a1bfdae0ca2588dd93160ad423aaa4208a94b|0.09576808655544278|35.157881615307893|00204665000003|FRESH PRODUCE|PRODUCE|-80.825175|80.825178217761746|258|1
35.152722|8517fed0a6668ec6c23bf46751a05725deb6efa2|14.940000000000001|2015-02-21 21:45:00|80.825044058860698|4|60888300005|160|35.154107980622896|0|29|31|-80.737839|4|35.297134|NON CARBONATED WATER|1.25|1|ETERNAL ARTISIAN WATER 1 LITER|f29a1bfdae0ca2588dd93160ad423aaa4208a94b|0.09576808655544278|35.157881615307893|00608883000058|BOTTLED WATER|G1 GROCERY|-80.825175|80.825178217761746|258|6
35.152722|fae124a6388be47edd5975d3c848cf0c5b8ac7a6|37.91|2014-12-24 18:16:00|80.825044058860698|4|20896300000|160|35.154107980622896|0|29|977|-80.737839|201|35.297134|FRESH HT CHICKEN|3.69|2|HT VALUE PK CHICKEN WINGS|f29a1bfdae0ca2588dd93160ad423aaa4208a94b|0.09576808655544278|35.157881615307893|00208963000000|POULTRY|MEAT|-80.825175|80.825178217761746|258|3
35.152722|8af259b9b0bfc0e9b16b1509c1ad36068b0d7f53|1.29|2015-01-21 21:58:00|80.825044058860698|4|7097000002|160|35.154107980622896|0|29|727|-80.737839|7|35.297134|SEASONAL CANDY-SINGLE FAC|0.65|1|I/O(V15)PEEPS CHICKS YELLW 5CT|f29a1bfdae0ca2588dd93160ad423aaa4208a94b|0.09576808655544278|35.157881615307893|00070970000027|CANDY|G1 GROCERY|-80.825175|80.825178217761746|258|1
35.152722|c5a986a0710b101d3006e0ca80ec1322fd543deb|8.99|2014-09-28 03:24:00|80.825044058860698|4|87126011085|160|35.154107980622896|0|29|740|-80.737839|87|35.297134|NFS-ROSE BQT|0.0|9|BUNCH- 10 CONSUMER ROSE|f29a1bfdae0ca2588dd93160ad423aaa4208a94b|0.09576808655544278|35.157881615307893|00871260110859|FLORAL|FLORAL|-80.825175|80.825178217761746|258|1
35.152722|658a5606b24ea264e9098e2019cb3151c7037992|5.38|2015-02-11 18:51:00|80.825044058860698|4|1450000253|160|35.154107980622896|0|29|1272|-80.737839|50|35.297134|BAG VEG STEAM|0.69|5|BE STEAMFRESH PREM BROCC FLRTS|f29a1bfdae0ca2588dd93160ad423aaa4208a94b|0.09576808655544278|35.157881615307893|00014500011831|VEGETABLES-FROZEN|FROZEN|-80.825175|80.825178217761746|258|2
35.152722|bdfd75c075f29493ea6ec7cb5dff0a9feab62063|9.99|2014-11-12 17:41:00|80.825044058860698|4|6574311308|160|35.154107980622896|0|29|3476|-80.737839|1040|35.297134|BRAND-PAUL MITCHELL|0.0|17|PAUL MITCHELL SHAMPOO 1|f29a1bfdae0ca2588dd93160ad423aaa4208a94b|0.09576808655544278|35.157881615307893|00065743113080|PROFESSIONAL HAIR & SCALP CARE|HBC|-80.825175|80.825178217761746|258|1
35.152722|4b2e1e9f4a7abc065bc524706744117d0833a57a|3.69|2014-10-20 20:08:00|80.825044058860698|4|1620033700|160|35.154107980622896|0|29|225|-80.737839|35|35.297134|SUGAR-GRANULATED|1.2|1|DIXIE CRYSTAL 4 LB GRAN SUGAR|f29a1bfdae0ca2588dd93160ad423aaa4208a94b|0.09576808655544278|35.157881615307893|00016200337006|SUGAR/SUBSTITUTES|G1 GROCERY|-80.825175|80.825178217761746|258|1
35.061685|eb115306df6ac7ab8b727f3d806476bd3821093d|5.99|2014-09-17 18:01:00|80.994598860450068|2|7732661225|475|35.071208776812753|0|53|3878|-80.97058|1070|35.03469|SOLID-UNISEX|2.49|17|TOM APRICOT LL DEOD STK|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00077326611258|DEODORANT|HBC|-80.994596|80.994598009133426|82|1
35.061685|457f4ae9c08847fc02cb8a955abb72e2cd880a2b|9.99|2015-02-02 08:39:00|80.994598860450068|2|9955536128|475|35.071208776812753|0|53|35|-80.97058|10|35.03469|PREMIUM WHOLE BEAN|0.0|1|NEWMAN'S ORG/COLOMBIAN W/B|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00099555361285|COFFEE|G1 GROCERY|-80.994596|80.994598009133426|82|1
35.061685|b83735f40acdc6e974bb1c4bc66976a60c4edaa3|5.15|2014-11-20 13:50:00|80.994598860450068|2||475|35.071208776812753|0|53|561|-80.97058|64|35.03469|FR PROD ORGANIC PRODUCE|1.44|4|ORG SWEET POTATOES|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00294091000005|FRESH PRODUCE|PRODUCE|-80.994596|80.994598009133426|82|1
35.061685|d217e3109200ee4f9c6ed18e05229700e3b72cc7|9.99|2014-11-26 14:36:00|1.4132775322775095|2|75122802115|475|0.611941844547108|0|58|36|-80.994596|10|35.061685|PREMIUM GROUND|2.0|1|ORGANIC COFFEE JAVA LOVE|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|0.61177642288969325|00751228552030|COFFEE|G1 GROCERY|-80.994596|1.4136223765226292|475|1
35.061685|68bcfcd5641b7ab7330e967d660ffc86af9df087|2.99|2015-03-03 16:24:00|80.994598860450068|2|20443000000|475|35.071208776812753|0|53|510|-80.97058|64|35.03469|FRESH PINEAPPLE|0.0|4|GOLD PINEAPPLES|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00643126072003|FRESH PRODUCE|PRODUCE|-80.994596|80.994598009133426|82|1
35.061685|9736a05a9265f036a10fe67aac2e872c980337ce|2.99|2014-12-11 13:02:00|80.994598860450068|2|20443000000|475|35.071208776812753|0|53|510|-80.97058|64|35.03469|FRESH PINEAPPLE|0.0|4|GOLD PINEAPPLES|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00643126072003|FRESH PRODUCE|PRODUCE|-80.994596|80.994598009133426|82|1
35.061685|a21cbbd6b54a0f8a199b8a2a330b608f5548ad84|9.99|2015-01-19 16:45:00|1.4132775322775095|2|75122802115|475|0.611941844547108|0|58|36|-80.994596|10|35.061685|PREMIUM GROUND|2.0|1|ORGANIC COFFEE JAVA LOVE|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|0.61177642288969325|00751228552030|COFFEE|G1 GROCERY|-80.994596|1.4136223765226292|475|1
35.061685|a4e31853f71460895a7a0295c60a1e041c53d415|2.25|2014-09-25 18:09:00|80.994598860450068|2||475|35.071208776812753|0|53|561|-80.97058|64|35.03469|FR PROD ORGANIC PRODUCE|0.23|4|ORG SWEET POTATOES|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00294091000005|FRESH PRODUCE|PRODUCE|-80.994596|80.994598009133426|82|1
35.061685|0ef77b089e34b24558af0efa3cd3b50c9174b9ab|3.56|2015-02-09 08:57:00|80.994598860450068|2||475|35.071208776812753|0|53|561|-80.97058|64|35.03469|FR PROD ORGANIC PRODUCE|0.0|4|ORG SWEET POTATOES|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00294091000005|FRESH PRODUCE|PRODUCE|-80.994596|80.994598009133426|82|1
35.061685|d3c17ba38f0bcce8048d82d17c8231e6949adb14|3.99|2015-01-25 18:31:00|1.4132775322775095|2||475|0.611941844547108|0|58|561|-80.994596|64|35.061685|FR PROD ORGANIC PRODUCE|0.0|4|ORG CAULIFLOWER|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|0.61177642288969325|00294079000003|FRESH PRODUCE|PRODUCE|-80.994596|1.4136223765226292|475|1
35.061685|feb48f8100c6c0d1f14acac07963291f910185a8|2.49|2015-01-26 09:07:00|80.994598860450068|2|72722322247|475|35.071208776812753|0|53|6987|-80.97058|1600|35.03469|VALENTINE HOME DECOR-IMPORT|0.0|18|I/O VAL GEL CLING ASSORTMENT|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00727223222476|SEASONAL MERCHANDISE|GM|-80.994596|80.994598009133426|82|1
35.061685|2ecec0e3589b0a325f5856fc509ad042915dde56|3.99|2014-11-13 20:10:00|80.994598860450068|2||475|35.071208776812753|0|53|561|-80.97058|64|35.03469|FR PROD ORGANIC PRODUCE|0.0|4|ORG CAULIFLOWER|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00294079000003|FRESH PRODUCE|PRODUCE|-80.994596|80.994598009133426|82|1
35.061685|ec2d5dfe3768e608b8d0be2de0b3e7a919801793|3.11|2015-02-14 19:10:00|1.4132775322775095|2||475|0.611941844547108|0|58|561|-80.994596|64|35.061685|FR PROD ORGANIC PRODUCE|0.0|4|ORG SWEET POTATOES|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|0.61177642288969325|00294091000005|FRESH PRODUCE|PRODUCE|-80.994596|1.4136223765226292|475|1
35.061685|c0113435de5430abc2d062b858463fad08454cd7|3.54|2014-10-25 19:37:00|80.994598860450068|2||475|35.071208776812753|0|53|561|-80.97058|64|35.03469|FR PROD ORGANIC PRODUCE|0.0|4|ORG SWEET POTATOES|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00294091000005|FRESH PRODUCE|PRODUCE|-80.994596|80.994598009133426|82|1
35.061685|0494ea066a982b7f56573c42ad8cb5b982191dc5|4.91|2015-02-17 17:46:00|80.994598860450068|2||475|35.071208776812753|0|53|561|-80.97058|64|35.03469|FR PROD ORGANIC PRODUCE|0.0|4|ORG SWEET POTATOES|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00294091000005|FRESH PRODUCE|PRODUCE|-80.994596|80.994598009133426|82|1
35.061685|b23094bdb3601a69c07330080983f7986d47bc50|3.39|2014-10-15 16:48:00|1.4132775322775095|2||475|0.611941844547108|0|58|561|-80.994596|64|35.061685|FR PROD ORGANIC PRODUCE|0.0|4|ORG SWEET POTATOES|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|0.61177642288969325|00294091000005|FRESH PRODUCE|PRODUCE|-80.994596|1.4136223765226292|475|1
35.061685|e50bfda69943e46797561069dfd8aaff9cf001b5|14.38|2015-02-06 09:07:00|80.994598860450068|2|3760035160|475|35.071208776812753|0|53|845|-80.97058|100|35.03469|NATURAL/ORGANIC BACON|3.6|19|HORMEL NATURAL CHOICE BACON|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00037600445955|BACON|CASE READY MEATS|-80.994596|80.994598009133426|82|2
35.061685|3fe4702ee153253db514a6dda3c42bb46621c0ba|7.99|2014-11-08 17:00:00|80.994598860450068|2|3760035160|475|35.071208776812753|0|53|845|-80.97058|100|35.03469|NATURAL/ORGANIC BACON|3.49|19|HORMEL NATURAL CHOICE BACON|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00037600445955|BACON|CASE READY MEATS|-80.994596|80.994598009133426|82|1
35.061685|ef90cbc87aba4443dc809c1bf849f4b0e0a6ccfd|1.49|2015-02-23 08:46:00|80.994598860450068|2|4113700761|475|35.071208776812753|0|53|387|-80.97058|65|35.03469|NFS-REMAIN CHAR/LOGS/ACC|0.0|1|"DURAFLAME 1"" MATCHES"|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00041137007616|CHARCOAL/LOGS/ACCESSORIES|G1 GROCERY|-80.994596|80.994598009133426|82|1
35.061685|ea10817f791831ddfdf22148b95b30cf50eda6bd|9.57|2014-10-12 19:13:00|80.994598860450068|2|75764561250|475|35.071208776812753|0|53|158|-80.97058|24|35.03469|NFS-DOG FOOD-WET|0.69|1|NEWMAN ORG DOG CHICKEN DINNER.|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00757645612500|PET FOOD/SUPPLIES|G1 GROCERY|-80.994596|80.994598009133426|82|3
35.061685|d751de1813c78a0fa49ae32637efca259f2c290d|6.38|2014-10-04 19:32:00|80.994598860450068|2|75764561250|475|35.071208776812753|0|53|158|-80.97058|24|35.03469|NFS-DOG FOOD-WET|0.69|1|NEWMAN ORG DOG CHICKEN DINNER.|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00757645612500|PET FOOD/SUPPLIES|G1 GROCERY|-80.994596|80.994598009133426|82|2
35.061685|1aa0db87c4f5c3315f0717a936d1bd4dc540e225|2.79|2014-12-16 16:21:00|1.4132775322775095|2|75764561250|475|0.611941844547108|0|58|158|-80.994596|24|35.061685|NFS-DOG FOOD-WET|0.0|1|NEWMAN ORG DOG CHICKEN DINNER.|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|0.61177642288969325|00757645612500|PET FOOD/SUPPLIES|G1 GROCERY|-80.994596|1.4136223765226292|475|1
35.061685|68a13c52c34d135f0017f5806f20ee95bf0b3c2d|8.370000000000001|2014-09-15 17:46:00|80.994598860450068|2|75764561200|475|35.071208776812753|0|53|158|-80.97058|24|35.03469|NFS-DOG FOOD-WET|0.79|1|NEWMAN ORG CAN DOG CH&BRWN RC|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00757645612005|PET FOOD/SUPPLIES|G1 GROCERY|-80.994596|80.994598009133426|82|3
35.061685|a14bfc377b7d0d26506c64b9c1e4d4fb134b7568|2.79|2015-01-04 18:05:00|80.994598860450068|2|75764561250|475|35.071208776812753|0|53|158|-80.97058|24|35.03469|NFS-DOG FOOD-WET|0.0|1|NEWMAN ORG DOG CHICKEN DINNER.|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00757645612500|PET FOOD/SUPPLIES|G1 GROCERY|-80.994596|80.994598009133426|82|1
35.061685|cc90c8b95ef53f8fe9b8894f5bf679ae71121122|11.16|2014-09-22 18:31:00|80.994598860450068|2|75764561200|475|35.071208776812753|0|53|158|-80.97058|24|35.03469|NFS-DOG FOOD-WET|3.16|1|NEWMAN ORG CAN DOG CH&BRWN RC|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00757645612005|PET FOOD/SUPPLIES|G1 GROCERY|-80.994596|80.994598009133426|82|4
35.061685|6adb3dc5c7f506125461dcf92da9d6fe3555f0b7|2.79|2014-12-29 12:54:00|80.994598860450068|2|75764561250|475|35.071208776812753|0|53|158|-80.97058|24|35.03469|NFS-DOG FOOD-WET|0.0|1|NEWMAN ORG DOG CHICKEN DINNER.|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00757645612500|PET FOOD/SUPPLIES|G1 GROCERY|-80.994596|80.994598009133426|82|1
35.061685|b53adecbd9b81198b9222b07e7c9dca99687fbf0|2.79|2015-03-09 08:34:00|80.994598860450068|2|75764561250|475|35.071208776812753|0|53|158|-80.97058|24|35.03469|NFS-DOG FOOD-WET|0.0|1|NEWMAN ORG DOG CHICKEN DINNER.|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00757645612500|PET FOOD/SUPPLIES|G1 GROCERY|-80.994596|80.994598009133426|82|1
35.061685|c095f23539669e48b1bb235b437af28dc216cab9|2.49|2014-09-12 13:57:00|80.994598860450068|2|7203698227|475|35.071208776812753|0|53|126|-80.97058|19|35.03469|PRESERVES/MARMALADE|0.0|1|HTO PRES APRICOT|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00072036982469|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.994596|80.994598009133426|82|1
35.061685|d7a873d9952d46c66e74f812f7b90bb8fac7bb70|5.0|2014-12-22 12:45:00|80.994598860450068|2|7203676367|475|35.071208776812753|0|53|243|-80.97058|39|35.03469|BAKED BEANS|0.0|1|HTO BAKED BEAN MAPLE|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00072036763679|VEGETABLES-CAN/JAR|G1 GROCERY|-80.994596|80.994598009133426|82|3
35.061685|80c1b9c3a29ce6edbeb61c0da1b0a07e1902c89e|2.99|2014-12-24 13:31:00|80.994598860450068|2|4667710630|475|35.071208776812753|0|53|6139|-80.97058|1546|35.03469|BULB-CARD NIGHT LIGHTS|0.0|18|(FE)(JHK)PHILIP 4W BC CLR S|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00046677106300|LIGHT BULBS/ELECTRICAL|GM|-80.994596|80.994598009133426|82|1
35.061685|60e919e433ee8336b8982f987c8c14a84075d2e4|2.29|2014-10-27 16:12:00|80.994598860450068|2|4150880012|475|35.071208776812753|0|53|30|-80.97058|4|35.03469|CARBONATED WATER|0.4|1|SAN PELLEGRINO 750ML|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00041508800129|BOTTLED WATER|G1 GROCERY|-80.994596|80.994598009133426|82|1
35.061685|b4ef5c04dbb2c26815c7f9e3628867978281d212|4.98|2015-01-28 09:22:00|80.994598860450068|2|4150880012|475|35.071208776812753|0|53|30|-80.97058|4|35.03469|CARBONATED WATER|0.49|1|SAN PELLEGRINO 750ML|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00041508800129|BOTTLED WATER|G1 GROCERY|-80.994596|80.994598009133426|82|2
35.061685|318e88b25386b3ef264906dde52578efae5d017c|2.49|2015-01-08 18:31:00|80.994598860450068|2|4150880012|475|35.071208776812753|0|53|30|-80.97058|4|35.03469|CARBONATED WATER|0.49|1|SAN PELLEGRINO 750ML|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00041508800129|BOTTLED WATER|G1 GROCERY|-80.994596|80.994598009133426|82|1
35.061685|7d526bba99c7e2249345ea6635807f31109eed84|17.49|2015-02-24 08:55:00|80.994598860450068|2|75764566010|475|35.071208776812753|0|53|156|-80.97058|24|35.03469|NFS-DOG FOOD-DRY|0.0|1|NEWMAN ORG ADLT DOG CHK RC DRY|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00757645660105|PET FOOD/SUPPLIES|G1 GROCERY|-80.994596|80.994598009133426|82|1
35.061685|f16c285ccb19a98fc707fad9c6d53e74f2ace16d|12.57|2014-10-22 20:18:00|80.994598860450068|2|74236531660|475|35.071208776812753|0|53|322|-80.97058|53|35.03469|SOUR CREAM|3.57|3|HORIZON SOUR CREAM 16 OZ|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00742365316609|CULTURES|DAIRY|-80.994596|80.994598009133426|82|3
35.061685|12a7d92f4e91364f5ea343cd7554b358f9417060|4.19|2014-09-30 17:19:00|80.994598860450068|2|74236531660|475|35.071208776812753|0|53|322|-80.97058|53|35.03469|SOUR CREAM|0.0|3|HORIZON SOUR CREAM 16 OZ|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00742365316609|CULTURES|DAIRY|-80.994596|80.994598009133426|82|1
35.061685|4b2a238bb4f6bfdff8ad0192c7353bb9a7b9f20a|3.29|2015-03-04 14:55:00|1.4132775322775095|2|65724350106|475|0.611941844547108|0|58|273|-80.994596|43|35.061685|PREMIUM NOVELTIES|0.0|5|PS CHOC FRUIT DIP BANANA|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|0.61177642288969325|00657243502060|FROZEN NOVELTIES|FROZEN|-80.994596|1.4136223765226292|475|1
35.061685|46f9b98e96026cb745ba13bd30d9ea193817b802|1.99|2015-01-15 19:03:00|80.994598860450068|2||475|35.071208776812753|0|53|561|-80.97058|64|35.03469|FR PROD ORGANIC PRODUCE|0.0|4|COO ORG RUSSET POTATO 50/60CT|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00294072000000|FRESH PRODUCE|PRODUCE|-80.994596|80.994598009133426|82|1
35.061685|4e1d587cbbe53535467aa925ea74afd7e30324d4|4.58|2014-12-05 13:38:00|80.994598860450068|2|7203676383|475|35.071208776812753|0|53|225|-80.97058|35|35.03469|SUGAR-GRANULATED|0.58|1|HTN ORGANIC SUGAR FT|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00072036763839|SUGAR/SUBSTITUTES|G1 GROCERY|-80.994596|80.994598009133426|82|2
35.061685|d99b29cc7ece47fe9fc545acd81b708a159312f6|4.59|2015-01-23 11:18:00|1.4132775322775095|2|5385200220|475|0.611941844547108|0|58|204|-80.994596|31|35.061685|TORTILLA CHIPS|0.6|1|GREEN MTN GRINGO WHITE TORTLLA|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|0.61177642288969325|00053852002203|SNACKS|G1 GROCERY|-80.994596|1.4136223765226292|475|1
35.061685|ac8fb9eb3060d689b3a53edf8389416616362885|2.49|2014-11-29 18:02:00|80.994598860450068|2||475|35.071208776812753|0|53|561|-80.97058|64|35.03469|FR PROD ORGANIC PRODUCE|0.0|4|ORG HASS AVOCADOS|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00294225000000|FRESH PRODUCE|PRODUCE|-80.994596|80.994598009133426|82|1
35.061685|7e84d29d751bc11b32f32adbfafb21e67f113efb|1.69|2014-11-21 18:47:00|80.994598860450068|2|7203698517|475|35.071208776812753|0|53|426|-80.97058|72|35.03469|NFS-PAPER TOWELS|0.35|1|YH ULT TOWEL 1RL SAS|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00072036985170|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.994596|80.994598009133426|82|1
35.061685|52996b1544e0441b5dd44c7231e21b5d0f50b7bd|4.99|2014-10-18 17:55:00|80.994598860450068|2|2840016473|475|35.071208776812753|0|53|201|-80.97058|31|35.03469|POTATO CHIPS|1.0|1|LAYS CLASSIC PARTY SIZE|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|35.072594466811061|00028400164733|SNACKS|G1 GROCERY|-80.994596|80.994598009133426|82|1
35.061685|f9d5b9f5d679331b49797948df0db6aeb1d0df6c|1.29|2015-03-08 21:19:00|1.4132775322775095|2|7203678692|475|0.611941844547108|0|58|1208|-80.994596|23|35.061685|WHSE PASTA VALUE ADD|0.0|1|HTO SPAGHETTI.|fb39e75903b150547e2f702dc4b0d40544d3d5fc|0.6580699884734476|0.61177642288969325|00072036707130|PASTA|G1 GROCERY|-80.994596|1.4136223765226292|475|1
35.006282|6adebd1a3c8ae9eb61b4597310306d9647788945|2.77|2014-09-12 13:38:00|1.4091206135396188|3|3338353030|60|0.6109748797816256|0|47|523|-80.562829|64|35.006282|FRESH POTATOES|0.0|4|RUSSET POTATO 8LB BAG|fc071cb340f590098059b243adcc4f3d508a1ea8|19.429895879212022|0.61242566243833529|00033383530307|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|1
35.006282|a9b035f0e6a034e9478caee894dd3f36108d27ba|6.68|2015-01-26 13:30:00|1.4091206135396188|3|7047043332|60|0.6109748797816256|0|47|685|-80.562829|61|35.006282|GREEK|1.6800000000000002|3|YOPLAIT GREEK 100 BLK CHERRY|fc071cb340f590098059b243adcc4f3d508a1ea8|19.429895879212022|0.61242566243833529|00070470435794|YOGURT|DAIRY|-80.562829|1.4060866207711706|60|5
35.006282|ba208af73d97f974e7f4caa857fc4fdbf7c683b4|1.24|2015-03-09 13:48:00|1.4091206135396188|3||60|0.6109748797816256|0|47|565|-80.562829|64|35.006282|REDUCED PRODUCE|0.0|4|PRODUCE REWRAP BY CT|fc071cb340f590098059b243adcc4f3d508a1ea8|19.429895879212022|0.61242566243833529|00204845000007|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|2
35.006282|319b731309dc2deab16994c8916ead554d03c5b7|1.98|2015-01-21 13:44:00|1.4091206135396188|3||60|0.6109748797816256|0|47|565|-80.562829|64|35.006282|REDUCED PRODUCE|0.0|4|PRODUCE REWRAP BY CT|fc071cb340f590098059b243adcc4f3d508a1ea8|19.429895879212022|0.61242566243833529|00204845000007|FRESH PRODUCE|PRODUCE|-80.562829|1.4060866207711706|60|2
35.006282|b3abfc88d9c055314d1c9419a65a68acd271a675|1.49|2015-02-09 13:30:00|1.4091206135396188|3|7203670302|60|0.6109748797816256|0|47|728|-80.562829|72|35.006282|NFS-PLASTIC FLATWARE|0.0|1|YH OCCASIONS FS FORKS|fc071cb340f590098059b243adcc4f3d508a1ea8|19.429895879212022|0.61242566243833529|00072036703019|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.562829|1.4060866207711706|60|1
35.006282|c64d3b1d1232defb4d7a45b298c466162e045e6a|8.370000000000001|2014-11-03 13:47:00|1.4091206135396188|3|7203670356|60|0.6109748797816256|0|47|442|-80.562829|76|35.006282|NFS-COOKING-STORAGE BAGS|5.37|1|YH FREEZER BAGS PINT 20CT|fc071cb340f590098059b243adcc4f3d508a1ea8|19.429895879212022|0.61242566243833529|00072036703569|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.562829|1.4060866207711706|60|3
35.006282|8c24216a18eb9ee39af3f9f6192b9e3da0bb1d39|3.89|2014-09-19 13:59:00|1.4091206135396188|3|4400003219|60|0.6109748797816256|0|47|1249|-80.562829|12|35.006282|CHOCOLATE CHIP COOKIES|1.94|1|CHIPS AHOY CHEWY|fc071cb340f590098059b243adcc4f3d508a1ea8|19.429895879212022|0.61242566243833529|00044000032234|COOKIES|G1 GROCERY|-80.562829|1.4060866207711706|60|1
35.006282|1482020a419462008888ad80a0f52a8b4ec937c8|179.89999999999998|2014-12-05 13:32:00|1.4091206135396188|3|7203678085|60|0.6109748797816256|0|47|665|-80.562829|145|35.006282|PACKAGED RAW|0.0|12|FISHERMANS SHRIMP 21/30 EZP WH|fc071cb340f590098059b243adcc4f3d508a1ea8|19.429895879212022|0.61242566243833529|00072036780850|SHRIMP|SEAFOOD|-80.562829|1.4060866207711706|60|5
35.006282|7e321c4bc18cfd152879879d82df011f21787eb5|4.19|2014-11-21 17:32:00|1.4091206135396188|3|2100000201|60|0.6109748797816256|0|47|317|-80.562829|52|35.006282|CHUNK AND BAR CHEESE|1.69|3|KRAFT SHARP CHEDDAR CHUNK|fc071cb340f590098059b243adcc4f3d508a1ea8|19.429895879212022|0.61242566243833529|00021000002016|CHEESE|DAIRY|-80.562829|1.4060866207711706|60|1
35.006282|0807aa0509ec3464b34da0760ab53735b8d93ec2|26.97|2014-12-16 17:40:00|1.4091206135396188|3|4900003165|60|0.6109748797816256|0|47|31|-80.562829|4|35.006282|NON CARBONATED WATER|4.5|1|DASANI .5 LITER 24 PK|fc071cb340f590098059b243adcc4f3d508a1ea8|19.429895879212022|0.61242566243833529|00049000031652|BOTTLED WATER|G1 GROCERY|-80.562829|1.4060866207711706|60|3
35.006282|79074166456a4585d70e6323eeea3289a3c05321|6.3|2015-02-25 13:55:00|1.4091206135396188|3|4060034500|60|0.6109748797816256|0|47|313|-80.562829|51|35.006282|MARGARINE|2.3|3|ICBINB SPREAD BOWL|fc071cb340f590098059b243adcc4f3d508a1ea8|19.429895879212022|0.61242566243833529|00040600345002|BUTTER & MARGARINE|DAIRY|-80.562829|1.4060866207711706|60|2
35.006282|02cd4239c39597c9fcdf74610c2265c48b413861|2.0|2014-12-08 13:53:00|1.4091206135396188|3|7203641150|60|0.6109748797816256|0|47|247|-80.562829|39|35.006282|VEGETABLES-FLANKER|0.0|1|HT SAUERKRAUT SHREDDED|fc071cb340f590098059b243adcc4f3d508a1ea8|19.429895879212022|0.61242566243833529|00072036411501|VEGETABLES-CAN/JAR|G1 GROCERY|-80.562829|1.4060866207711706|60|2
35.006282|709b047245863f94cbb1b529d92e9d5da2b93c39|4.38|2014-10-31 17:43:00|1.4091206135396188|3|4900005010|60|0.6109748797816256|0|47|55|-80.562829|8|35.006282|REGULAR|0.4|23|CLASSIC COKE 2 LT CONTOUR|fc071cb340f590098059b243adcc4f3d508a1ea8|19.429895879212022|0.61242566243833529|00049000050103|CARBONATED BEVERAGES|BEVERAGE|-80.562829|1.4060866207711706|60|2
35.006282|557a71275f861fd0cf6808a9ffde5e20620fba0e|6.78|2014-11-14 17:45:00|1.4091206135396188|3|20165700000|60|0.6109748797816256|0|47|297|-80.562829|49|35.006282|GROUND BEEF|1.51|2|HT GROUND BEEF CHUCK 80% LEAN|fc071cb340f590098059b243adcc4f3d508a1ea8|19.429895879212022|0.61242566243833529|00201657000003|BEEF|MEAT|-80.562829|1.4060866207711706|60|1
35.006282|b229cf6983831b4fa879b5ab89c5ab43b4f6aef8|40.89|2014-12-17 13:43:00|1.4091206135396188|3|20140400000|60|0.6109748797816256|0|47|296|-80.562829|49|35.006282|RANCHER BEEF|17.05|2|BEEF LOIN NY STRIP STEAK BNLS|fc071cb340f590098059b243adcc4f3d508a1ea8|19.429895879212022|0.61242566243833529|00201404000003|BEEF|MEAT|-80.562829|1.4060866207711706|60|3
35.006282|30b8d0dffe7a3c0a84a3592b675727a588ab6bd6|6.02|2015-03-06 17:22:00|1.4091206135396188|3|20165700000|60|0.6109748797816256|0|47|297|-80.562829|49|35.006282|GROUND BEEF|1.34|2|HT GROUND BEEF CHUCK 80% LEAN|fc071cb340f590098059b243adcc4f3d508a1ea8|19.429895879212022|0.61242566243833529|00201657000003|BEEF|MEAT|-80.562829|1.4060866207711706|60|1
35.006282|3d46f46374b9a66d0b798f467f5bc9f33ccb160e|2.59|2014-10-16 17:50:00|1.4091206135396188|3|5100017520|60|0.6109748797816256|0|47|1201|-80.562829|33|35.006282|RTS CANNED|1.09|1|CAM HOMESTYLE CHICKEN NOODLE|fc071cb340f590098059b243adcc4f3d508a1ea8|19.429895879212022|0.61242566243833529|00051000016591|SOUP|G1 GROCERY|-80.562829|1.4060866207711706|60|1
35.006282|1c0653088189e0c24cce0f56cbcc535d1840b8fd|6.25|2014-11-17 13:41:00|1.4091206135396188|3|2400016286|60|0.6109748797816256|0|47|245|-80.562829|39|35.006282|VEGETABLES-CORE|0.0|1|DEL MONTE GRN BEANS CUT|fc071cb340f590098059b243adcc4f3d508a1ea8|19.429895879212022|0.61242566243833529|00024000162865|VEGETABLES-CAN/JAR|G1 GROCERY|-80.562829|1.4060866207711706|60|5
35.006282|14db77c762b82a1be5814bcb637efb0f71970383|19.98|2015-02-13 13:52:00|1.4091206135396188|3|7203695262|60|0.6109748797816256|0|47|1671|-80.562829|383|35.006282|CHEESE CAKE|6.0|14|HAZELNUT CHEESECAKE|fc071cb340f590098059b243adcc4f3d508a1ea8|19.429895879212022|0.61242566243833529|00072036953285|PASTRY CASE|BAKERY|-80.562829|1.4060866207711706|60|2
35.006282|74c196debae868cbf97c1d4b7557d7d457665e51|4.69|2014-09-25 13:41:00|1.4091206135396188|3|4900002468|60|0.6109748797816256|0|47|55|-80.562829|8|35.006282|REGULAR|2.34|23|CLASSIC COKE .5 LITER/6 PK.|fc071cb340f590098059b243adcc4f3d508a1ea8|19.429895879212022|0.61242566243833529|00049000024685|CARBONATED BEVERAGES|BEVERAGE|-80.562829|1.4060866207711706|60|1
35.006282|82667d948d551d6db849db4e76221e7813ed55c0|7.36|2015-02-11 13:33:00|1.4091206135396188|3|20191100000|60|0.6109748797816256|0|47|299|-80.562829|49|35.006282|ANGUS BEEF|0.0|2|ANGUS BEEF BNLS CHUCKEYE STEAK|fc071cb340f590098059b243adcc4f3d508a1ea8|19.429895879212022|0.61242566243833529|00201911000008|BEEF|MEAT|-80.562829|1.4060866207711706|60|1
35.444064|e4c0f946739b20253def55b61a422d2daf19a5ad|1.26|2014-12-01 11:23:00|80.995508130988839|4||121|35.534326613896404|0|40|558|-80.895009|64|35.603432|SPECIALTY-VEGETABLES|0.0|4|COO GINGER ROOT, BULK|fcfb95bba64a3f99397eb8a57df3422c598930e4|6.236942512230774|35.466476270328783|00204612000001|FRESH PRODUCE|PRODUCE|-80.995484|80.995717779578086|274|1
35.444064|ea093c85b13986dd8de282a12f81bd858edcac9c|5.2|2015-01-13 11:46:00|1.4102725052409182|3||121|0.6186156170875914|0|1|500|-80.995484|64|35.444064|FRESH APPLES|0.0|4|HONEY CRISP APPLE|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00233283000003|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|293c92ce71ebf6ec46d90e553fcd82360cd62948|3.89|2015-01-20 17:40:00|1.4102725052409182|3|7247000222|121|0.6186156170875914|0|1|1641|-80.995484|377|35.444064|PACKAGED DONUTS|0.0|14|K K 6 ORIG GLAZED DONUT  PP|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00072470002228|DONUTS|BAKERY|-80.995484|1.413637875046387|121|1
35.444064|9ad6e39b53d2ff640d88542b2b9e3090efb2ff39|3.89|2014-09-27 20:26:00|1.4102725052409182|3|7247000222|121|0.6186156170875914|0|1|1641|-80.995484|377|35.444064|PACKAGED DONUTS|0.0|14|K K 6 ORIG GLAZED DONUT  PP|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00072470002228|DONUTS|BAKERY|-80.995484|1.413637875046387|121|1
35.444064|1558ee043aaa3106fa7c91dc9afb12b4980cf4d5|3.89|2015-01-29 11:41:00|1.4102725052409182|3|7247000222|121|0.6186156170875914|0|1|1641|-80.995484|377|35.444064|PACKAGED DONUTS|0.0|14|K K 6 ORIG GLAZED DONUT  PP|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00072470002228|DONUTS|BAKERY|-80.995484|1.413637875046387|121|1
35.444064|0d73870420486ab6a5479528e66e52146cf6ad6e|2.69|2014-12-14 20:26:00|80.995508130988839|3|7940073830|121|35.516991377409113|0|40|3545|-80.945176|1045|35.323246|SHAMPOO-VALUE|0.0|17|SUAVE MEN DAILY CLN OCEAN SHAM|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|35.466476270328783|00079400128041|HAIR & SCALP CARE|HBC|-80.995484|80.995575828289404|166|1
35.444064|c95080c3f57ae8cf6ded127d7878813a0d692860|11.1|2014-12-08 18:30:00|1.4102725052409182|3|20895700000|121|0.6186156170875914|0|1|977|-80.995484|201|35.444064|FRESH HT CHICKEN|3.87|2|HT VALUE PK CHCKN LEG QUARTERS|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00208957000009|POULTRY|MEAT|-80.995484|1.413637875046387|121|1
35.444064|7199fdb3b874ad3ce476f2feef48b31b9d4da0e2|6.25|2014-11-28 12:03:00|1.4102725052409182|3|2400016286|121|0.6186156170875914|0|1|245|-80.995484|39|35.444064|VEGETABLES-CORE|0.0|1|DEL MONTE GRN BEANS LS|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00024000566670|VEGETABLES-CAN/JAR|G1 GROCERY|-80.995484|1.413637875046387|121|5
35.444064|3a8442509fa1ae74c239ec9bc3518c677ff62be1|4.29|2014-10-24 12:02:00|1.4102725052409182|3|2840016014|121|0.6186156170875914|0|1|201|-80.995484|31|35.444064|POTATO CHIPS|2.15|1|LAYS CLASSIC|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00028400160148|SNACKS|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|3d101fd0b386e78a0724decbb41a13ad68270ca0|3.25|2014-11-16 19:47:00|1.4102725052409182|3|3120020007|121|0.6186156170875914|0|1|130|-80.995484|20|35.444064|CRANBERRY JUICE/DRINKS-SHELF|1.63|1|OSPRAY CRANBERRY JUICE|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00031200200075|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|1f897a1274d88ba3c734ddedeac1887df45c3488|4.49|2015-02-19 16:29:00|80.995508130988839|3|70897191777|121|35.516991377409113|0|40|1703|-80.945176|387|35.323246|SEASONAL COOKIES|0.0|14|VALENTINE PINK FRSTD CHOC COOK|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|35.466476270328783|00708971917777|COOKIES|BAKERY|-80.995484|80.995575828289404|166|1
35.444064|39212430d9b581757acffdead459b14b16d569b9|3.98|2015-02-21 19:23:00|1.4102725052409182|3|88439506246|121|0.6186156170875914|0|1|115|-80.995484|16|35.444064|REMAINING FRUIT|0.0|1|LUCKS FRIED APPLES|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00884395062467|FRUIT-CAN/JAR|G1 GROCERY|-80.995484|1.413637875046387|121|2
35.444064|ed14fc799865e698c7e7a4b5523712ee87c8da23|3.98|2014-09-20 17:39:00|1.4102725052409182|3|88439506246|121|0.6186156170875914|0|1|115|-80.995484|16|35.444064|REMAINING FRUIT|0.98|1|LUCKS FRIED APPLES|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00884395062467|FRUIT-CAN/JAR|G1 GROCERY|-80.995484|1.413637875046387|121|2
35.444064|bdcedae4988be7c8959a9ca5bef677cc6eadc6da|3.25|2014-12-16 16:06:00|1.4102725052409182|3|7203656080|121|0.6186156170875914|0|1|318|-80.995484|52|35.444064|SHREDDED/GRATED CHEESE|3.25|3|HT NACHO TACO MEXICAN BLEND|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00072036560834|CHEESE|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|4bd3ab237d7a05db450d1095015faacf34f651e0|2.89|2014-11-14 16:53:00|1.4102725052409182|3|7203663102|121|0.6186156170875914|0|1|339|-80.995484|57|35.444064|EGGNOGS/DRINKS|0.39|3|I/O HARRIS TEETER EGG NOG|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00072036631022|MILK|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|188d89211b2019221a29053ed1617bc2f15163fa|5.78|2014-12-27 13:47:00|1.4102725052409182|3|7203663102|121|0.6186156170875914|0|1|339|-80.995484|57|35.444064|EGGNOGS/DRINKS|0.78|3|I/O HARRIS TEETER EGG NOG|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00072036631022|MILK|DAIRY|-80.995484|1.413637875046387|121|2
35.444064|04ee770ac100fa6fd3521998d5189d42a6850ca0|2.89|2014-11-22 19:32:00|80.995508130988839|3|7203663102|121|35.516991377409113|0|40|339|-80.945176|57|35.323246|EGGNOGS/DRINKS|0.39|3|I/O HARRIS TEETER EGG NOG|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|35.466476270328783|00072036631022|MILK|DAIRY|-80.995484|80.995575828289404|166|1
35.444064|1027a16f20c362249c132176ce686bbfefae9ac6|5.78|2014-12-06 12:10:00|1.4102725052409182|3|7203663102|121|0.6186156170875914|0|1|339|-80.995484|57|35.444064|EGGNOGS/DRINKS|1.78|3|I/O HARRIS TEETER EGG NOG|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00072036631022|MILK|DAIRY|-80.995484|1.413637875046387|121|2
35.444064|bee9196bc52a6bbda5891835c897d8bc7692c232|2.29|2015-02-01 20:58:00|1.4102725052409182|3|7203663996|121|0.6186156170875914|0|1|342|-80.995484|57|35.444064|FRESH MILK|0.82|3|HARRIS TEETER WHOLE MILK|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00072036639967|MILK|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|6216a6303ddced9c075ab63b872fda2c7384a55c|2.29|2015-01-09 18:46:00|1.4102725052409182|3|7203663996|121|0.6186156170875914|0|1|342|-80.995484|57|35.444064|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00072036631299|MILK|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|c585e155b114605fbdb355dcda2a55c2bb52fc4f|2.19|2014-09-13 18:22:00|1.4102725052409182|3|7203670343|121|0.6186156170875914|0|1|443|-80.995484|76|35.444064|NFS-GARBAGE BAGS|0.41|1|YH SMALL GARBAGE TWST TIE 4 GL|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00072036704955|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|aa9ba0c52bbff58f226c8a8ec5c6ff7a8ec2b229|3.69|2014-09-24 20:41:00|1.4102725052409182|3|7127925101|121|0.6186156170875914|0|1|555|-80.995484|64|35.444064|PACKAGED SALADS|0.0|4|F.E. AMERICAN SALAD|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00071279241005|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|6184f205b4f65c89fdeb239368aaf0a99d53c99d|3.58|2014-11-04 20:19:00|1.4102725052409182|3|5100001047|121|0.6186156170875914|0|1|212|-80.995484|33|35.444064|CONDENSED SOUP|1.58|1|CAMP COND CREAM OF ONION|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00051000016171|SOUP|G1 GROCERY|-80.995484|1.413637875046387|121|2
35.444064|daaca57f9080b5b928756e53735ac618c6b3e730|1.94|2014-11-18 19:06:00|1.4102725052409182|3|5210007086|121|0.6186156170875914|0|1|217|-80.995484|34|35.444064|EXTRACTS FOOD COLORING|0.58|1|E  MCCORMICK VANILLA EXTRACT|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00052100070865|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.995484|1.413637875046387|121|2
35.444064|dece9c136c0d8cbae14d01539bc06b07481294f4|1.27|2014-09-16 16:39:00|80.995508130988839|3|5963500189|121|35.516991377409113|0|40|1461|-80.945176|40|35.323246|FROZEN GARLIC TOAST AND BRD|0.0|5|FURLANI TEXAS TOAST|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|35.466476270328783|00059635001890|FROZEN DOUGH|FROZEN|-80.995484|80.995575828289404|166|1
35.444064|f3faa097e10d632e9af159f107e9e6b61029b304|1.27|2014-10-08 20:56:00|1.4102725052409182|3|5963500189|121|0.6186156170875914|0|1|1461|-80.995484|40|35.444064|FROZEN GARLIC TOAST AND BRD|0.0|5|FURLANI TEXAS TOAST|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00059635001890|FROZEN DOUGH|FROZEN|-80.995484|1.413637875046387|121|1
35.444064|815124ec54a12e1029beb1ae7b8c36cceecd15c3|3.99|2014-11-11 14:19:00|1.4102725052409182|3|7127930108|121|0.6186156170875914|0|1|555|-80.995484|64|35.444064|PACKAGED SALADS|0.0|4|F.E. BACON CAESAR KIT|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00071279301082|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|efa2b56269d96064f3319312048f696ddff720e4|1.69|2015-01-06 18:05:00|80.995508130988839|3|7203688003|121|35.516991377409113|0|40|527|-80.945176|64|35.323246|FRESH CARROTS|0.0|4|HT BABY CARROTS 1LB BAG|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|35.466476270328783|00072036880031|FRESH PRODUCE|PRODUCE|-80.995484|80.995575828289404|166|1
35.444064|978835bc56af3589e29ccaa3a2f891cbbef91526|7.69|2015-03-03 09:50:00|1.4102725052409182|3|1380010334|121|0.6186156170875914|0|1|1280|-80.995484|48|35.444064|MULTI SERVE MEALS|0.0|5|STOUFFER FM/STYLE MAC/CHEESE|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00013800103345|FROZEN MEALS|FROZEN|-80.995484|1.413637875046387|121|1
35.444064|9aca3cecf14de105885955fc62c9670799e648e0|2.99|2015-02-08 14:29:00|80.995508130988839|3|7433610102|121|35.516991377409113|0|40|342|-80.945176|57|35.323246|FRESH MILK|0.0|3|HIGHLAND CREST WHOLE MILK|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|35.466476270328783|00074336879203|MILK|DAIRY|-80.995484|80.995575828289404|166|1
35.444064|b449d90cd0df3c4f17d7febc45fbb49eb0a041c8|2.99|2015-03-08 19:49:00|1.4102725052409182|3|7433610102|121|0.6186156170875914|0|1|342|-80.995484|57|35.444064|FRESH MILK|0.0|3|HIGHLAND CREST WHOLE MILK|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00074336879203|MILK|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|45bf0342b0d5f7b99389507fe121b869ece85306|7.47|2015-01-11 19:16:00|1.4102725052409182|3|20140400000|121|0.6186156170875914|0|1|296|-80.995484|49|35.444064|RANCHER BEEF|0.0|2|BEEF LOIN NY STRIP STEAK BNLS|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00201404000003|BEEF|MEAT|-80.995484|1.413637875046387|121|1
35.444064|0b8c96b3114c752a1a7d157c8f22535bb9f7b781|3.34|2015-02-28 14:07:00|1.4102725052409182|3|7203643010|121|0.6186156170875914|0|1|252|-80.995484|45|35.444064|PREMIUM ICE CREAM|1.37|5|HT PREM BANANA PUDDING IC|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00072036430311|ICE CREAM|FROZEN|-80.995484|1.413637875046387|121|1
35.444064|5c10358dc73b75b170ef465298d3b3cbd3e6bc22|3.34|2014-10-06 19:48:00|1.4102725052409182|3|7203643010|121|0.6186156170875914|0|1|252|-80.995484|45|35.444064|PREMIUM ICE CREAM|0.84|5|HT PREM BANANA PUDDING IC|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00072036430311|ICE CREAM|FROZEN|-80.995484|1.413637875046387|121|1
35.444064|83c406c3b8dba83b1054ff03fd11254f782126bc|7.89|2015-02-03 19:43:00|1.4102725052409182|3|1380014333|121|0.6186156170875914|0|1|1280|-80.995484|48|35.444064|MULTI SERVE MEALS|0.9|5|STOUF LIMITED ED MAC N CHS|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00013800713049|FROZEN MEALS|FROZEN|-80.995484|1.413637875046387|121|1
35.444064|699024adc3b4abbed6d0345055fa64a72f0c5532|2.77|2014-10-14 21:15:00|1.4102725052409182|3|3338353030|121|0.6186156170875914|0|1|523|-80.995484|64|35.444064|FRESH POTATOES|0.0|4|RUSSET POTATO 8LB BAG|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00033383530307|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|074e245b181d0aae949e07740f716cc70d1ca723|2.77|2015-01-04 19:36:00|1.4102725052409182|3|3338353030|121|0.6186156170875914|0|1|523|-80.995484|64|35.444064|FRESH POTATOES|0.0|4|RUSSET POTATO 8LB BAG|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00033383530307|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|7fcc43a811394a039282d0b1caf5f96b89054f55|3.99|2014-10-18 17:41:00|1.4102725052409182|3|4000015140|121|0.6186156170875914|0|1|46|-80.995484|7|35.444064|PKG CHOC|0.49|1|3 MUSKETEER FUN SIZE|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00040000151227|CANDY|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|757ea8cd5079db76ce389f68dd455a5f2f63d13b|21.98|2014-10-26 20:01:00|1.4102725052409182|3|3040077569|121|0.6186156170875914|0|1|427|-80.995484|72|35.444064|NFS-TOILET TISSUE|6.0|1|ANGEL SOFT SOFT/STRONG 16R|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00030400775697|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.995484|1.413637875046387|121|2
35.444064|cd6da362b3a6fe15b1cfeb0fa63233116e73caf3|3.49|2015-01-18 19:40:00|1.4102725052409182|3|7203663995|121|0.6186156170875914|0|1|342|-80.995484|57|35.444064|FRESH MILK|0.92|3|HARRIS TEETER WHOLE MILK|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00072036639950|MILK|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|1ca3913b1c65e77ba0e6d6bb796d00226e83a866|3.99|2014-10-12 19:48:00|1.4102725052409182|3|7203663995|121|0.6186156170875914|0|1|342|-80.995484|57|35.444064|FRESH MILK|1.02|3|HARRIS TEETER WHOLE MILK|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00072036639950|MILK|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|993c6c26bae5b31b6921dfe6668a06ec3b3bd76d|1.19|2014-11-13 14:57:00|1.4102725052409182|3|4144310211|121|0.6186156170875914|0|1|247|-80.995484|39|35.444064|VEGETABLES-FLANKER|0.0|1|M HOLMES COLLARD GREENS|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00041443102111|VEGETABLES-CAN/JAR|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|bb13e71ebfb33b21536cca957ffbd6021a88b4c3|4.69|2014-11-24 19:51:00|1.4102725052409182|3|4900002468|121|0.6186156170875914|0|1|55|-80.995484|8|35.444064|REGULAR|4.69|23|M MAID LIGHT LEMONADE 6PK .5L|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00025000058738|CARBONATED BEVERAGES|BEVERAGE|-80.995484|1.413637875046387|121|1
35.444064|445b9c57eb6ae525e8076189d893a0bb4c0e60ad|6.99|2015-01-24 18:35:00|1.4102725052409182|3|30031873512|121|0.6186156170875914|0|1|4236|-80.995484|1200|35.444064|DEX ADULT/CHILDREN|0.0|17|ROBITUSSIN PK M-SYM COLD NT LQ|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00300318735121|COUGH/COLD/SINUS|HBC|-80.995484|1.413637875046387|121|1
35.444064|bce994c1a34d5d35b09629e823e54812f4c77cd6|0.5|2014-12-30 13:24:00|1.4102725052409182|3||121|0.6186156170875914|0|1|543|-80.995484|64|35.444064|FRESH GARLIC|0.0|4|COO GARLIC, WHITE, BULK|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00204608000008|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|66859f68c317c3e0794eb835449a3530ff6ae854|6.99|2014-10-28 19:30:00|80.995508130988839|3|2370001450|121|35.516991377409113|0|40|291|-80.945176|48|35.323246|FROZEN POUTLRY|0.0|5|TYSON CHICKEN NUGGETS 32OZ|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|35.466476270328783|00023700028471|FROZEN MEALS|FROZEN|-80.995484|80.995575828289404|166|1
35.444064|2e9e5f48767572576189d7d2f9f7bb79b3570231|0.97|2015-01-22 16:04:00|80.995508130988839|3|7203604053|121|35.516991377409113|0|40|51|-80.945176|7|35.323246|MARSHMALLOWS|0.0|1|HT MINI MARSHMALLOW|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|35.466476270328783|00072036040534|CANDY|G1 GROCERY|-80.995484|80.995575828289404|166|1
35.444064|0cff10fc8b8bf7840190ac24b7609d912e8e267d|1.49|2014-11-17 16:55:00|80.995508130988839|3|7203653022|121|35.516991377409113|0|40|1273|-80.945176|50|35.323246|BAG VEG NON STEAM|0.0|5|HT CHOPPED BROCCOLI|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|35.466476270328783|00072036530783|VEGETABLES-FROZEN|FROZEN|-80.995484|80.995575828289404|166|1
35.444064|a141f64407ef41f4e73e4f88a3393b968b1a40f3|12.19|2014-09-20 17:48:00|1.4102725052409182|3|1380023260|121|0.6186156170875914|0|1|1280|-80.995484|48|35.444064|MULTI SERVE MEALS|3.22|5|STOUFFER LASAGNA|fd858fd3e8fcc494574aab53184261e7e66e3d41|5.039108314631327|0.61833652052202714|00013800232601|FROZEN MEALS|FROZEN|-80.995484|1.413637875046387|121|1
35.17739|e2eda0c09c33c2eb1403ce1b86131804ad9ec187|0.79|2015-02-23 16:10:00|1.4094857484078087|4||208|0.613961277758128|0|26|532|-80.80146|64|35.17739|FRESH CUCUMBERS|0.0|4|COO CUCUMBERS S/S|0c1614152cefab11d7f01e51c313347a9ea2af16|1.379660302971585|0.61471665291522548|00204062000002|FRESH PRODUCE|PRODUCE|-80.80146|1.4102515174184975|208|1
35.17739|6d0bb512e462417821d5b5395db0c76137e7eca2|1.39|2014-11-30 14:55:00|1.4094857484078087|4|2200000488|208|0.613961277758128|0|26|48|-80.80146|7|35.17739|REGISTER GUM|0.0|1|(FE)ORBIT MINT GUM 14PC|0c1614152cefab11d7f01e51c313347a9ea2af16|1.379660302971585|0.61471665291522548|00022000004833|CANDY|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|e4a9bbad693718b672bc0b45b456385ef4c97fcf|1.49|2015-01-03 15:20:00|1.4094857484078087|4||208|0.613961277758128|0|26|525|-80.80146|64|35.17739|FRESH LETTUCE|0.0|4|ICEBERG LETTUCE|0c1614152cefab11d7f01e51c313347a9ea2af16|1.379660302971585|0.61471665291522548|00204061000003|FRESH PRODUCE|PRODUCE|-80.80146|1.4102515174184975|208|1
35.17739|73722887bffedacc9d57a4ef6148b52c52665493|1.89|2015-03-09 13:48:00|1.4094857484078087|4|2700038249|208|0.613961277758128|0|26|70|-80.80146|11|35.17739|KETCHUP|0.89|1|HUNTS KETCHUP 24|0c1614152cefab11d7f01e51c313347a9ea2af16|1.379660302971585|0.61471665291522548|00027000382493|CONDIMENTS|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|609fae523fbe4ad4cd931c77b72922cd6251ec7d|3.08|2014-12-13 17:04:00|1.4094857484078087|4|7203636010|208|0.613961277758128|0|26|30|-80.80146|4|35.17739|CARBONATED WATER|0.68|1|HT SIMPLY CLR + B VIT KEY LIME|0c1614152cefab11d7f01e51c313347a9ea2af16|1.379660302971585|0.61471665291522548|00072036983671|BOTTLED WATER|G1 GROCERY|-80.80146|1.4102515174184975|208|4
35.17739|025cc2de0d3634cd082f85844c68e9c5220ec7bc|7.99|2014-11-25 13:11:00|1.4094857484078087|4|5200020805|208|0.613961277758128|0|26|171|-80.80146|20|35.17739|ISOTONIC DRINKS|2.99|1|GATORADE COOL BLUE 8PK|0c1614152cefab11d7f01e51c313347a9ea2af16|1.379660302971585|0.61471665291522548|00052000208443|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|dc95311a529539804064664b3bd647d4fd5bcebb|3.98|2014-10-17 13:53:00|80.801203185414451|4|4900004574|208|35.197356838147783|0|24|171|-80.844274|20|35.204336|ISOTONIC DRINKS|2.4|1|POWERADE LEMON LIME|0c1614152cefab11d7f01e51c313347a9ea2af16|1.379660302971585|35.194272495053255|00049000045734|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.80146|80.801462110476464|61|2
35.17739|cd96b2e3eab30339f47ec465d17ccdf4dd3693ab|3.98|2015-02-11 19:46:00|80.801203185414451|4|4900004574|208|35.197356832805845|0|24|171|-80.824767|20|35.116751|ISOTONIC DRINKS|2.4|1|POWERADE GRAPE|0c1614152cefab11d7f01e51c313347a9ea2af16|1.379660302971585|35.194272495053255|00049000045239|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.80146|80.801477995337251|294|2
35.17739|334682fe2d872d388542d2c0d8d8b5fa8cf548ee|9.99|2014-11-19 17:22:00|80.801203185414451|4|1820011047|208|35.197356837664685|0|24|455|-80.85013|82|35.175855|DOMESTIC PREMIUM 12PK&>|0.0|16|BUD 12PK 12OZ CAN|0c1614152cefab11d7f01e51c313347a9ea2af16|1.379660302971585|35.194272495053255|00018200110474|DOMESTIC BEER|BEER|-80.80146|80.801465773820624|218|1
35.17739|1985383f3b7f53b93a9ffe5fb2e7d723dec18acf|7.99|2014-10-06 19:10:00|1.4094857484078087|4|5200020805|208|0.613961277758128|0|26|171|-80.80146|20|35.17739|ISOTONIC DRINKS|3.99|1|GATORADE GLACIER CHERRY 8PK|0c1614152cefab11d7f01e51c313347a9ea2af16|1.379660302971585|0.61471665291522548|00052000102451|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|136936bc25b7608aaf351cb4f19c3a139addfc66|2.31|2014-11-08 18:30:00|1.4094857484078087|4|7203636010|208|0.613961277758128|0|26|30|-80.80146|4|35.17739|CARBONATED WATER|0.0|1|HT SIMPLY CLEAR KEY LIME|0c1614152cefab11d7f01e51c313347a9ea2af16|1.379660302971585|0.61471665291522548|00072036360250|BOTTLED WATER|G1 GROCERY|-80.80146|1.4102515174184975|208|3
35.17739|2cef5b243882828ca8964c08004bbca81a61148a|1.54|2014-11-17 17:30:00|1.4094857484078087|4|7203636010|208|0.613961277758128|0|26|30|-80.80146|4|35.17739|CARBONATED WATER|0.34|1|HT SIMPLY CLEAR KEY LIME|0c1614152cefab11d7f01e51c313347a9ea2af16|1.379660302971585|0.61471665291522548|00072036360250|BOTTLED WATER|G1 GROCERY|-80.80146|1.4102515174184975|208|2
35.17739|bf98addc8a5277472da4c7f92979fed208a9f37d|6.57|2014-10-19 11:07:00|1.4094857484078087|4|5100013458|208|0.613961277758128|0|26|1499|-80.80146|33|35.17739|RTS MICROWAVE|1.57|1|CAMP MW BOWLS HR CHICKEN NOODL|0c1614152cefab11d7f01e51c313347a9ea2af16|1.379660302971585|0.61471665291522548|00051000195784|SOUP|G1 GROCERY|-80.80146|1.4102515174184975|208|3
34.977331|247ad00fe2cdddff2728834f006ad57366ccdeee|7.98|2015-02-06 18:59:00|81.02739863253349|3|85591900302|149|35.014573965463335|0|14|41|-80.847383|6|35.024464|BREAKFAST BARS|2.0|1|S BCH CEREAL BAR FIBER DK CHOC|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00855919003051|BREAKFAST FOODS|G1 GROCERY|-81.027334|81.027393142178198|317|2
34.977331|bae383edbf4ba1e13889c90687cfea4581ad74bd|3.99|2015-01-27 16:22:00|81.02739863253349|3|85420800508|149|35.014573965463335|0|14|577|-80.847383|136|35.024464|OTHER MERCH FR MSC JUICE|0.0|4|ORG. SUJA BERRY GOODNESS|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00854208005103|OTHER MERCHANDISE|PRODUCE|-81.027334|81.027393142178198|317|1
34.977331|064c6249d9657fe159438b759f1f88fa53d8b3c0|2.39|2014-11-25 06:10:00|81.02739863253349|3|78616250700|149|35.014573965463335|0|14|31|-80.847383|4|35.024464|NON CARBONATED WATER|0.4|1|CB GLACEAU SMART WATER|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00786162507006|BOTTLED WATER|G1 GROCERY|-81.027334|81.027393142178198|317|1
34.977331|45fe1712a4dc20c968829954dc1aff7e13b9f3ea|6.99|2014-10-18 07:27:00|81.02739863253349|3|1820005989|149|35.014573965463335|0|14|455|-80.847383|82|35.024464|DOMESTIC PREMIUM 12PK&>|0.0|16|MICHELOB ULTRA 6PK 12OZ  BTL|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00018200059896|DOMESTIC BEER|BEER|-81.027334|81.027393142178198|317|1
34.977331|bd73f7aafc5466d1a937cc7aa677edbebf71a661|2.99|2014-09-28 17:22:00|81.02739863253349|3|1380004717|149|35.014573965463335|0|14|1278|-80.847383|48|35.024464|SINGLE SERVE NUTRITIONAL|0.0|5|LC CAFE CLSSC 4 CHEESE PIZZA|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00013800047199|FROZEN MEALS|FROZEN|-81.027334|81.027393142178198|317|1
34.977331|b5eb2a62552ddfc1c0b97802b58446d1db2ee1f6|2.99|2014-10-13 15:43:00|81.02739863253349|3|1380004717|149|35.014573965463335|0|14|1278|-80.847383|48|35.024464|SINGLE SERVE NUTRITIONAL|0.0|5|LC CAFE CLSSC 4 CHEESE PIZZA|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00013800047199|FROZEN MEALS|FROZEN|-81.027334|81.027393142178198|317|1
34.977331|862615b5e291a4ee9b18e0c82915cf9fde993fdf|6.58|2014-12-13 09:56:00|81.02739863253349|3|79285014099|149|35.014573965463335|0|14|3272|-80.847383|1023|35.024464|NATURAL/ORGANIC PRODUCT|0.0|17|BURT B HONEY LIP BALM TUBE|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00792850136991|NATURAL PERSONAL CARE|HBC|-81.027334|81.027393142178198|317|2
34.977331|673660084168d78c94e29ef9933dd835cccc3e43|4.49|2014-12-06 12:20:00|81.02739863253349|3|85968600400|149|35.014573965463335|0|14|46|-80.847383|7|35.024464|PKG CHOC|0.0|1|BARKTHINS DRK CHOCOLATE MINT|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00859686004037|CANDY|G1 GROCERY|-81.027334|81.027393142178198|317|1
34.977331|f5ae6b13a8838f03aac73b9b01e8b5d16245455e|6.99|2014-12-23 16:07:00|81.02739863253349|3|3680009234|149|35.014573965463335|0|14|4353|-80.847383|1205|35.024464|SLEEPING AID|0.0|17|TC NIGHTTIME SLEEP AID CAPS|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00036800092341|PAIN RELIEF|HBC|-81.027334|81.027393142178198|317|1
34.977331|db8735f42fe6415843f4620085ce4b132aadc733|8.99|2014-12-21 16:07:00|81.02739863253349|3|76604700434|149|35.014573965463335|0|14|37|-80.847383|10|35.024464|PODS/CUPS/SINGLES|1.6|1|PANERA CUPS HAZELNUT 12CT|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00766047004363|COFFEE|G1 GROCERY|-81.027334|81.027393142178198|317|1
34.977331|608051d257bd4e93d5a36a46e28802f5f7cf1071|1.88|2014-10-05 18:58:00|81.02739863253349|3||149|35.014573965463335|0|14|502|-80.847383|64|35.024464|FRESH BANANAS|0.0|4|BANANAS, YELLOW|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00204011000008|FRESH PRODUCE|PRODUCE|-81.027334|81.027393142178198|317|1
34.977331|7c53c2d5926956ab44c46a136378e2bd3a21ce91|1.89|2015-02-18 20:12:00|81.02739863253349|3||149|35.014573965463335|0|14|502|-80.847383|64|35.024464|FRESH BANANAS|0.0|4|BANANAS, YELLOW|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00204011000008|FRESH PRODUCE|PRODUCE|-81.027334|81.027393142178198|317|1
34.977331|5bbeaff2b6c663e7e5909e6e5984ee964bb73640|2.22|2014-11-02 11:43:00|81.02739863253349|3||149|35.014573965463335|0|14|502|-80.847383|64|35.024464|FRESH BANANAS|0.0|4|BANANAS, YELLOW|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00204011000008|FRESH PRODUCE|PRODUCE|-81.027334|81.027393142178198|317|1
34.977331|b7ae85572105fe3b3674845563c86680da8a29e6|1.95|2014-09-24 19:15:00|81.02739863253349|3||149|35.014573948188662|0|14|502|-80.8062|64|35.037115|FRESH BANANAS|0.0|4|BANANAS, YELLOW|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00204011000008|FRESH PRODUCE|PRODUCE|-81.027334|81.027407588011428|27|1
34.977331|1fbcf9ca027bfffe39e12cb23f7c19647f42c342|3.99|2014-11-25 17:04:00|81.02739863253349|3|4667716926|149|35.014573965463335|0|14|6137|-80.847383|1546|35.024464|BULB-CARD FAN LIGHT|0.0|18|PHILIP 40 W DURAMAX LLBC FAN W|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00046677169268|LIGHT BULBS/ELECTRICAL|GM|-81.027334|81.027393142178198|317|1
34.977331|952d16a6af8a52b9ed7089b780a51a213cd2fc19|2.99|2014-10-23 19:07:00|81.02739863253349|3|3800035900|149|35.014573948188662|0|14|42|-80.8062|6|35.037115|GRANOLA/YOGURT BARS|0.0|1|KLG NUTRI GRN BAR FC APPLE COB|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00038000724145|BREAKFAST FOODS|G1 GROCERY|-81.027334|81.027407588011428|27|1
34.977331|ca53a2ba97ebf590485a8cdcb258a8e4c9cd4a32|2.52|2014-10-25 14:08:00|81.02739863253349|3||149|35.014573965463335|0|14|502|-80.847383|64|35.024464|FRESH BANANAS|0.0|4|BANANAS, YELLOW|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00204011000008|FRESH PRODUCE|PRODUCE|-81.027334|81.027393142178198|317|1
34.977331|73cdf9f198548f98d2246a23a30be5537c8e25e7|2.48|2015-03-03 16:06:00|81.02739863253349|3||149|35.014573965463335|0|14|502|-80.847383|64|35.024464|FRESH BANANAS|0.0|4|BANANAS, YELLOW|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00204011000008|FRESH PRODUCE|PRODUCE|-81.027334|81.027393142178198|317|1
34.977331|2b0a089f0fd0384a5eba72f26d4f088f58c0f264|2.29|2014-10-20 19:07:00|81.02739863253349|3||149|35.014573948188662|0|14|502|-80.8062|64|35.037115|FRESH BANANAS|0.0|4|BANANAS, YELLOW|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00204011000008|FRESH PRODUCE|PRODUCE|-81.027334|81.027407588011428|27|1
34.977331|ab30ff02adf32c458ace9e4bce642609470e3c41|1.94|2014-11-25 16:12:00|81.02739863253349|3||149|35.014573965463335|0|14|502|-80.847383|64|35.024464|FRESH BANANAS|0.0|4|BANANAS, YELLOW|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00204011000008|FRESH PRODUCE|PRODUCE|-81.027334|81.027393142178198|317|1
34.977331|d4e46dd24c0e41f50a56f7ce37670a9da5468ac2|1.66|2014-09-11 17:10:00|81.02739863253349|3||149|35.014573965463335|0|14|502|-80.847383|64|35.024464|FRESH BANANAS|0.0|4|BANANAS, YELLOW|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00204011000008|FRESH PRODUCE|PRODUCE|-81.027334|81.027393142178198|317|1
34.977331|a09bebcef30525120ebc92e4cb67a32e90cca7ba|1.81|2014-12-07 17:38:00|81.02739863253349|3||149|35.014573965463335|0|14|502|-80.847383|64|35.024464|FRESH BANANAS|0.0|4|BANANAS, YELLOW|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00204011000008|FRESH PRODUCE|PRODUCE|-81.027334|81.027393142178198|317|1
34.977331|454fccb33b7c17ddf3ca5577eaf9ecedeea6c6dd|1.77|2014-10-11 09:19:00|81.02739863253349|3||149|35.014573965463335|0|14|502|-80.847383|64|35.024464|FRESH BANANAS|0.0|4|BANANAS, YELLOW|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00204011000008|FRESH PRODUCE|PRODUCE|-81.027334|81.027393142178198|317|1
34.977331|d71651d8cb46691fc9224d3e35dca3b5b905c231|1.85|2014-11-19 18:50:00|81.02739863253349|3||149|35.014573965463335|0|14|502|-80.847383|64|35.024464|FRESH BANANAS|0.0|4|BANANAS, YELLOW|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00204011000008|FRESH PRODUCE|PRODUCE|-81.027334|81.027393142178198|317|1
34.977331|52e7f26c82cd15de1688d3ae2840c05322781256|8.99|2015-03-07 17:26:00|81.02739863253349|3|76604700405|149|35.014573965463335|0|14|36|-80.847383|10|35.024464|PREMIUM GROUND|2.0|1|PANERA HAZELNUT CREME COFFEE|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00766047004097|COFFEE|G1 GROCERY|-81.027334|81.027393142178198|317|1
34.977331|e190189d709772be99bfb2265005161e9b8ed724|3.99|2014-11-26 20:51:00|81.02739863253349|3|7203698715|149|35.014573965463335|0|14|4353|-80.847383|1205|35.024464|SLEEPING AID|0.0|17|HT REST SIMPLY CAPS|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00072036987150|PAIN RELIEF|HBC|-81.027334|81.027393142178198|317|1
34.977331|5acb3ba0da2312eb2be6acc067782ea88d943a44|5.99|2014-10-08 16:25:00|81.02739863253349|3|8500001752|149|35.014573965463335|0|14|9938|-80.847383|885|35.024464|NFS POP PINOT GRS/GRIGIO|0.0|13|THE NAKED GRAPE PINOT GRIGIO|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00085000017524|POPULAR (4-$7.99)|WINE|-81.027334|81.027393142178198|317|1
34.977331|748212ac8e0ed5a911b91141526daf520bfa4d68|2.78|2014-12-10 18:56:00|81.02739863253349|3|7203676368|149|35.014573948188662|0|14|1212|-80.8062|272|35.037115|HISP BEANS/PEPPERS|0.0|1|HTO REFRIED BLACK BEANS|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00072036976710|HISPANIC PREP. FOODS|G1 GROCERY|-81.027334|81.027407588011428|27|2
34.977331|1953fb39de6c1b408cbfb5bf75cd809a13a22730|0.97|2014-11-26 18:51:00|81.02739863253349|3|4300020431|149|35.014573965463335|0|14|94|-80.847383|14|35.024464|PUDDING MIXES|0.22|1|JELL-O BUTTERSCOTCH PUDDING|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00043000206539|DESSERTS/GELS/SYRUPS|G1 GROCERY|-81.027334|81.027393142178198|317|1
34.977331|59d55d86915ed61dc70bb583347b138fac3a4ac6|3.39|2015-01-28 06:36:00|81.02739863253349|3|4000042065|149|35.014573965463335|0|14|46|-80.847383|7|35.024464|PKG CHOC|0.0|1|I/O MM MILK CHOCOLATE BONUS|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00040000420651|CANDY|G1 GROCERY|-81.027334|81.027393142178198|317|1
34.977331|df17f71b9bb34b1a5304761913d39c9c7d55af5e|7.99|2014-10-30 16:01:00|81.02739863253349|3|1820013986|149|35.014573965463335|0|14|458|-80.847383|82|35.024464|CRAFT BEER|0.0|16|SHOCK TOP ALE 6PK|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00018200139864|DOMESTIC BEER|BEER|-81.027334|81.027393142178198|317|1
34.977331|b4594716340e35bbc95c0161815e3883091b62e2|7.89|2014-09-16 16:18:00|81.02739863253349|3|1910003108|149|35.014573965463335|0|14|3246|-80.847383|1020|35.024464|FACIAL CARE|0.0|17|BIORE ULTRA DEEP PORE STRIPS|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00019100031098|FACIAL CLEANSER & MOISTURIZER|HBC|-81.027334|81.027393142178198|317|1
34.977331|0cc5c18b3bfdd1256c1338af60b05b5536c3e65c|3.75|2014-11-29 17:17:00|81.02739863253349|3|1600048796|149|35.014573965463335|0|14|74|-80.847383|9|35.024464|RTE CEREAL ALL FAMILY|1.25|1|GM RICE CHEX|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00016000487949|CEREAL|G1 GROCERY|-81.027334|81.027393142178198|317|1
34.977331|000b982b52bbcf8c8c99468ff659af4dc5932302|1.78|2015-01-12 18:52:00|81.02739863253349|3||149|35.014573965463335|0|14|532|-80.847383|64|35.024464|FRESH CUCUMBERS|0.0|4|COO CUCUMBERS S/S|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00204062000002|FRESH PRODUCE|PRODUCE|-81.027334|81.027393142178198|317|2
34.977331|dbae31113a078de16053c0600f6c48e69f9a36fa|2.0|2014-09-15 19:19:00|81.02739863253349|3||149|35.014573965463335|0|14|500|-80.847383|64|35.024464|FRESH APPLES|0.0|4|RED DEL APPLE EASTERN|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00204168000005|FRESH PRODUCE|PRODUCE|-81.027334|81.027393142178198|317|1
34.977331|204348b2eca2695d848161e5cf158bcaedccbc9e|5.99|2014-11-08 12:15:00|81.02739863253349|3|8500001849|149|35.014573965463335|0|14|9944|-80.847383|885|35.024464|NFS POP OTHER RED|0.0|13|BAREFOOT SWEET RED|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00085000018491|POPULAR (4-$7.99)|WINE|-81.027334|81.027393142178198|317|1
34.977331|1edede5e1b69948d120fb359daa985aa76ed0fc3|2.85|2014-10-02 19:10:00|81.02739863253349|3|2580002320|149|35.014573965463335|0|14|1278|-80.847383|48|35.024464|SINGLE SERVE NUTRITIONAL|0.0|5|WW SMART ONES CHICKEN PARMESAN|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00025800023981|FROZEN MEALS|FROZEN|-81.027334|81.027393142178198|317|1
34.977331|7187a3093fa65b184c5f85575964e4e0724a2709|8.79|2014-10-09 18:10:00|81.02739863253349|3|9955508520|149|35.014573965463335|0|14|37|-80.847383|10|35.024464|PODS/CUPS/SINGLES|0.0|1|CARIBOU BLEND K-CUPS|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00099555089929|COFFEE|G1 GROCERY|-81.027334|81.027393142178198|317|1
34.977331|946922e8bd6ce00b113023a1d8d1c3fe01a6e95c|8.79|2014-10-01 16:31:00|81.02739863253349|3|9955508520|149|35.014573965463335|0|14|37|-80.847383|10|35.024464|PODS/CUPS/SINGLES|0.0|1|CARIBOU BLEND K-CUPS|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00099555089929|COFFEE|G1 GROCERY|-81.027334|81.027393142178198|317|1
34.977331|873a889fe7d45345ab71c246f83db9309f452584|1.99|2014-12-04 06:44:00|81.02739863253349|3|78616233800|149|35.014573965463335|0|14|31|-80.847383|4|35.024464|NON CARBONATED WATER|0.99|1|CB SMARTWATER 1 LTR PET SINGLE|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00786162338006|BOTTLED WATER|G1 GROCERY|-81.027334|81.027393142178198|317|1
34.977331|ea52b37a4c0f7e02ac8c120c1d9b3ab58299401e|3.99|2014-12-04 16:26:00|81.02739863253349|3|66559609990|149|35.014573965463335|0|14|326|-80.847383|54|35.024464|COOKIES/BROWNIES-REFRIGERATED|0.0|3|IMMACULATE BAKE GF CHOC CHUNK|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00665596099908|DOUGH PRODUCTS|DAIRY|-81.027334|81.027393142178198|317|1
34.977331|433000237f42c5cb9349049675dc4144d27d4160|5.99|2014-09-12 18:55:00|81.02739863253349|3|8500001444|149|35.014573965463335|0|14|9938|-80.847383|885|35.024464|NFS POP PINOT GRS/GRIGIO|0.0|13|CB-BAREFOOT PINOT GRIGIO|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00085000014448|POPULAR (4-$7.99)|WINE|-81.027334|81.027393142178198|317|1
34.977331|3eabf8d8d5900522ae2078f072990007c71b0792|7.89|2014-12-30 19:32:00|81.02739863253349|3|9955508205|149|35.014573965463335|0|14|37|-80.847383|10|35.024464|PODS/CUPS/SINGLES|0.0|1|EIGHT O'CLOCK HAZELNUT K-CUPS|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00099555082067|COFFEE|G1 GROCERY|-81.027334|81.027393142178198|317|1
34.977331|e29fffa5e2f84dd488fda645a5686dd548144f88|1.39|2014-09-14 15:05:00|81.02739863253349|3|1254667609|149|35.014573948188662|0|14|48|-80.8062|7|35.037115|REGISTER GUM|0.0|1|TRIDENT WHITE PEPPERMINT|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00012546676090|CANDY|G1 GROCERY|-81.027334|81.027407588011428|27|1
34.977331|87a4ad2887f8872419673b37b7660ca700bf3636|1.39|2014-09-27 14:42:00|81.02739863253349|3|1254667609|149|35.014573965463335|0|14|48|-80.847383|7|35.024464|REGISTER GUM|0.0|1|TRIDENT WHITE PEPPERMINT|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00012546676090|CANDY|G1 GROCERY|-81.027334|81.027393142178198|317|1
34.977331|3ea2df1db665acdae908beb536596605b5697459|3.5|2015-02-22 11:43:00|81.02739863253349|3|96824|149|35.014573965463335|0|14|1581|-80.847383|369|35.024464|NFS BEVERAGE BREWED|0.0|22|BREWED  COFFEE TALL.|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00000000968240|NFS STARBUCKS|COFFEE SHOP|-81.027334|81.027393142178198|317|2
34.977331|f992ec9a9ccebf63761f6a185c21b1c16f45f422|3.85|2014-09-20 18:08:00|81.02739863253349|3|3800001611|149|35.014573965463335|0|14|61|-80.847383|9|35.024464|RTE CEREAL ADULT|1.36|1|KELLOGG SPECIAL K 12 OZ BOX|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00038000016110|CEREAL|G1 GROCERY|-81.027334|81.027393142178198|317|1
34.977331|07db9c1d87b61250a162f3f3d5dfc33314c0cc87|2.99|2014-12-02 18:53:00|81.02739863253349|3|1570007200|149|35.014573965463335|0|14|1147|-80.847383|229|35.024464|HOT COCOA MIX|0.0|1|SWISS MISS NO SUGAR HOT COCOA|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00015700072004|COCOAS CREAMERS SYRUPS|G1 GROCERY|-81.027334|81.027393142178198|317|1
34.977331|728fb9cf960dd1126a8522d33ed13b092bd66e12|1.49|2015-02-06 06:38:00|81.02739863253349|3|7203670302|149|35.014573965463335|0|14|728|-80.847383|72|35.024464|NFS-PLASTIC FLATWARE|0.0|1|E  YH OCCASIONS FS SPOONS|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00072036703026|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-81.027334|81.027393142178198|317|1
34.977331|1dac95692aaf2565f02c5a95c43c2876893b9cb4|9.99|2014-11-26 12:48:00|81.02739863253349|3|7023666021|149|35.014573948188662|0|14|751|-80.8062|87|35.037115|NFS-BOUQUETS|0.0|9|LOVE IN BLOOM|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00070236660217|FLORAL|FLORAL|-81.027334|81.027407588011428|27|1
34.977331|ac0d7ebc3cf76349e999ff1562db4f128b9b805b|3.79|2015-02-27 15:31:00|81.02739863253349|3|4950800600|149|35.014573965463335|0|14|1981|-80.847383|480|35.024464|CHIPS|1.29|6|ORIGINAL PRETZEL CRISPS|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00049508006008|DRY GOODS|DELI|-81.027334|81.027393142178198|317|1
34.977331|30129382b1d4a67a2026ad844a9dba4a74a2a1fd|5.35|2014-12-26 19:58:00|81.02739863253349|3|3700041759|149|35.014573965463335|0|14|388|-80.847383|66|35.024464|NFS-DISHWASH PWDR/LIQUID|1.06|1|CASCADE DAWN FRESH SCENT 20CT|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00037000417590|DETERGENTS|G1 GROCERY|-81.027334|81.027393142178198|317|1
34.977331|fc2f318c4c0ac1f7a00bb536009685d0b58d514a|2.67|2015-01-15 19:00:00|81.02739863253349|3|7203698754|149|35.014573935960946|0|14|1265|-80.816172|57|35.059823|ALMOND MILK|0.0|3|HT ALMOND DRINK UNSWT VANILLA|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00072036987563|MILK|DAIRY|-81.027334|81.027416294623393|66|1
34.977331|4bebd8c83aed65650b7a3caf19d9cdeac190199d|3.15|2015-03-03 06:40:00|81.02739863253349|3|7265500105|149|35.014573965463335|0|14|1278|-80.847383|48|35.024464|SINGLE SERVE NUTRITIONAL|0.0|5|HC CAFE STEAMERS CHKN MARINARA|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00072655001015|FROZEN MEALS|FROZEN|-81.027334|81.027393142178198|317|1
34.977331|498a930f2c44e58f4d9fd24e0467b6e559e2c314|3.69|2014-10-29 16:35:00|81.02739863253349|3|38151905501|149|35.014573965463335|0|14|3530|-80.847383|1045|35.024464|SHAMPOO-MID PRICE|0.7|17|HERBAL ESS SHAM COLOR ME HAPPY|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00381519055058|HAIR & SCALP CARE|HBC|-81.027334|81.027393142178198|317|1
34.977331|ac789ffef7edc1c48f3f69a393989aa51145771e|3.69|2014-11-23 16:32:00|81.02739863253349|3|38151905501|149|35.014573965463335|0|14|3530|-80.847383|1045|35.024464|SHAMPOO-MID PRICE|0.7|17|HERBAL ESS SHAM COLOR ME HAPPY|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00381519055058|HAIR & SCALP CARE|HBC|-81.027334|81.027393142178198|317|1
34.977331|2fabc5c57c8ebf86034fd8c6080f855563d2b5d6|4.15|2014-11-22 17:29:00|81.02739863253349|3|980089500|149|35.014573965463335|0|14|1435|-80.847383|19|35.024464|SHELF STABLE SPREADS|1.15|1|NUTELLA HAZELNUT SPREAD|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00009800895007|JAMS/JELLIES/SPREADS|G1 GROCERY|-81.027334|81.027393142178198|317|1
34.977331|3028f4085af207cf0cc160361d43d8ba85b8fb06|1.2|2014-09-12 06:25:00|81.02739863253349|3|3663203732|149|35.014573965463335|0|14|685|-80.847383|61|35.024464|GREEK|0.0|3|DANNON LNF GREEK STRAWBERRY|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00036632037312|YOGURT|DAIRY|-81.027334|81.027393142178198|317|1
34.977331|ec4fa2bcbb113d2bcbd7525140a02d7984f6fe6e|1.2|2015-02-25 08:04:00|81.02739863253349|3|3663203732|149|35.014573965463335|0|14|685|-80.847383|61|35.024464|GREEK|0.2|3|DANNON LNF GREEK STRAWBERRY|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00036632037312|YOGURT|DAIRY|-81.027334|81.027393142178198|317|1
34.977331|702961bc359799efc0b2e21a9b6fddf2c26d2fcf|5.98|2015-03-05 16:09:00|81.02739863253349|3|4300002825|149|35.014573965463335|0|14|121|-80.847383|20|35.024464|ASEPTIC JUICES|0.98|1|KOOLAID JAMMERS TROP/PUNCH|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00043000028254|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-81.027334|81.027393142178198|317|2
34.977331|a7686f8feb64583ffa7915268f4c80396f79c3b4|2.1|2014-10-28 06:36:00|81.02739863253349|3|96825|149|35.014573965463335|0|14|1581|-80.847383|369|35.024464|NFS BEVERAGE BREWED|0.0|22|BREWED COFFEE GRANDE|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00000000968250|NFS STARBUCKS|COFFEE SHOP|-81.027334|81.027393142178198|317|1
34.977331|de0304d9d051c431b139b121dfc9e2a16085133a|2.69|2014-10-19 19:11:00|81.02739863253349|3|7203663996|149|35.014573965463335|0|14|342|-80.847383|57|35.024464|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|0c25962eb9bc8cce1ac1e782fce57b6e697ed354|2.573401152459771|35.014943729270243|00072036631299|MILK|DAIRY|-81.027334|81.027393142178198|317|1
35.23102|3262f1f711e030ee92fbefb5ba014e041226ebf4|6.69|2014-11-25 10:16:00|1.4094857484078087|4|7790050209|205|0.6148972978359727|0|26|1271|-80.8438|41|35.23102|PROTEIN BREAKFAST|0.0|5|J D SAUS/EGG/CHS CROSSIANT 4CT|1324b55b17c59430c753c3944b7cc6592e2157f3|0.4218690723014831|0.61471665291522548|00077900502101|BREAKFAST FOODS FROZEN|FROZEN|-80.8438|1.4109904898237917|205|1
35.23102|f6155ebfd26f44d642e50af8265ea057e58d8362|6.69|2015-01-21 13:12:00|1.4094857484078087|4|7790050209|205|0.6148972978359727|0|26|1271|-80.8438|41|35.23102|PROTEIN BREAKFAST|0.0|5|J D SAUS/EGG/CHS CROSSIANT 4CT|1324b55b17c59430c753c3944b7cc6592e2157f3|0.4218690723014831|0.61471665291522548|00077900502101|BREAKFAST FOODS FROZEN|FROZEN|-80.8438|1.4109904898237917|205|1
35.23102|f8eedab555e62c9ad259fefdb8b3228dd9a0eba0|6.69|2014-12-22 16:58:00|1.4094857484078087|4|7790050209|205|0.6148972978359727|0|26|1271|-80.8438|41|35.23102|PROTEIN BREAKFAST|0.0|5|J D SAUS/EGG/CHS CROSSIANT 4CT|1324b55b17c59430c753c3944b7cc6592e2157f3|0.4218690723014831|0.61471665291522548|00077900502101|BREAKFAST FOODS FROZEN|FROZEN|-80.8438|1.4109904898237917|205|1
35.23102|b7d50c21ff69922ba8a0ce11d1a24fc629b95959|2.29|2014-09-30 10:47:00|1.4094857484078087|4|1200000410|205|0.6148972978359727|0|26|854|-80.8438|32|35.23102|LIQUID ICED COFFEES|0.0|1|STARBUCKS FRAPPUCCINO VANILLA|1324b55b17c59430c753c3944b7cc6592e2157f3|0.4218690723014831|0.61471665291522548|00012000004100|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.8438|1.4109904898237917|205|1
35.23102|c91914b8e1acccba3a9912b08d7db01e56ce93ab|2.29|2014-09-27 21:30:00|1.4094857484078087|4|1200000410|205|0.6148972978359727|0|26|854|-80.8438|32|35.23102|LIQUID ICED COFFEES|0.0|1|STARBUCKS FRAPPUCCINO VANILLA|1324b55b17c59430c753c3944b7cc6592e2157f3|0.4218690723014831|0.61471665291522548|00012000004100|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.8438|1.4109904898237917|205|1
35.23102|bf0a14ca210ab3ffe42defaef5b73176e18e5b27|3.35|2015-02-22 20:53:00|1.4094857484078087|4|1312000286|205|0.6148972978359727|0|26|1469|-80.8438|278|35.23102|REGULAR CUT FRIES|0.0|5|ORE-IDA CTRY STYLE HASH BROWNS|1324b55b17c59430c753c3944b7cc6592e2157f3|0.4218690723014831|0.61471665291522548|00013120008337|FROZEN POTATO|FROZEN|-80.8438|1.4109904898237917|205|1
35.23102|4a6c88c1d025bb1ce247679a75ddf39630f8da1d|3.75|2015-01-09 20:10:00|1.4094857484078087|4|1600048796|205|0.6148972978359727|0|26|74|-80.8438|9|35.23102|RTE CEREAL ALL FAMILY|0.0|1|GM HONEY NUT CHEX|1324b55b17c59430c753c3944b7cc6592e2157f3|0.4218690723014831|0.61471665291522548|00016000487925|CEREAL|G1 GROCERY|-80.8438|1.4109904898237917|205|1
35.23102|cf3fcb7b4ca2ab7a44b391636334bf61de95be52|1.57|2014-12-21 15:23:00|1.4094857484078087|4|7203661018|205|0.6148972978359727|0|26|221|-80.8438|34|35.23102|SALT SALT SUBSTITUTES|0.0|1|HT GARLIC SALT|1324b55b17c59430c753c3944b7cc6592e2157f3|0.4218690723014831|0.61471665291522548|00072036610188|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.8438|1.4109904898237917|205|1
35.23102|ca5093197ddc6414585a18bfdfdb59f0dadcbb39|3.29|2015-02-21 15:25:00|1.4094857484078087|4|7203698555|205|0.6148972978359727|0|26|427|-80.8438|72|35.23102|NFS-TOILET TISSUE|0.5|1|HT 1000 SHEET BATHTISSUE 4 RL|1324b55b17c59430c753c3944b7cc6592e2157f3|0.4218690723014831|0.61471665291522548|00072036985552|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.8438|1.4109904898237917|205|1
35.23102|42a0eb4f1822f3e7496ec73c2a7bbd1bef43ff8d|2.69|2015-02-17 21:55:00|1.4094857484078087|4|1380016610|205|0.6148972978359727|0|26|1278|-80.8438|48|35.23102|SINGLE SERVE NUTRITIONAL|0.19|5|LC STEAK TIPS PORTABELLO|1324b55b17c59430c753c3944b7cc6592e2157f3|0.4218690723014831|0.61471665291522548|00013800156501|FROZEN MEALS|FROZEN|-80.8438|1.4109904898237917|205|1
35.23102|d245b4cc120e29dd4d33f7f18c8687f2ededcac1|4.49|2015-01-16 21:30:00|1.4094857484078087|4|85804600400|205|0.6148972978359727|0|26|1279|-80.8438|48|35.23102|SINGLE SERVE FLAVOR|0.0|5|MOMMA B CKN ALFREDO|1324b55b17c59430c753c3944b7cc6592e2157f3|0.4218690723014831|0.61471665291522548|00858046004083|FROZEN MEALS|FROZEN|-80.8438|1.4109904898237917|205|1
35.23102|40baf816175f70e2df47cf386b5e66630ab364d9|2.63|2014-09-26 20:33:00|1.4094857484078087|4||205|0.6148972978359727|0|26|505|-80.8438|64|35.23102|FRESH SOFT FRUIT|0.0|4|EASTERN PEACHES|1324b55b17c59430c753c3944b7cc6592e2157f3|0.4218690723014831|0.61471665291522548|00204403000005|FRESH PRODUCE|PRODUCE|-80.8438|1.4109904898237917|205|1
35.23102|229c5069e350f6cd238a002c29cc65e2d5911d73|1.79|2015-01-21 13:15:00|1.4094857484078087|4|8079380770|205|0.6148972978359727|0|26|99|-80.8438|32|35.23102|LIQUID TEA|0.0|1|D FUZE SLENDER TROPICAL PUNCH|1324b55b17c59430c753c3944b7cc6592e2157f3|0.4218690723014831|0.61471665291522548|00080793807765|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.8438|1.4109904898237917|205|1
35.23102|734a9556d326a026a28bd20b211a43a992d05277|4.29|2014-10-02 14:40:00|1.4094857484078087|4|2840015938|205|0.6148972978359727|0|26|201|-80.8438|31|35.23102|POTATO CHIPS|0.0|1|RUFFLES ULTIMATE BCN CHED SKIN|1324b55b17c59430c753c3944b7cc6592e2157f3|0.4218690723014831|0.61471665291522548|00028400208949|SNACKS|G1 GROCERY|-80.8438|1.4109904898237917|205|1
35.23102|2b65b4e16cf3b6d76275d1eb0637bd44023ebe5c|3.99|2014-09-30 10:46:00|1.4094857484078087|4|75491808201|205|0.6148972978359727|0|26|197|-80.8438|31|35.23102|POPPED POPCORN|0.0|1|POPPYCOCK ORIGINAL|1324b55b17c59430c753c3944b7cc6592e2157f3|0.4218690723014831|0.61471665291522548|00754918082015|SNACKS|G1 GROCERY|-80.8438|1.4109904898237917|205|1
35.603432|3636dc4b1b7b162dacf0bbd7757649e77fbc2b43|5.29|2014-10-30 17:50:00|80.891462859624312|4|5209220388|274|35.647045933837617|0|45|5827|-80.875654|1536|35.585842|FOILWARE CASSEROLE|1.06|18|CNC GIANT ALL PURPOSE PAN/LID|14497c7397bdafc5c997b3d6157d59910f6a06d5|3.0136175176124556|35.636605227883024|00052092203883|FOILWARE|GM|-80.895009|80.895014043343394|99|1
35.603432|ac4b1310ffc5773de74d77c51898afe4f09bfb6b|14.99|2014-10-02 11:11:00|80.891462859624312|4|1820053218|274|35.647045933837617|0|45|455|-80.875654|82|35.585842|DOMESTIC PREMIUM 12PK&>|0.0|16|BUD LIGHT 18PK 12OZ CAN|14497c7397bdafc5c997b3d6157d59910f6a06d5|3.0136175176124556|35.636605227883024|00018200532184|DOMESTIC BEER|BEER|-80.895009|80.895014043343394|99|1
35.603432|b3f736ed02df42b6bc2ca5df56f7a7ccb8bce5de|5.96|2014-12-19 15:27:00|80.891462859624312|4|3890000473|274|35.647045933837617|0|45|115|-80.875654|16|35.585842|REMAINING FRUIT|0.96|1|DOLE PINEAPPLE 20 CHUNKS JC.|14497c7397bdafc5c997b3d6157d59910f6a06d5|3.0136175176124556|35.636605227883024|00038900004736|FRUIT-CAN/JAR|G1 GROCERY|-80.895009|80.895014043343394|99|4
35.603432|bf38b049bce3293647281aea35636eb74461d56f|3.25|2014-11-13 11:10:00|80.891462859624312|4|7203656080|274|35.647045933837617|0|45|318|-80.875654|52|35.585842|SHREDDED/GRATED CHEESE|3.25|3|HT SHRED SHARP CHED CHEESE 2%|14497c7397bdafc5c997b3d6157d59910f6a06d5|3.0136175176124556|35.636605227883024|00072036590466|CHEESE|DAIRY|-80.895009|80.895014043343394|99|1
35.603432|2b3cb1e97d42926769f0fb8b218e2005ac564e23|21.98|2014-10-30 14:19:00|80.891462859624312|4|7203683001|274|35.647045933837617|0|45|352|-80.875654|110|35.585842|IQF CHICKEN|5.5|19|HT 2.5 LB CHICKEN TENDR BRST|14497c7397bdafc5c997b3d6157d59910f6a06d5|3.0136175176124556|35.636605227883024|00072036830029|FROZEN CASE MEAT|CASE READY MEATS|-80.895009|80.895014043343394|99|2
35.603432|fe9c09286aa500fba0ad9a18644998c425804917|25.38|2014-11-24 14:19:00|80.891462859624312|4|20009200000|274|35.647045933837617|0|45|974|-80.875654|201|35.585842|FRESH TURKEY|6.36|2|BUTTERBALL FRSH TURKEY BREAST|14497c7397bdafc5c997b3d6157d59910f6a06d5|3.0136175176124556|35.636605227883024|00200092000005|POULTRY|MEAT|-80.895009|80.895014043343394|99|1
35.603432|c2965c8fde545aaf8da4819c5ceb55cf463fb201|4.99|2015-01-16 12:12:00|80.891462859624312|4|7336070341|274|35.647045933837617|0|45|30|-80.875654|4|35.585842|CARBONATED WATER|1.49|1|LACROIX WTR GRPEFRT 12PK|14497c7397bdafc5c997b3d6157d59910f6a06d5|3.0136175176124556|35.636605227883024|00012993102012|BOTTLED WATER|G1 GROCERY|-80.895009|80.895014043343394|99|1
35.603432|6edfd08ae932caa9b4a58c3e2a6dd7dbd03abfc8|6.43|2015-02-25 13:20:00|80.891462859624312|4|20169200000|274|35.647045933837617|0|45|297|-80.875654|49|35.585842|GROUND BEEF|0.0|2|GROUND BEEF 96% LEAN|14497c7397bdafc5c997b3d6157d59910f6a06d5|3.0136175176124556|35.636605227883024|00201692000006|BEEF|MEAT|-80.895009|80.895014043343394|99|1
35.603432|b2eef5a05994e892054cf7b7b9349f54f6812a13|2.79|2015-01-29 14:08:00|80.891462859624312|4|4127800005|274|35.647045933837617|0|45|221|-80.875654|34|35.585842|SALT SALT SUBSTITUTES|1.3|1|JANES KRAZY MIXED UP SALT|14497c7397bdafc5c997b3d6157d59910f6a06d5|3.0136175176124556|35.636605227883024|00041278000057|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.895009|80.895014043343394|99|1
35.603432|7262fa6582eb5405410fb58fe0a2225f84dfa4b6|13.58|2014-09-20 12:28:00|80.891462859624312|4|4900002890|274|35.647045933837617|0|45|54|-80.875654|8|35.585842|DIET|3.4|23|DIET COKE 12OZ 12PK FRIDGE CAN|14497c7397bdafc5c997b3d6157d59910f6a06d5|3.0136175176124556|35.636605227883024|00049000028911|CARBONATED BEVERAGES|BEVERAGE|-80.895009|80.895014043343394|99|2
35.603432|0cb0fb4fd07e15095ceff522e10748912ae16b2d|4.78|2014-12-29 14:25:00|80.891462859624312|4|7342000011|274|35.647045933837617|0|45|322|-80.875654|53|35.585842|SOUR CREAM|0.78|3|DAISY LIGHT SOUR CREAM|14497c7397bdafc5c997b3d6157d59910f6a06d5|3.0136175176124556|35.636605227883024|00073420000158|CULTURES|DAIRY|-80.895009|80.895014043343394|99|2
35.603432|b12d4d27aaee7107d9a3cf644617fc62ed7b3e96|13.98|2015-03-05 21:12:00|80.891462859624312|4|4900002890|274|35.647045933837617|0|45|54|-80.875654|8|35.585842|DIET|3.5|23|FRESCA 12OZ 12PK FRIDGEPACK CN|14497c7397bdafc5c997b3d6157d59910f6a06d5|3.0136175176124556|35.636605227883024|00049000031058|CARBONATED BEVERAGES|BEVERAGE|-80.895009|80.895014043343394|99|2
35.323246|199e34f88df3f6164678042934fa79fa1d471bff|14.7|2014-09-14 15:01:00|1.4102725052409182|4|3040077377|166|0.6165069451919168|0|1|427|-80.945176|72|35.323246|NFS-TOILET TISSUE|2.72|1|ANGEL SOFT SOFT/STRONG 12DR|14c6ed8bd59d63a74fc39a74f553b840ec5879d8|2.4606716167626996|0.61833652052202714|00030400773778|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.945176|1.4127598348062935|166|2
35.323246|040e075b5057a1c26718611c1725fc80d58f156b|4.29|2014-11-26 07:41:00|80.945255278477163|4|2840016014|166|35.35885744302513|0|13|201|-80.848528|31|35.053394|POTATO CHIPS|2.15|1|LAYS BBQ|14c6ed8bd59d63a74fc39a74f553b840ec5879d8|2.4606716167626996|35.37387923947206|00028400160131|SNACKS|G1 GROCERY|-80.945176|80.945279402759297|11|1
35.323246|5788c149be0babc4b5eaff7a847d2383fe1bd5f7|14.97|2015-02-07 16:55:00|1.4102725052409182|4|6827493471|166|0.6165069451919168|0|1|31|-80.945176|4|35.323246|NON CARBONATED WATER|6.0|1|NESTLE PURE LIFE .5L 24PK|14c6ed8bd59d63a74fc39a74f553b840ec5879d8|2.4606716167626996|0.61833652052202714|00068274934711|BOTTLED WATER|G1 GROCERY|-80.945176|1.4127598348062935|166|3
35.323246|6ae84ca12a5398a50b80d40a737bc17c9b8ecc30|9.98|2014-11-15 14:28:00|1.4102725052409182|4|6827493471|166|0.6165069451919168|0|1|31|-80.945176|4|35.323246|NON CARBONATED WATER|1.2|1|NESTLE PURE LIFE .5L 24PK|14c6ed8bd59d63a74fc39a74f553b840ec5879d8|2.4606716167626996|0.61833652052202714|00068274934711|BOTTLED WATER|G1 GROCERY|-80.945176|1.4127598348062935|166|2
35.323246|8d6a3cc4ee79fff2df972e6e22bc229f27119191|4.99|2015-01-18 18:40:00|1.4102725052409182|4|6827493471|166|0.6165069451919168|0|1|31|-80.945176|4|35.323246|NON CARBONATED WATER|2.0|1|NESTLE PURE LIFE .5L 24PK|14c6ed8bd59d63a74fc39a74f553b840ec5879d8|2.4606716167626996|0.61833652052202714|00068274934711|BOTTLED WATER|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|87d259f5a1567a64a423261f8d4382cd6eafd2a0|4.99|2015-02-15 17:38:00|1.4102725052409182|4|6827493471|166|0.6165069451919168|0|1|31|-80.945176|4|35.323246|NON CARBONATED WATER|1.0|1|NESTLE PURE LIFE .5L 24PK|14c6ed8bd59d63a74fc39a74f553b840ec5879d8|2.4606716167626996|0.61833652052202714|00068274934711|BOTTLED WATER|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|1e76f8754766130c585dd0215844255585a3f843|4.99|2014-11-24 17:34:00|80.945255278477163|4|20165500000|166|35.35885744302513|0|13|297|-80.848528|49|35.053394|GROUND BEEF|0.0|2|HT PREMIUM GRND BEEF 80% LEAN|14c6ed8bd59d63a74fc39a74f553b840ec5879d8|2.4606716167626996|35.37387923947206|00201655000005|BEEF|MEAT|-80.945176|80.945279402759297|11|1
35.323246|199181fb7afb80473c651de5a9f31d67afb5d6a7|30.67|2014-12-31 13:13:00|80.945255278477163|4|20926400000|166|35.35885744302513|0|13|668|-80.848528|146|35.053394|LEGS/CLUSTERS|12.280000000000001|12|PRE BAGGED SNOW CRAB CLUSTERS|14c6ed8bd59d63a74fc39a74f553b840ec5879d8|2.4606716167626996|35.37387923947206|00209264000003|CRAB|SEAFOOD|-80.945176|80.945279402759297|11|2
35.323246|630b8558698e04446e3082181dfdc7cca0141030|4.58|2015-01-31 20:26:00|1.4102725052409182|4|7203663996|166|0.6165069451919168|0|1|342|-80.945176|57|35.323246|FRESH MILK|0.82|3|HARRIS TEETER 2%   MILK|14c6ed8bd59d63a74fc39a74f553b840ec5879d8|2.4606716167626996|0.61833652052202714|00072036639998|MILK|DAIRY|-80.945176|1.4127598348062935|166|2
35.323246|ad195111bf08a9c3e5a6c8615d168b242239b069|21.98|2014-12-14 18:02:00|1.4102725052409182|4|3040077569|166|0.6165069451919168|0|1|427|-80.945176|72|35.323246|NFS-TOILET TISSUE|5.0|1|ANGEL SOFT SOFT/STRONG 16R|14c6ed8bd59d63a74fc39a74f553b840ec5879d8|2.4606716167626996|0.61833652052202714|00030400775697|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.945176|1.4127598348062935|166|2
35.323246|8fe50d3d01ee98b372e3aae33bde3e8babcd903c|7.94|2014-12-14 18:08:00|1.4102725052409182|4|3040077569|166|0.6165069451919168|0|1|427|-80.945176|72|35.323246|NFS-TOILET TISSUE|0.0|1|ANGEL SOFT SOFT/STRONG 16R|14c6ed8bd59d63a74fc39a74f553b840ec5879d8|2.4606716167626996|0.61833652052202714|00030400775697|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.945176|1.4127598348062935|166|2
35.323246|7e35867dfdbac567402a75600203a6fecc4ea7ab|3.99|2014-09-27 19:17:00|80.945255278477163|4|7203663995|166|35.358857538486085|0|13|342|-80.8438|57|35.23102|FRESH MILK|1.02|3|HARRIS TEETER 2% MILK|14c6ed8bd59d63a74fc39a74f553b840ec5879d8|2.4606716167626996|35.37387923947206|00072036639981|MILK|DAIRY|-80.945176|80.945197777645774|205|1
35.323246|ec74de7f994eff15ea49558b6b6367c540d59aeb|12.99|2015-01-15 07:41:00|80.945255278477163|4|7023666348|166|35.35885744302513|0|13|751|-80.848528|87|35.053394|NFS-BOUQUETS|0.0|9|$12.99 SIMPLY ELEGANT BOUQUET|14c6ed8bd59d63a74fc39a74f553b840ec5879d8|2.4606716167626996|35.37387923947206|00070236663485|FLORAL|FLORAL|-80.945176|80.945279402759297|11|1
35.323246|7ab156c4ce85064c8eb7402ed41ec8895d41ca23|4.3|2015-01-06 18:07:00|1.4102725052409182|4|7142909849|166|0.6165069451919168|0|1|238|-80.945176|38|35.323246|RICE FLAVORED|0.16|1|ZAT RICE JAMBALAYA MIX.|14c6ed8bd59d63a74fc39a74f553b840ec5879d8|2.4606716167626996|0.61833652052202714|00071429095236|RICE GRAINS AND BEANS|G1 GROCERY|-80.945176|1.4127598348062935|166|2
35.17335|fd6e2f94679e9bfd11c35c3ccc69d5f92707e476|5.78|2014-12-17 19:52:00|80.709059419360486|2|7203663102|174|35.18473217051357|0|31|339|-80.654118|57|35.123768|EGGNOGS/DRINKS|1.78|3|I/O HARRIS TEETER EGG NOG|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|35.187384292804154|00072036631022|MILK|DAIRY|-80.70901|80.709013723936394|473|2
35.17335|2d589514ac1894221977987c5a662b226fd7e185|2.89|2015-01-14 19:13:00|1.4094857484078087|2|7203655029|174|0.6138907664563474|0|26|331|-80.70901|52|35.17335|NATURAL SLICED|1.22|3|HT SLICED MUENSTER CHEESE|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00072036600387|CHEESE|DAIRY|-80.70901|1.4086379605250285|174|1
35.17335|955d022dadbe8a8adcd7e8c11a0ba04028d1596b|2.89|2015-01-25 18:07:00|1.4094857484078087|2|7203655029|174|0.6138907664563474|0|26|331|-80.70901|52|35.17335|NATURAL SLICED|0.0|3|HT SLICED MUENSTER CHEESE|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00072036600387|CHEESE|DAIRY|-80.70901|1.4086379605250285|174|1
35.17335|e3933cfecac29dcbaef8b8f954a8d16b4e7c3e8b|3.39|2014-12-23 21:54:00|1.4094857484078087|2|7102231552|174|0.6138907664563474|0|26|117|-80.70901|17|35.17335|DRIED REMAINING FRUIT|1.7|1|MARIANI CRANBERRIES|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00071022315526|FRUIT-DRIED|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|7cef5f771e054a80a5a5fc9685b897e2f2c61be4|4.15|2014-12-01 17:16:00|1.4094857484078087|2|4400000488|174|0.6138907664563474|0|26|89|-80.70901|12|35.17335|GRAHAM CRACKERS|0.65|1|HONEYMAID GRAHAMS|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00044000004637|COOKIES|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|b42939dfc553b536120ff19e0c0bae6335f2d4cb|3.99|2014-10-10 13:36:00|1.4094857484078087|2|4157005982|174|0.6138907664563474|0|26|1148|-80.70901|21|35.17335|ALMONDS|0.99|1|BLUE DIAM HNY RST ALMONDS CAN|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00041570072561|NUTS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|a5fd809a7e65b8819ea14c3eb6493f68dc81dca7|4.89|2014-10-28 19:53:00|1.4094857484078087|2|3700084609|174|0.6138907664563474|0|26|3592|-80.70901|1050|35.17335|HAIR STYLING HAIR SPRAY|1.4|17|VS FLEXIBLE HOLD HAIR SPRAY|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00037000846925|HAIR STYLING|HBC|-80.70901|1.4086379605250285|174|1
35.17335|46823b7d8ca5189da74f031a14f203e39868487f|3.99|2014-10-19 20:01:00|80.709059419360486|2|4000015140|174|35.184732164768299|0|31|46|-80.64817|7|35.04711|PKG CHOC|0.49|1|3 MUSKETEER FUN SIZE|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|35.187384292804154|00040000151227|CANDY|G1 GROCERY|-80.70901|80.709024478830585|129|1
35.17335|b29b03f20d8700b8dfa4fb7818506cc1a9121b97|3.79|2014-09-23 21:13:00|1.4094857484078087|2|4000047070|174|0.6138907664563474|0|26|46|-80.70901|7|35.17335|PKG CHOC|0.0|1|M&M MILK CHOCOLATE|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00040000470700|CANDY|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|418df222c2d6179563fa4d901df2ea8353ce110e|4.69|2014-11-06 20:55:00|80.709059419360486|2|3700088763|174|35.184732169464603|0|31|393|-80.709466|68|35.124987|NFS-AIR FRESHENERS|0.0|1|FEBREZE AE HVY DUTY CRISP CLN|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|35.187384292804154|00037000887669|FRESHENERS/DEODORIZERS|G1 GROCERY|-80.70901|80.709017043522778|157|1
35.17335|36c7ae32d516d208ae3495be85c26fed11790152|2.99|2014-12-26 20:50:00|1.4094857484078087|2|8630221549|174|0.6138907664563474|0|26|7422|-80.70901|1600|35.17335|CHRISTMAS BOWS|2.24|18|"I/O6"" CONFETTI BOWS HDAY COLOR"|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00086302215496|SEASONAL MERCHANDISE|GM|-80.70901|1.4086379605250285|174|1
35.17335|75a8f703d61e84ff6bde3ad4b281eb9f2d44bb0b|3.94|2014-11-13 17:22:00|80.709059419360486|2|7203695946|174|35.184732169464603|0|31|1295|-80.709466|383|35.124987|PIES PASTRY CASE TAX|0.0|14|"9"" CHOCOLATE SILK PIE"|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|35.187384292804154|00072036959461|PASTRY CASE|BAKERY|-80.70901|80.709017043522778|157|2
35.17335|34235f2a486766daecad8a81d102fa1f4bb90c2a|2.19|2015-01-13 19:19:00|80.709059419360486|2|7418226090|174|35.184732169464603|0|31|722|-80.709466|73|35.124987|NFS-HAND SOAPS|1.19|1|SS HAND COUNTRY DESIGNS|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|35.187384292804154|00074182260125|PERSONAL SOAP/BATH ADDITIVES|G1 GROCERY|-80.70901|80.709017043522778|157|1
35.17335|f9cfc51d8ade9b9ab61a6311f702a72e88280993|6.7|2014-09-28 17:33:00|80.709059419360486|2|7203656080|174|35.184732167794387|0|31|318|-80.825175|52|35.152722|SHREDDED/GRATED CHEESE|2.58|3|HT FANCY SHRED MEXICAN CHEESE|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|35.187384292804154|00072036590442|CHEESE|DAIRY|-80.70901|80.709020321020603|160|2
35.17335|ac5b51f0929170a873689ecf38e98c5cc276faf4|6.5|2015-03-05 18:58:00|1.4094857484078087|2|7203656080|174|0.6138907664563474|0|26|318|-80.70901|52|35.17335|SHREDDED/GRATED CHEESE|0.0|3|HT FANCY SHRED MEXICAN CHEESE|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00072036590442|CHEESE|DAIRY|-80.70901|1.4086379605250285|174|2
35.17335|648e67d5e083d4a9461082978807ea03250a2534|27.56|2014-12-13 17:32:00|1.4094857484078087|2|3040077377|174|0.6138907664563474|0|26|427|-80.70901|72|35.17335|NFS-TOILET TISSUE|3.6|1|ANGEL SOFT SOFT/STRONG 12DR|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00030400773778|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.70901|1.4086379605250285|174|4
35.17335|af0bd06def1b070792d72492f3a3ce058502100d|3.98|2014-10-21 21:09:00|80.709059419360486|2|2920000307|174|35.184732169464603|0|31|149|-80.709466|23|35.124987|WHSE PASTA CORE|1.98|1|MUELLER FETTUCCINE|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|35.187384292804154|00029200002058|PASTA|G1 GROCERY|-80.70901|80.709017043522778|157|2
35.17335|ad89646b38058d50417f4dade2b19852c2fcb963|2.29|2015-02-14 18:56:00|80.709059419360486|2|2670012915|174|35.184732164768299|0|31|1267|-80.64817|53|35.04711|DIPS AND SPREADS|0.79|3|DEAN'S FRENCH ONION DIP|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|35.187384292804154|00026700129155|CULTURES|DAIRY|-80.70901|80.709024478830585|129|1
35.17335|7f620f9b1bc9f38deae9fb051c6fa3676225c4e0|3.29|2015-01-17 19:01:00|1.4094857484078087|2|2840004768|174|0.6138907664563474|0|26|202|-80.70901|31|35.17335|PRETZELS|1.65|1|ROLD GOLD PRETZEL TINY TWIST|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00028400047685|SNACKS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|c69e2d59cad34ae31f42e0f25642b825442df3f4|3.79|2015-01-10 22:16:00|1.4094857484078087|2|2100062503|174|0.6138907664563474|0|26|318|-80.70901|52|35.17335|SHREDDED/GRATED CHEESE|1.29|3|KRAFT 2% MEXICAN FOUR CHEESE|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00021000024612|CHEESE|DAIRY|-80.70901|1.4086379605250285|174|1
35.17335|ce1baec7f4d35639a4fe70829842fe46cf85f6a6|7.38|2014-11-25 18:58:00|1.4094857484078087|2|2100062503|174|0.6138907664563474|0|26|318|-80.70901|52|35.17335|SHREDDED/GRATED CHEESE|1.84|3|KRAFT 2% MEXICAN FOUR CHEESE|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00021000024612|CHEESE|DAIRY|-80.70901|1.4086379605250285|174|2
35.17335|abee5417db320e8fec39fc3b11cf10ffe82b4df8|7.38|2014-11-23 19:10:00|1.4094857484078087|2|2100062503|174|0.6138907664563474|0|26|318|-80.70901|52|35.17335|SHREDDED/GRATED CHEESE|1.84|3|KRAFT 2% MEXICAN FOUR CHEESE|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00021000024612|CHEESE|DAIRY|-80.70901|1.4086379605250285|174|2
35.17335|82fbf18c5ed5abe9b3eacf05cda145756a15068d|7.58|2015-01-30 21:57:00|1.4094857484078087|2|2100062503|174|0.6138907664563474|0|26|318|-80.70901|52|35.17335|SHREDDED/GRATED CHEESE|1.89|3|KRAFT 2% MEXICAN FOUR CHEESE|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00021000024612|CHEESE|DAIRY|-80.70901|1.4086379605250285|174|2
35.17335|2a8b16fb15e27f94d4b62206aea025aca560506b|2.49|2014-11-03 19:32:00|1.4094857484078087|2|4137620228|174|0.6138907664563474|0|26|727|-80.70901|7|35.17335|SEASONAL CANDY-SINGLE FAC|1.25|1|I/O(H14)KRABBY PATTIES|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00041376202285|CANDY|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|13555212a7366e47f5e2f11766c08498eebfafe5|1.39|2015-02-19 21:23:00|1.4094857484078087|2|5210076069|174|0.6138907664563474|0|26|80|-80.70901|34|35.17335|SEASONING PACKETS|0.0|1|MC GRILL MATES MESQUITE MARNDE|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00052100025780|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|1cd3260a15d909115597f25526e0140a31d3702f|3.87|2015-02-25 19:15:00|1.4094857484078087|2|4800000245|174|0.6138907664563474|0|26|190|-80.70901|29|35.17335|TUNA-CANNED|0.8699999999999999|1|COS TUNA CHUNK LIGHT|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00048000002457|SEAFOOD-CANNED|G1 GROCERY|-80.70901|1.4086379605250285|174|3
35.17335|9460e36809b17e33b3b70e0779a444bb72125586|4.69|2014-11-09 18:17:00|1.4094857484078087|2|4900002468|174|0.6138907664563474|0|26|54|-80.70901|8|35.17335|DIET|2.35|23|DIET COKE .5 LITER/6 PK.|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.70901|1.4086379605250285|174|1
35.17335|be3046ed62087530e6ed2353993298ce4c2f57bb|24.950000000000003|2015-01-07 21:56:00|1.4094857484078087|2|4900002468|174|0.6138907664563474|0|26|54|-80.70901|8|35.17335|DIET|14.950000000000001|23|DIET COKE .5 LITER/6 PK.|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.70901|1.4086379605250285|174|5
35.17335|4cc877a76196e7d9088646f0eaf0be2fdbcd7ea1|1.99|2014-12-30 20:35:00|1.4094857484078087|2|7069027166|174|0.6138907664563474|0|26|141|-80.70901|21|35.17335|TRAIL MIXES AND BLENDS|0.0|1|FISHER ENERGY TRAIL MIX|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00070690271684|NUTS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|8fa063ecd4b4369373ff83299ba9f67a1ca70da1|1.99|2014-12-21 16:33:00|1.4094857484078087|2|7069027166|174|0.6138907664563474|0|26|141|-80.70901|21|35.17335|TRAIL MIXES AND BLENDS|0.0|1|FISHER ENERGY TRAIL MIX|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00070690271684|NUTS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|5b934caa37c9dd56af29dd56372a44b12e675a21|1.2|2015-02-22 19:57:00|1.4094857484078087|2|7047000641|174|0.6138907664563474|0|26|688|-80.70901|61|35.17335|LIGHT|0.2|3|YOPLAIT LIGHT BLUEBERRY|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00070470006529|YOGURT|DAIRY|-80.70901|1.4086379605250285|174|2
35.17335|1c882202d0294a4992986bac8aba8dc90b199ff8|1.99|2014-09-30 19:14:00|80.709059419360486|2|7069027166|174|35.18473217051357|0|31|141|-80.654118|21|35.123768|TRAIL MIXES AND BLENDS|0.99|1|FISHER ENERGY TRAIL MIX|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|35.187384292804154|00070690271684|NUTS|G1 GROCERY|-80.70901|80.709013723936394|473|1
35.17335|5eeba87d552e27229e56900c1cbd863cb29852f1|3.59|2014-12-22 20:07:00|1.4094857484078087|2|4150022020|174|0.6138907664563474|0|26|164|-80.70901|39|35.17335|VEGETABLES-SPECIALTY|1.8|1|FRENCHS FRIED ONION 6 OZ|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00041500220208|VEGETABLES-CAN/JAR|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|1c1446d2a25418e3a5870fb03f3bfcc332301aa8|4.99|2014-11-13 22:18:00|1.4094857484078087|2|3700039316|174|0.6138907664563474|0|26|726|-80.70901|73|35.17335|NFS-BODY WASHES|1.0|1|OLD SPC RED ZN SWAGGER BDYWASH|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00037000167709|PERSONAL SOAP/BATH ADDITIVES|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|5f93e985932d4ca51ed86ef261bc2537722f8c34|4.79|2014-10-15 21:11:00|1.4094857484078087|2|85641600001|174|0.6138907664563474|0|26|1433|-80.70901|9|35.17335|GRANOLA|1.79|1|BEAR NAKED GRN FIT TRIPLE BERY|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00856416000703|CEREAL|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|d35f97d709c0bd431b7e12fda872912c0afcd9fa|4.35|2015-03-03 19:08:00|1.4094857484078087|2|85641600001|174|0.6138907664563474|0|26|1433|-80.70901|9|35.17335|GRANOLA|0.0|1|BEAR NAKED GRN FIT TRIPLE BERY|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00856416000703|CEREAL|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|253c65dc13e772f1cd6acd92a4c0550358b2ab82|1.99|2015-01-13 21:42:00|1.4094857484078087|2|1111033407|174|0.6138907664563474|0|26|6654|-80.70901|1564|35.17335|HOME/OFFICE-GLUE|0.0|18|OFFICE WORKS SUPR GLUE GEL 2PK|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00011110334077|SCHOOL & OFFICE SUPPLY|GM|-80.70901|1.4086379605250285|174|1
35.17335|473fa321a01eb0f6dc66d3d94c861bc4308dc795|4.19|2014-10-13 18:50:00|1.4094857484078087|2|4812110208|174|0.6138907664563474|0|26|1037|-80.70901|164|35.17335|ENGLISH MUFFINS|2.1|7|THOMAS ENG MUFFN ORIG 6 PK PP|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00048121102081|BREAKFAST|COMMERCIAL BAKERY|-80.70901|1.4086379605250285|174|1
35.17335|6bb9acc574a46087d89df87120f8d8231cb2effd|2.49|2015-01-20 10:01:00|1.4094857484078087|2|8079380391|174|0.6138907664563474|0|26|97|-80.70901|8|35.17335|ENERGY DRINKS|0.0|23|NOS 16 OZ REG CAN|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00080793803910|CARBONATED BEVERAGES|BEVERAGE|-80.70901|1.4086379605250285|174|1
35.17335|0219e36a7810c90f7764689b1b5840a079bbc426|9.96|2014-09-18 19:29:00|80.709059419360486|2|8079380391|174|35.184732169659284|0|31|97|-80.739|8|35.141204|ENERGY DRINKS|4.96|23|NOS 16 OZ REG CAN|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|35.187384292804154|00080793803910|CARBONATED BEVERAGES|BEVERAGE|-80.70901|80.70901655571835|171|4
35.17335|356b2c51bc1d36e722ea4cd0122b38a297e819f3|4.98|2014-12-13 10:37:00|1.4094857484078087|2|8079380391|174|0.6138907664563474|0|26|97|-80.70901|8|35.17335|ENERGY DRINKS|2.48|23|NOS 16 OZ REG CAN|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00080793803910|CARBONATED BEVERAGES|BEVERAGE|-80.70901|1.4086379605250285|174|2
35.17335|4c7d6d9a72c66aae7702d56a8c90dfa7607c4947|2.49|2014-11-15 22:23:00|1.4094857484078087|2|8079380391|174|0.6138907664563474|0|26|97|-80.70901|8|35.17335|ENERGY DRINKS|1.24|23|NOS 16 OZ REG CAN|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00080793803910|CARBONATED BEVERAGES|BEVERAGE|-80.70901|1.4086379605250285|174|1
35.17335|8198c15619ea95b97fd541f7f7ad0acde19f03cc|7.470000000000001|2014-11-14 16:01:00|1.4094857484078087|2|8079380391|174|0.6138907664563474|0|26|97|-80.70901|8|35.17335|ENERGY DRINKS|3.7199999999999998|23|NOS 16 OZ REG CAN|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00080793803910|CARBONATED BEVERAGES|BEVERAGE|-80.70901|1.4086379605250285|174|3
35.17335|956b5584ee91b4da72fcf36b1ac36441daac068b|0.97|2015-01-09 21:32:00|1.4094857484078087|2|7203697849|174|0.6138907664563474|0|26|1251|-80.70901|12|35.17335|WHOLESOME COOKIES|0.0|1|HT FIG BARS|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00072036978493|COOKIES|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|2a94ca93986a7129a33eabb5ec986ffae6296a28|1.69|2015-01-29 10:23:00|1.4094857484078087|2|1200000129|174|0.6138907664563474|0|26|55|-80.70901|8|35.17335|REGULAR|0.0|23|CB PEPSI COLA 20 0Z|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00012000001291|CARBONATED BEVERAGES|BEVERAGE|-80.70901|1.4086379605250285|174|1
35.17335|d105ff38496fa7970865801bc62d796619e62267|4.99|2014-12-02 13:26:00|1.4094857484078087|2|3700047984|174|0.6138907664563474|0|26|726|-80.70901|73|35.17335|NFS-BODY WASHES|1.0|1|GILL DRY SKIN HYDRATOR&BDYWSH|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00037000479840|PERSONAL SOAP/BATH ADDITIVES|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|a65222634fecdc611243d11480228f8529f1193f|4.19|2014-10-03 18:36:00|1.4094857484078087|2|81793900734|174|0.6138907664563474|0|26|725|-80.70901|66|35.17335|NFS-DISHWASHING LIQUID|2.22|1|METHOD DISH SOAP CLEMENTINE|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00817939007358|DETERGENTS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|e8a6c0b42cc07ce42cb0894291981eb4dcb87de6|2.69|2014-12-03 20:28:00|1.4094857484078087|2|7203688023|174|0.6138907664563474|0|26|555|-80.70901|64|35.17335|PACKAGED SALADS|0.0|4|HT CURLY SPINACH,PKG|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00072036880239|FRESH PRODUCE|PRODUCE|-80.70901|1.4086379605250285|174|1
35.17335|c53578457ae8a46165115a138ce6a4d86906d3a2|5.78|2015-01-01 19:27:00|1.4094857484078087|2|7203663102|174|0.6138907664563474|0|26|339|-80.70901|57|35.17335|EGGNOGS/DRINKS|0.78|3|I/O HARRIS TEETER LT EGG NOG|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00072036631039|MILK|DAIRY|-80.70901|1.4086379605250285|174|2
35.17335|cf1a723b025863931ec6034bbc5acbf25e8a8543|7.38|2014-12-05 20:33:00|80.709059419360486|2|73291322733|174|35.18473217051357|0|31|725|-80.654118|66|35.123768|NFS-DISHWASHING LIQUID|2.38|1|7TH GEN DISH LIQ ULTRA POWER|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|35.187384292804154|00732913229284|DETERGENTS|G1 GROCERY|-80.70901|80.709013723936394|473|2
35.17335|d15342b9706a85e6a8aec067c3d58588aa692046|5.99|2014-09-20 16:24:00|80.709059419360486|2|7203695643|174|35.184732164768299|0|31|1663|-80.64817|381|35.04711|CREME CAKE|0.0|14|44 OZ CHOC CREME CAKE|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|35.187384292804154|00072036956644|CAKES|BAKERY|-80.70901|80.709024478830585|129|1
35.17335|f10ffc9b4129740190bf0ca57d684062753ba3af|4.29|2015-03-04 18:18:00|1.4094857484078087|2|3000006119|174|0.6138907664563474|0|26|74|-80.70901|9|35.17335|RTE CEREAL ALL FAMILY|0.0|1|QUAKER CINNAMON LIFE|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00030000060834|CEREAL|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|1cad6f1d946bdd70e6a161f31e2c8220964e5d7b|3.35|2015-02-01 20:01:00|1.4094857484078087|2|2840005597|174|0.6138907664563474|0|26|199|-80.70901|31|35.17335|DIPS & SALSAS|1.67|1|TOSTITOS HOT SALSA|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00028400055994|SNACKS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|7bbdee65ea4707067d75d8a2b9756259fc189cb9|0.33|2015-01-30 12:04:00|80.709059419360486|2||174|35.18473217040431|0|31|502|-80.826724|64|35.195689|FRESH BANANAS|0.0|4|BANANAS, YELLOW|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|35.187384292804154|00204011000008|FRESH PRODUCE|PRODUCE|-80.70901|80.7090141941556|412|1
35.17335|815846c115c2d215230dd12dc45ab4be09fc8416|2.29|2014-10-18 15:24:00|80.709059419360486|2|1900008501|174|35.18473217040431|0|31|50|-80.826724|7|35.195689|PEG CANDY|0.29|1|LIFESAVERS GUMMIES COOLERS PEG|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|35.187384292804154|00022000122643|CANDY|G1 GROCERY|-80.70901|80.7090141941556|412|1
35.17335|955e5827fbff9d9f5636d9f80a28d729031f4dcb|6.99|2014-12-07 18:29:00|1.4094857484078087|2|3700013885|174|0.6138907664563474|0|26|389|-80.70901|66|35.17335|NFS-LAUNDRY DETERGENTS|0.5|1|TIDE HE ORIGINAL W/BLEACH|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00037000875482|DETERGENTS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|33cad61fda3c3829eacf114e23850d6c41322a32|3.0|2014-11-18 19:39:00|1.4094857484078087|2|7047000100|174|0.6138907664563474|0|26|687|-80.70901|61|35.17335|BLENDED|0.5|3|YOPLAIT ORG MIXED BERRY|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00070470003108|YOGURT|DAIRY|-80.70901|1.4086379605250285|174|5
35.17335|1e63675f8b0c379e6900849728763b1938d22df4|8.97|2014-11-01 17:42:00|80.709059419360486|2|3993805735|174|35.184732164768299|0|31|7278|-80.64817|1600|35.04711|HALLOWEEN PARTY GOODS/DECOR|6.720000000000001|18|SPIDER ZIPPER BAG|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|35.187384292804154|00039938057374|SEASONAL MERCHANDISE|GM|-80.70901|80.709024478830585|129|3
35.17335|c9692f36ae9808cd3c11ba20a3a0410233ec010c|3.89|2014-12-26 20:52:00|1.4094857484078087|2|4127101787|174|0.6138907664563474|0|26|341|-80.70901|57|35.17335|CREAMERS|0.42|3|DUNKIN DONUTS EXTRA EXTRA 32OZ|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00041271017885|MILK|DAIRY|-80.70901|1.4086379605250285|174|1
35.17335|9e90206c16fd6b38dcabc67b48d2113d5858e46d|1.37|2014-12-21 22:27:00|80.709059419360486|2|7203627034|174|35.184732169659284|0|31|155|-80.739|24|35.141204|NFS-DOG TREATS|0.0|1|HT YOURPET WVY BACON CHEESE|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|35.187384292804154|00072036270337|PET FOOD/SUPPLIES|G1 GROCERY|-80.70901|80.70901655571835|171|1
35.17335|070855ad7d4e541078cbb2d0c0fcd99cc597c3c7|4.99|2014-10-14 21:20:00|1.4094857484078087|2|82744400099|174|0.6138907664563474|0|26|4954|-80.70901|1245|35.17335|EYE-SOFT LENS SALINES|1.0|17|REVITALENS MP SOL TRAVEL|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00827444000997|EYE & EAR CARE|HBC|-80.70901|1.4086379605250285|174|1
35.17335|252b891fc445ef936de97d6bae706d951d22e0df|0.76|2014-10-11 20:19:00|1.4094857484078087|2||174|0.6138907664563474|0|26|502|-80.70901|64|35.17335|FRESH BANANAS|0.0|4|BANANAS, YELLOW|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00204011000008|FRESH PRODUCE|PRODUCE|-80.70901|1.4086379605250285|174|1
35.17335|fcd6adbf83fe3e1e429592df4046873122c6b656|0.46|2014-11-15 14:04:00|1.4094857484078087|2||174|0.6138907664563474|0|26|502|-80.70901|64|35.17335|FRESH BANANAS|0.0|4|BANANAS, YELLOW|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00204011000008|FRESH PRODUCE|PRODUCE|-80.70901|1.4086379605250285|174|1
35.17335|6a907a37576a0189d1916714488f29646a32cef2|0.72|2014-12-05 15:05:00|1.4094857484078087|2||174|0.6138907664563474|0|26|502|-80.70901|64|35.17335|FRESH BANANAS|0.0|4|BANANAS, YELLOW|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00204011000008|FRESH PRODUCE|PRODUCE|-80.70901|1.4086379605250285|174|1
35.17335|a17fd21dfd0d6d849bfd7070951dce11be2f3d23|0.53|2015-02-24 21:05:00|1.4094857484078087|2||174|0.6138907664563474|0|26|502|-80.70901|64|35.17335|FRESH BANANAS|0.0|4|BANANAS, YELLOW|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00204011000008|FRESH PRODUCE|PRODUCE|-80.70901|1.4086379605250285|174|1
35.17335|e4e2318c75d5265855fe8281d31014718031f77e|0.73|2015-02-22 18:48:00|1.4094857484078087|2||174|0.6138907664563474|0|26|502|-80.70901|64|35.17335|FRESH BANANAS|0.0|4|BANANAS, YELLOW|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00204011000008|FRESH PRODUCE|PRODUCE|-80.70901|1.4086379605250285|174|1
35.17335|e0d62bbb4fe22e8c3a634b685f6e5bdfaa347b77|2.49|2014-11-29 10:26:00|1.4094857484078087|2|1200001643|174|0.6138907664563474|0|26|97|-80.70901|8|35.17335|ENERGY DRINKS|1.0|23|MTN DEW AMP TALL  BOY|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00012000016431|CARBONATED BEVERAGES|BEVERAGE|-80.70901|1.4086379605250285|174|1
35.17335|d41b7b4b76301aa5e959505e9a7a907e6e60ab7f|2.35|2014-12-10 20:25:00|1.4094857484078087|2|1480000010|174|0.6138907664563474|0|26|104|-80.70901|16|35.17335|APPLESAUCE-CUPS|0.0|1|MOTTS 6PK APLSC CINNAMON|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00014800000238|FRUIT-CAN/JAR|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|421e161a884e0e8aba513defa723d52cd4762436|1.59|2015-03-03 20:55:00|1.4094857484078087|2|4650073332|174|0.6138907664563474|0|26|393|-80.70901|68|35.17335|NFS-AIR FRESHENERS|0.59|1|GLADE AEROSOL APPLE CINNAMON|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00046500733437|FRESHENERS/DEODORIZERS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|5eaa822d169499e3148be8d2ec78167b452cdc3b|1.59|2015-02-08 13:20:00|1.4094857484078087|2|4650073332|174|0.6138907664563474|0|26|393|-80.70901|68|35.17335|NFS-AIR FRESHENERS|0.59|1|GLADE AEROSOL APPLE CINNAMON|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00046500733437|FRESHENERS/DEODORIZERS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|d12c23a88a216599bf7e6135898c153b0647ca03|3.39|2014-10-17 15:11:00|1.4094857484078087|2|8705212799|174|0.6138907664563474|0|26|400|-80.70901|69|35.17335|NFS-LIQUID CLEANERS|0.89|1|CITRUS MAGIC NTRL ALL PURP CLN|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00087052127992|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|84b67c25e247234f90f8dc7af7fd350bd9abc58b|3.99|2015-02-10 09:09:00|80.709059419360486|2|4400002854|174|35.18473217091757|0|31|1248|-80.810056|12|35.219587|SANDWICH COOKIES|0.49|1|OREO|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|35.187384292804154|00044000032029|COOKIES|G1 GROCERY|-80.70901|80.709010318724438|401|1
35.17335|2f37851d545f4c9a65aadd2e79b435c4a80a6ecc|2.99|2015-03-09 21:11:00|1.4094857484078087|2|7433610102|174|0.6138907664563474|0|26|342|-80.70901|57|35.17335|FRESH MILK|0.0|3|HIGHLAND CREST SKIM MILK|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00074336101083|MILK|DAIRY|-80.70901|1.4086379605250285|174|1
35.17335|ef836065e49d938e97dc5c1e82acec4a683c7116|7.1|2014-11-29 17:08:00|1.4094857484078087|2|7433610102|174|0.6138907664563474|0|26|342|-80.70901|57|35.17335|FRESH MILK|2.16|3|HIGHLAND CREST SKIM MILK|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00074336101083|MILK|DAIRY|-80.70901|1.4086379605250285|174|2
35.17335|964b98cb203a1a6ab62f13693a4375d6fe246e19|3.15|2014-12-08 17:46:00|1.4094857484078087|2|7225003706|174|0.6138907664563474|0|26|1026|-80.70901|162|35.17335|WHEAT|0.66|7|NATOWN HONEYWHEAT BRD|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00072250037068|SLICED BREAD|COMMERCIAL BAKERY|-80.70901|1.4086379605250285|174|1
35.17335|68e51b0628a76908f4d610702a4eb88544b15458|3.19|2014-09-27 13:50:00|1.4094857484078087|2|3680018458|174|0.6138907664563474|0|26|4010|-80.70901|1080|35.17335|DENTURE CLEANER PRODUCT|0.0|17|TC MINT DENTURE TABS 18458|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00036800184589|ORAL HYGIENE|HBC|-80.70901|1.4086379605250285|174|1
35.17335|c64ac56a0ec646361a088d9a83d18a0535a52e81|3.99|2014-10-02 20:30:00|1.4094857484078087|2|74447391224|174|0.6138907664563474|0|26|1265|-80.70901|57|35.17335|ALMOND MILK|1.99|3|SO DELICIOUS VAN ALMOND MILK|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00744473912247|MILK|DAIRY|-80.70901|1.4086379605250285|174|1
35.17335|1387a1ca47e7eb6a24f0e70779d3ceb2d14de361|5.99|2014-11-25 19:02:00|1.4094857484078087|2|85822200126|174|0.6138907664563474|0|26|7209|-80.70901|1600|35.17335|BACK TO SCHOOL|0.0|18|I/OIPHONE 5 COMPATIBLE CABLE|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00858222001264|SEASONAL MERCHANDISE|GM|-80.70901|1.4086379605250285|174|1
35.17335|383fc536d72498a73286fdc9b5bbe72dcf17dfa0|5.99|2014-11-09 18:23:00|1.4094857484078087|2|85822200126|174|0.6138907664563474|0|26|7209|-80.70901|1600|35.17335|BACK TO SCHOOL|0.0|18|I/OIPHONE 5 COMPATIBLE CABLE|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00858222001264|SEASONAL MERCHANDISE|GM|-80.70901|1.4086379605250285|174|1
35.17335|89ad1a3c4ac691ac9cb9decaa9904539f771c3d5|2.99|2014-12-02 21:28:00|1.4094857484078087|2|2529360050|174|0.6138907664563474|0|26|339|-80.70901|57|35.17335|EGGNOGS/DRINKS|0.3|3|I/O SILK NOG|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00025293600508|MILK|DAIRY|-80.70901|1.4086379605250285|174|1
35.17335|074b9a8d32d2147e26f599be8fa3c81268801372|2.99|2014-12-20 20:04:00|1.4094857484078087|2|2529360050|174|0.6138907664563474|0|26|339|-80.70901|57|35.17335|EGGNOGS/DRINKS|0.3|3|I/O SILK NOG|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00025293600508|MILK|DAIRY|-80.70901|1.4086379605250285|174|1
35.17335|c10bedf4d10470b2b9e5c8eb7d3249603a517d1e|2.99|2014-12-18 21:52:00|1.4094857484078087|2|2529360050|174|0.6138907664563474|0|26|339|-80.70901|57|35.17335|EGGNOGS/DRINKS|0.3|3|I/O SILK NOG|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00025293600508|MILK|DAIRY|-80.70901|1.4086379605250285|174|1
35.17335|336d6c5ba2bb0641c403b57c3792e951d25e7fec|2.99|2014-11-23 19:27:00|1.4094857484078087|2|2529360050|174|0.6138907664563474|0|26|339|-80.70901|57|35.17335|EGGNOGS/DRINKS|0.3|3|I/O SILK NOG|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00025293600508|MILK|DAIRY|-80.70901|1.4086379605250285|174|1
35.17335|3bb4e1726e4c1fbec85d8476c216bb564f328ae8|5.98|2014-11-25 21:48:00|1.4094857484078087|2|2529360050|174|0.6138907664563474|0|26|339|-80.70901|57|35.17335|EGGNOGS/DRINKS|0.6|3|I/O SILK NOG|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00025293600508|MILK|DAIRY|-80.70901|1.4086379605250285|174|2
35.17335|8ca787b66523393ba79ea1fa117738bd97dd9dfa|2.99|2014-10-31 22:47:00|1.4094857484078087|2|2529360050|174|0.6138907664563474|0|26|339|-80.70901|57|35.17335|EGGNOGS/DRINKS|0.3|3|I/O SILK NOG|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00025293600508|MILK|DAIRY|-80.70901|1.4086379605250285|174|1
35.17335|60def405a3c4dc5e19a739b6bce95f4091dc5c7d|7.99|2015-01-05 22:04:00|1.4094857484078087|2|8079380924|174|0.6138907664563474|0|26|97|-80.70901|8|35.17335|ENERGY DRINKS|3.0|23|NOS 12 OZ 6PK CANS|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00080793809240|CARBONATED BEVERAGES|BEVERAGE|-80.70901|1.4086379605250285|174|1
35.17335|6d582047bfa9049a1530e66eb7ff6ea76e506b35|7.99|2015-01-26 08:59:00|1.4094857484078087|2|8079380924|174|0.6138907664563474|0|26|97|-80.70901|8|35.17335|ENERGY DRINKS|3.0|23|NOS 12 OZ 6PK CANS|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00080793809240|CARBONATED BEVERAGES|BEVERAGE|-80.70901|1.4086379605250285|174|1
35.17335|cfa03ac7e6d9106a16ece47cf09e44a9d2c6c278|4.99|2014-12-20 14:54:00|80.709059419360486|2|71575620002|174|35.18473217043951|0|31|504|-80.844274|64|35.204336|FRESH BERRIES|0.0|4|STRAWBERRIES 1LB CLAM|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|35.187384292804154|00812049005102|FRESH PRODUCE|PRODUCE|-80.70901|80.709014048636988|61|1
35.17335|b592ab6fb22b2b7a283e4e5476ec07c923ae100a|5.97|2015-01-07 21:11:00|1.4094857484078087|2|7069027166|174|0.6138907664563474|0|26|141|-80.70901|21|35.17335|TRAIL MIXES AND BLENDS|2.9699999999999998|1|FISHER HUNGER FIGHTR TRAIL MIX|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00070690271837|NUTS|G1 GROCERY|-80.70901|1.4086379605250285|174|3
35.17335|4ec2042e7e19e54def8eee7219c9542871e38bb6|1.99|2014-12-14 18:27:00|1.4094857484078087|2|7069027166|174|0.6138907664563474|0|26|141|-80.70901|21|35.17335|TRAIL MIXES AND BLENDS|0.0|1|FISHER HUNGER FIGHTR TRAIL MIX|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00070690271837|NUTS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|9c04968ba272088521353271e7912cdd11d77841|1.99|2014-11-22 18:18:00|1.4094857484078087|2|7069027166|174|0.6138907664563474|0|26|141|-80.70901|21|35.17335|TRAIL MIXES AND BLENDS|0.49|1|FISHER HUNGER FIGHTR TRAIL MIX|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00070690271837|NUTS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|5b535e04b9169a7e09761b36a0c974bd75c86580|1.99|2014-10-10 19:20:00|1.4094857484078087|2|7069027166|174|0.6138907664563474|0|26|141|-80.70901|21|35.17335|TRAIL MIXES AND BLENDS|0.0|1|FISHER HUNGER FIGHTR TRAIL MIX|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00070690271837|NUTS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|0bc64e498fb11bbe1897496399d415039f063032|3.98|2014-10-07 19:49:00|1.4094857484078087|2|7069027166|174|0.6138907664563474|0|26|141|-80.70901|21|35.17335|TRAIL MIXES AND BLENDS|1.98|1|FISHER HUNGER FIGHTR TRAIL MIX|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00070690271837|NUTS|G1 GROCERY|-80.70901|1.4086379605250285|174|2
35.17335|f6aae3f14fb52155682a39b0ad7080022d015309|1.99|2014-12-03 17:28:00|1.4094857484078087|2|7069027166|174|0.6138907664563474|0|26|141|-80.70901|21|35.17335|TRAIL MIXES AND BLENDS|0.0|1|FISHER HUNGER FIGHTR TRAIL MIX|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00070690271837|NUTS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|65e2a96443fbba80573ba70706b8a9ab3bdbd647|3.15|2014-12-04 13:13:00|1.4094857484078087|2|3000001190|174|0.6138907664563474|0|26|60|-80.70901|9|35.17335|HOT CEREAL|0.65|1|QUAKER OATML CINN SPICE|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00030000312087|CEREAL|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|5314c43328f4e2bfcc4be076d8f0034958a3b83a|6.98|2014-10-19 21:36:00|1.4094857484078087|2|3000001190|174|0.6138907664563474|0|26|60|-80.70901|9|35.17335|HOT CEREAL|0.99|1|QUAKER OATML CINN SPICE|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00030000312087|CEREAL|G1 GROCERY|-80.70901|1.4086379605250285|174|2
35.17335|84dfb5a790387936d8076b9389f8eab46178973a|3.15|2014-11-01 22:12:00|1.4094857484078087|2|3000001190|174|0.6138907664563474|0|26|60|-80.70901|9|35.17335|HOT CEREAL|0.36|1|QUAKER OATML CINN SPICE|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00030000312087|CEREAL|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|a36506b8ce1802ae481c3cc732691a2ccd12a37b|4.29|2014-09-11 20:39:00|1.4094857484078087|2|2840006399|174|0.6138907664563474|0|26|204|-80.70901|31|35.17335|TORTILLA CHIPS|1.79|1|TOSTITOS SCOOPS 10 OZ|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00028400064088|SNACKS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|9038d7a7456724d7ca37631f93ef0f3418540362|3.95|2014-12-14 18:24:00|1.4094857484078087|2|7203663995|174|0.6138907664563474|0|26|342|-80.70901|57|35.17335|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00072036631282|MILK|DAIRY|-80.70901|1.4086379605250285|174|1
35.17335|14c6021ae261eaad48b91c6925393466ae759d5b|6.98|2015-02-08 13:18:00|1.4094857484078087|2|7203663995|174|0.6138907664563474|0|26|342|-80.70901|57|35.17335|FRESH MILK|1.72|3|HARRIS TEETER FF SKIM MILK|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00072036631282|MILK|DAIRY|-80.70901|1.4086379605250285|174|2
35.17335|d6a192248cae2fa81ecb3ba9984d880dcb1bd0c1|2.39|2015-02-14 15:56:00|1.4094857484078087|2|7084781116|174|0.6138907664563474|0|26|97|-80.70901|8|35.17335|ENERGY DRINKS|0.0|23|MONSTER ENERGY CAN|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|0.61471665291522548|00070847811169|CARBONATED BEVERAGES|BEVERAGE|-80.70901|1.4086379605250285|174|1
35.17335|98d3d72568d9c553537e7432eb4721d5f04f58fa|2.99|2014-12-16 16:50:00|80.709059419360486|2|20443000000|174|35.18473217043951|0|31|510|-80.844274|64|35.204336|FRESH PINEAPPLE|0.0|4|GOLD PINEAPPLES|20ae36c4b3d87834aa1107b125dfc9f10e128f20|0.7864805236518413|35.187384292804154|00643126072003|FRESH PRODUCE|PRODUCE|-80.70901|80.709014048636988|61|1
35.297134|b6fa85c9c876303b455876a26faae34d80b5b986|3.79|2015-01-07 13:09:00|1.4094857484078087|4|2100062503|258|0.6160512048176361|0|26|318|-80.737839|52|35.297134|SHREDDED/GRATED CHEESE|1.29|3|KRAFT 2% SHARP SHRED|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00021000024605|CHEESE|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|f2e20fd132631534c4d834935e24213d04e3b4f6|1.27|2014-09-25 10:48:00|1.4094857484078087|4|7203628032|258|0.6160512048176361|0|26|163|-80.737839|25|35.297134|RELISHES|0.0|1|HT RELISH SWEET 16|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00072036280329|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.737839|1.409141121495086|258|1
35.297134|0aba3658f0b2decdeddbf94c0d77ac3a0a0909ef|2.79|2014-12-11 10:41:00|1.4094857484078087|4|7365111706|258|0.6160512048176361|0|26|160|-80.737839|25|35.297134|OLIVES|1.4|1|MARIO OLIVE MANZ 5.75|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00073651117069|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.737839|1.409141121495086|258|1
35.297134|ae9cd4a49f33fb5dffb3ac0287ccd6530bc8f0ee|2.75|2014-11-13 11:07:00|1.4094857484078087|4|930018709|258|0.6160512048176361|0|26|162|-80.737839|25|35.297134|PICKLES|1.38|1|MT OLV CHIPS BREAD & BUTR 24FP|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00009300000772|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.737839|1.409141121495086|258|1
35.297134|5f03587091481af5d7ab2d1e651f6c1614d960b3|7.78|2014-12-06 11:49:00|1.4094857484078087|4|5450019352|258|0.6160512048176361|0|26|359|-80.737839|101|35.297134|MEAT WIENERS|1.94|19|BALL PARK FRANKS|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00054500193526|WIENERS|CASE READY MEATS|-80.737839|1.409141121495086|258|2
35.297134|312f6dbaa6d1f032435cb2391169de015c6fe876|6.5|2014-10-31 11:47:00|1.4094857484078087|4|5150025362|258|0.6160512048176361|0|26|195|-80.737839|30|35.297134|SALAD & COOKING OIL|0.92|1|CRISCO CANOLA OIL|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00051500251515|SHORTENING/OIL|G1 GROCERY|-80.737839|1.409141121495086|258|2
35.297134|2ed07c6f9d7d406c4e5f5ae4bce1a2019b029d70|1.57|2014-12-16 10:31:00|80.737901233649083|4|7203601075|258|35.348004019597305|0|46|1267|-80.70901|53|35.17335|DIPS AND SPREADS|0.0|3|HT FRENCH ONION DIP 16 OZ|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|35.349871187060224|00072036010759|CULTURES|DAIRY|-80.737839|80.73791116456448|174|1
35.297134|a039e21e8ede386b476b0e0988c3acd4390f75fb|1.29|2015-03-06 11:26:00|1.4094857484078087|4|4920005675|258|0.6160512048176361|0|26|224|-80.737839|35|35.297134|SUGAR-BROWN|0.0|1|DOMINO LT BRWN SUGAR-BOX|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00049200056752|SUGAR/SUBSTITUTES|G1 GROCERY|-80.737839|1.409141121495086|258|1
35.297134|43821b0ccf9e79ad6ad241f0905f80f631d15e61|7.89|2015-01-29 10:45:00|1.4094857484078087|4|2770067902|258|0.6160512048176361|0|26|270|-80.737839|307|35.297134|DESSERTS FROZEN|6.9|5|I/O M SMITHS FLKY CRUST SW POT|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00027700679060|DESSERTS FROZEN|FROZEN|-80.737839|1.409141121495086|258|1
35.297134|9ace665f375a0dcf92e7b1f88f8d6bfcc3b6a32c|4.99|2014-12-20 11:15:00|1.4094857484078087|4|7203688058|258|0.6160512048176361|0|26|562|-80.737839|64|35.297134|FRESH CUT FRUIT|1.0|4|HT CORED GOLDEN PINEAPPLE|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00072036880581|FRESH PRODUCE|PRODUCE|-80.737839|1.409141121495086|258|1
35.297134|e1c42b59dbdd73b95f4a147a886d335378985379|19.98|2015-02-12 12:08:00|1.4094857484078087|4|7203661016|258|0.6160512048176361|0|26|297|-80.737839|49|35.297134|GROUND BEEF|14.0|2|GROUND CHUCK 80% LEAN 2 LB|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00072036610164|BEEF|MEAT|-80.737839|1.409141121495086|258|2
35.297134|bee9ad95abe18cc66bad22e3983ca0a396b8fcf4|3.63|2015-03-05 10:32:00|1.4094857484078087|4||258|0.6160512048176361|0|26|503|-80.737839|64|35.297134|FRESH GRAPES|2.08|4|RED GRAPES,SEEDLESS 12/16|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00204023000003|FRESH PRODUCE|PRODUCE|-80.737839|1.409141121495086|258|1
35.297134|2ededcdf22c1dc4df029071580caa52596ace8ca|3.35|2014-09-18 11:15:00|1.4094857484078087|4|7203656080|258|0.6160512048176361|0|26|318|-80.737839|52|35.297134|SHREDDED/GRATED CHEESE|1.35|3|HT FANCY SHRED MILD CHED CHES|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00072036560810|CHEESE|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|e7b3d22610ba6b2c33dac37e0b407fb2ce0807ad|3.35|2014-10-23 11:30:00|1.4094857484078087|4|7203656080|258|0.6160512048176361|0|26|318|-80.737839|52|35.297134|SHREDDED/GRATED CHEESE|1.68|3|HT FANCY SHRED SHARP CHED CHE|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00072036550262|CHEESE|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|0dfd8a37a69f929dccc3a343a29dee7364c5fc48|3.99|2015-01-22 12:14:00|1.4094857484078087|4|1090000015|258|0.6160512048176361|0|26|440|-80.737839|76|35.297134|NFS-ALUMINUM FOIL|0.0|1|REYNOLDS FOIL 75 FT|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00010900000154|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.737839|1.409141121495086|258|1
35.297134|f578f84d9ae6499f11851e388a6cd443a4461076|3.99|2014-11-25 11:07:00|1.4094857484078087|4|7203688049|258|0.6160512048176361|0|26|562|-80.737839|64|35.297134|FRESH CUT FRUIT|0.0|4|HT MIXED FRUIT CHUNKS 16OZ|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00072036880499|FRESH PRODUCE|PRODUCE|-80.737839|1.409141121495086|258|1
35.297134|62cecacc319fcac72ad18af1edd0fd440b8d99f6|2.45|2014-10-16 10:54:00|1.4094857484078087|4|7203663217|258|0.6160512048176361|0|26|330|-80.737839|55|35.297134|EGGS|0.45|3|HT GRADE A LARGE EGGS 18 CT|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00072036632173|EGGS FRESH|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|f79fbd5b46b516009430d8b0e1b4dc6aa79fde08|3.99|2014-10-13 10:40:00|1.4094857484078087|4|7203663995|258|0.6160512048176361|0|26|342|-80.737839|57|35.297134|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00072036631282|MILK|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|eb6fc1cc3cc1f161b5e02c35061d0a4ba4e654bb|14.98|2014-11-20 10:56:00|1.4094857484078087|4|7203661029|258|0.6160512048176361|0|26|671|-80.737839|147|35.297134|OYSTERS|2.0|12|FISHERMAN'S MKT STND OYSTERS|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00072036610294|MOLLUSK|SEAFOOD|-80.737839|1.409141121495086|258|2
35.297134|9fc9d8073e6ce28fb3bf2c51c3417ac43b6aa439|2.69|2014-10-09 10:01:00|80.737901233649083|4|7203663996|258|35.348004020931938|0|46|342|-80.810056|57|35.219587|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|35.349871187060224|00072036631299|MILK|DAIRY|-80.737839|80.737909737224996|401|1
35.297134|26697f05f77448558e68fd04650c0660755c7ff2|2.59|2014-12-06 11:57:00|1.4094857484078087|4|7203663996|258|0.6160512048176361|0|26|342|-80.737839|57|35.297134|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00072036631299|MILK|DAIRY|-80.737839|1.409141121495086|258|1
35.297134|6b3ba0092f7eb73eb4fbd7a4e7c4261a66c8247f|4.79|2015-01-10 10:26:00|1.4094857484078087|4|75703751313|258|0.6160512048176361|0|26|420|-80.737839|71|35.297134|NFS-SOIL/SPOT/STAIN REMO|0.0|1|OXI CLEAN STAIN REMOVER 28LOAD|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00757037513132|LAUNDRY SUPPLIES|G1 GROCERY|-80.737839|1.409141121495086|258|1
35.297134|aedea3e009b97eea41041154683ca82da8e02067|1.47|2015-02-09 11:45:00|1.4094857484078087|4|7203625014|258|0.6160512048176361|0|26|145|-80.737839|22|35.297134|MILK-CANNED|0.0|1|HT SWEETENED CONDENSED MILK|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00072036250148|PACKAGED MILKS & MODIFIERS|G1 GROCERY|-80.737839|1.409141121495086|258|1
35.297134|bc14ad090bb6b29ad511a0a32426d8285d3aa5cf|4.99|2014-11-07 11:35:00|1.4094857484078087|4|2073511020|258|0.6160512048176361|0|26|252|-80.737839|45|35.297134|PREMIUM ICE CREAM|1.99|5|TURKEY HILL DUTCH CHOC IC|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00020735420959|ICE CREAM|FROZEN|-80.737839|1.409141121495086|258|1
35.297134|916ea2f67fbd0c8b4dc472d76eb5267b23b071f3|5.99|2014-10-25 11:01:00|80.737901233649083|4|7203688134|258|35.348004053647294|0|46|563|-80.780702|64|35.318911|FRESH VEGETABLE/FRUIT TRAYS|0.0|4|HT VEGETABLE TRAY, SMALL|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|35.349871187060224|00072036881342|FRESH PRODUCE|PRODUCE|-80.737839|80.737840969163074|167|1
35.297134|a5b18c64fd457faf21e3c012255853a2dd83dcf2|2.45|2014-11-21 11:13:00|1.4094857484078087|4|1450000253|258|0.6160512048176361|0|26|1273|-80.737839|50|35.297134|BAG VEG NON STEAM|1.23|5|BE BABY WHITE CORN|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00014500002907|VEGETABLES-FROZEN|FROZEN|-80.737839|1.409141121495086|258|1
35.297134|3ba7e1e3fa87a5dce87364e43593e485a80b49ed|4.9|2014-10-31 12:02:00|1.4094857484078087|4|1450000253|258|0.6160512048176361|0|26|1273|-80.737839|50|35.297134|BAG VEG NON STEAM|1.56|5|BE BABY WHITE CORN|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00014500002907|VEGETABLES-FROZEN|FROZEN|-80.737839|1.409141121495086|258|2
35.297134|74f3e45d1b89b25ea0c7cc9b96d9c62009befbbb|7.89|2015-01-29 10:53:00|1.4094857484078087|4|2770067902|258|0.6160512048176361|0|26|270|-80.737839|307|35.297134|DESSERTS FROZEN|6.9|5|I/O M SMITHS FLKY CRUST PMPKN|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00027700679077|DESSERTS FROZEN|FROZEN|-80.737839|1.409141121495086|258|1
35.297134|fd1d20622ce4b61d3818ce622076457e6ab4071a|3.5|2014-09-29 09:53:00|1.4094857484078087|4|2920000212|258|0.6160512048176361|0|26|149|-80.737839|23|35.297134|WHSE PASTA CORE|0.88|1|MUELLER POT SZ SPAGHETTI THIN|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00029200907957|PASTA|G1 GROCERY|-80.737839|1.409141121495086|258|2
35.297134|1a774edd324a3858d6244306884c764567c1a1ac|3.69|2014-10-13 10:47:00|1.4094857484078087|4|1620033700|258|0.6160512048176361|0|26|225|-80.737839|35|35.297134|SUGAR-GRANULATED|1.2|1|DIXIE CRYSTAL 4 LB GRAN SUGAR|22e72c8bf7973945acd6b3c89196c06cc4aa8886|3.514997861999427|0.61471665291522548|00016200337006|SUGAR/SUBSTITUTES|G1 GROCERY|-80.737839|1.409141121495086|258|1
35.297134|0ce205e15b9554560521819620cd273837cb8050|3.19|2014-09-28 09:00:00|80.728244613218536|4|4667501350|258|35.319865533884958|0|5|682|-80.764523|61|35.341927|KIDS|0.0|3|YOCRUNCH BAN/NILLA WAFER 4PK|23c8afa312d6f4fe8796310fc552c82b10a6a7a9|1.5706941898861861|35.296297200616316|00046675013297|YOGURT|DAIRY|-80.737839|80.737848592077654|220|1
35.297134|da85a8abd4d8ca51c6038db7d6d841cd545d4b07|3.89|2015-02-15 18:51:00|1.4094857484078087|4|7045900555|258|0.6160512048176361|0|26|1461|-80.737839|40|35.297134|FROZEN GARLIC TOAST AND BRD|0.0|5|NY SOFT GARLIC PULL APARTS|23c8afa312d6f4fe8796310fc552c82b10a6a7a9|1.5706941898861861|0.61471665291522548|00070459005277|FROZEN DOUGH|FROZEN|-80.737839|1.409141121495086|258|1
35.297134|63a1526f569f60b31eb2bffb46e1f322effa0172|4.29|2015-02-18 06:13:00|1.4094857484078087|4|1380010067|258|0.6160512048176361|0|26|1280|-80.737839|48|35.297134|MULTI SERVE MEALS|0.95|5|STOUFFER MEAT LOVERS LASAGNA|23c8afa312d6f4fe8796310fc552c82b10a6a7a9|1.5706941898861861|0.61471665291522548|00013800869807|FROZEN MEALS|FROZEN|-80.737839|1.409141121495086|258|1
35.297134|d6313016e7dbeb9f3b025402a643bbc42e0bc7fd|2.99|2015-03-06 13:52:00|80.728244613218536|4|81097900392|258|35.31986551305868|0|5|1246|-80.762919|34|35.442529|SPICE BLENDS|1.0|1|TRUE LIME GARLIC & CILANTRO|23c8afa312d6f4fe8796310fc552c82b10a6a7a9|1.5706941898861861|35.296297200616316|00810979003922|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.737839|80.737877907524648|471|1
35.297134|d6684b9353068fab5f8021268956077ed0459cbf|4.69|2014-10-07 06:09:00|1.4094857484078087|4|3736300612|258|0.6160512048176361|0|26|1279|-80.737839|48|35.297134|SINGLE SERVE FLAVOR|1.36|5|MICH ANGELO CHCKN PARMESAN|23c8afa312d6f4fe8796310fc552c82b10a6a7a9|1.5706941898861861|0.61471665291522548|00037363571243|FROZEN MEALS|FROZEN|-80.737839|1.409141121495086|258|1
35.297134|8ff633d8e08af3e373c4b3a257b7e84506b1374d|7.99|2014-10-18 06:45:00|80.728244613218536|4|1114110526|258|35.319865533884958|0|5|36|-80.764523|10|35.341927|PREMIUM GROUND|0.0|1|EIGHT OCLOCK DECAF GRND COFF|23c8afa312d6f4fe8796310fc552c82b10a6a7a9|1.5706941898861861|35.296297200616316|00011141105264|COFFEE|G1 GROCERY|-80.737839|80.737848592077654|220|1
35.297134|7f62e6b10cd86ab7aa0c32184a1415e312bf4973|5.19|2014-10-07 06:08:00|1.4094857484078087|4|89162700903|258|0.6160512048176361|0|26|1279|-80.737839|48|35.297134|SINGLE SERVE FLAVOR|3.19|5|EVOL ZITI BOLOGNESE|23c8afa312d6f4fe8796310fc552c82b10a6a7a9|1.5706941898861861|0.61471665291522548|00891627002962|FROZEN MEALS|FROZEN|-80.737839|1.409141121495086|258|1
35.03469|9362f1a0bb0afec4bcda96d4c6e9390c4f30fa6a|1.64|2014-12-09 14:39:00|1.4132775322775095|1||82|0.6114706929155321|0|58|502|-80.97058|64|35.03469|FRESH BANANAS|0.0|4|BANANAS, YELLOW|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00204011000008|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|124dd106615005451b72212cc382f7617f0bd4bd|1.59|2014-11-18 15:06:00|1.4132775322775095|1||82|0.6114706929155321|0|58|502|-80.97058|64|35.03469|FRESH BANANAS|0.0|4|BANANAS, YELLOW|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00204011000008|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|f3ed8eb7436a36f1015a571a348fc7c56a548e65|1.22|2015-01-19 18:10:00|80.970593795509558|1||82|35.050189210146748|0|4|502|-80.994596|64|35.061685|FRESH BANANAS|0.0|4|BANANAS, YELLOW|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|35.073829668338668|00204011000008|FRESH PRODUCE|PRODUCE|-80.97058|80.970583268867514|475|1
35.03469|414a530e992cad9445d4b571be0bf0bc43ebb2de|1.66|2014-12-03 15:46:00|1.4132775322775095|1||82|0.6114706929155321|0|58|502|-80.97058|64|35.03469|FRESH BANANAS|0.0|4|BANANAS, YELLOW|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00204011000008|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|832f2881bb1490757fe8baf29f9e48dc92c14074|1.57|2014-11-12 15:10:00|1.4132775322775095|1||82|0.6114706929155321|0|58|502|-80.97058|64|35.03469|FRESH BANANAS|0.0|4|BANANAS, YELLOW|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00204011000008|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|8e7bc5d911499b5d87b89a7a148c89abf52be143|1.39|2015-01-27 18:34:00|1.4132775322775095|1||82|0.6114706929155321|0|58|502|-80.97058|64|35.03469|FRESH BANANAS|0.0|4|BANANAS, YELLOW|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00204011000008|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|1243724e3ee2401e02e3d5fc47da78c7e653e976|1.16|2014-12-20 15:44:00|1.4132775322775095|1||82|0.6114706929155321|0|58|502|-80.97058|64|35.03469|FRESH BANANAS|0.0|4|BANANAS, YELLOW|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00204011000008|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|97db1edea3a552337fef4833b6573c96fbcc841c|1.56|2014-12-14 13:52:00|1.4132775322775095|1||82|0.6114706929155321|0|58|502|-80.97058|64|35.03469|FRESH BANANAS|0.0|4|BANANAS, YELLOW|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00204011000008|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|3f59a8288cc940ddbf3de6e1ac261e28d3678529|0.7|2014-10-26 11:11:00|1.4132775322775095|1||82|0.6114706929155321|0|58|502|-80.97058|64|35.03469|FRESH BANANAS|0.0|4|BANANAS, YELLOW|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00204011000008|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|ce37ac1846e937e2c6f9b4a7ec07555d6d1ef3cf|0.78|2014-10-29 15:00:00|1.4132775322775095|1||82|0.6114706929155321|1|58|502|-80.97058|64|35.03469|FRESH BANANAS|0.0|4|BANANAS, YELLOW|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00204011000008|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|a6e846524f66b7c632c96d480bf00f6017f0e7d3|0.91|2014-10-16 17:44:00|1.4132775322775095|1||82|0.6114706929155321|0|58|502|-80.97058|64|35.03469|FRESH BANANAS|0.0|4|BANANAS, YELLOW|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00204011000008|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|ccebb2fc6087d5dcf8f42f55393e062a3e7216d9|1.2|2014-09-21 20:02:00|1.4132775322775095|1||82|0.6114706929155321|0|58|502|-80.97058|64|35.03469|FRESH BANANAS|0.0|4|BANANAS, YELLOW|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00204011000008|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|90d74819f195e5d6420646d7ff393c19491b99dd|0.99|2015-01-30 17:25:00|1.4132775322775095|1||82|0.6114706929155321|0|58|502|-80.97058|64|35.03469|FRESH BANANAS|0.0|4|BANANAS, YELLOW|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00204011000008|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|a55f31262850de7466f61c970c9a5cc5dbc537e2|1.62|2014-11-07 12:41:00|1.4132775322775095|1||82|0.6114706929155321|0|58|502|-80.97058|64|35.03469|FRESH BANANAS|0.0|4|BANANAS, YELLOW|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00204011000008|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|651a6438e2a354f9171905ab4ca798f4a77e1b46|1.03|2015-01-12 14:48:00|1.4132775322775095|1||82|0.6114706929155321|0|58|502|-80.97058|64|35.03469|FRESH BANANAS|0.0|4|BANANAS, YELLOW|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00204011000008|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|bf584a4ba2170c6fc4c76d0e9a27cc1ea4b6058b|3.35|2014-09-22 17:54:00|80.970593795509558|1|7203656080|82|35.050189210146748|0|4|318|-80.994596|52|35.061685|SHREDDED/GRATED CHEESE|1.35|3|HT GOURMENT SHARP BLEND|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|35.073829668338668|00072036600783|CHEESE|DAIRY|-80.97058|80.970583268867514|475|1
35.03469|343aaccfddcb438ce7a79b99b05028b528b0a4be|9.99|2014-12-05 14:49:00|1.4132775322775095|1|8500001443|82|0.6114706929155321|0|58|9938|-80.97058|885|35.03469|NFS POP PINOT GRS/GRIGIO|0.0|13|CB-BAREFOOT PINOT GRIGIO 1.5L|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00085000014431|POPULAR (4-$7.99)|WINE|-80.97058|1.4132032182494703|82|1
35.03469|20e5c1429e4387cf0599c7696813d77d65294eaa|10.0|2014-10-13 16:16:00|1.4132775322775095|1|8143403123|82|0.6114706929155321|0|58|9934|-80.97058|885|35.03469|NFS POP CHARDONNAY|0.0|13|CB-REX GOLIATH CHARDONNAY|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00081434031235|POPULAR (4-$7.99)|WINE|-80.97058|1.4132032182494703|82|2
35.03469|a095b588af50a5977c7a6198e43522a52e2685d0|3.99|2015-02-15 12:36:00|1.4132775322775095|1|7835470843|82|0.6114706929155321|0|58|317|-80.97058|52|35.03469|CHUNK AND BAR CHEESE|0.4|3|CABOT EXTRA SHARP WHITE CHEDD|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00078354703182|CHEESE|DAIRY|-80.97058|1.4132032182494703|82|1
35.03469|016f0667fc4b7a93a9608ea7b2fc1756e292d4e5|3.99|2015-03-06 18:06:00|1.4132775322775095|1|7835470843|82|0.6114706929155321|0|58|317|-80.97058|52|35.03469|CHUNK AND BAR CHEESE|0.4|3|CABOT EXTRA SHARP WHITE CHEDD|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00078354703182|CHEESE|DAIRY|-80.97058|1.4132032182494703|82|1
35.03469|7b2e23848bdede0096a7b55ec66d1e1adc7f15cf|3.99|2014-11-02 17:04:00|1.4132775322775095|1|7835470843|82|0.6114706929155321|0|58|317|-80.97058|52|35.03469|CHUNK AND BAR CHEESE|1.49|3|CABOT EXTRA SHARP WHITE CHEDD|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00078354703182|CHEESE|DAIRY|-80.97058|1.4132032182494703|82|1
35.03469|73ab7c140de653f49ebcbfd7374ea9108cd1b354|3.99|2015-01-02 12:48:00|1.4132775322775095|1|7835470843|82|0.6114706929155321|0|58|317|-80.97058|52|35.03469|CHUNK AND BAR CHEESE|0.4|3|CABOT EXTRA SHARP WHITE CHEDD|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00078354703182|CHEESE|DAIRY|-80.97058|1.4132032182494703|82|1
35.03469|fdc88014ece51e10be300342b6c88806a65882fa|1.99|2014-10-12 11:02:00|1.4132775322775095|1|7203688096|82|0.6114706929155321|0|58|526|-80.97058|64|35.03469|FRESH MUSHROOMS|0.0|4|HT SLICED WHITE MUSHROOMS|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00072036880963|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|6d2b21b67cb000734e415bf77861c029f901c720|1.99|2014-09-25 12:55:00|1.4132775322775095|1|7203688096|82|0.6114706929155321|0|58|526|-80.97058|64|35.03469|FRESH MUSHROOMS|0.49|4|HT SLICED WHITE MUSHROOMS|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00072036880963|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|890d95f543bf4af605e086219172bccbfb5cccb2|1.99|2015-01-24 13:22:00|1.4132775322775095|1|7203688096|82|0.6114706929155321|0|58|526|-80.97058|64|35.03469|FRESH MUSHROOMS|0.0|4|HT SLICED WHITE MUSHROOMS|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00072036880963|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|8b11bd895bcbc8ba1c4f01f82b84b96982cb4ba0|3.99|2014-11-10 15:31:00|1.4132775322775095|1|7403010300|82|0.6114706929155321|0|58|321|-80.97058|53|35.03469|RICOTTA/FARMERS CHEESE|0.0|3|SORRENTO WHOLE MILK RICOTTA|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00074030103000|CULTURES|DAIRY|-80.97058|1.4132032182494703|82|1
35.03469|dc24280d0c24a253580d636051e5f12fdd5115ab|0.44|2015-01-10 14:32:00|1.4132775322775095|1||82|0.6114706929155321|0|58|534|-80.97058|64|35.03469|FRESH CHILI PEPPERS|0.0|4|COO POBLANO CHILI PEPPER|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00204701000004|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|f162c00b7f5d4d45c95ca11d3c0b6355010bb1c5|2.99|2014-12-07 10:59:00|1.4132775322775095|1||82|0.6114706929155321|0|58|561|-80.97058|64|35.03469|FR PROD ORGANIC PRODUCE|0.0|4|ORG CELERY|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00294070000002|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|39237987da747e3a1d6dced5a3ba9487f192db42|7.99|2014-12-28 15:14:00|1.4132775322775095|1|2100061161|82|0.6114706929155321|0|58|314|-80.97058|52|35.03469|CHEESE-PROCESSED-OTHER|0.0|3|KRAFT VELVEETA CHEESE|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00021000611614|CHEESE|DAIRY|-80.97058|1.4132032182494703|82|1
35.03469|9718f67d1497c4161d64d362629495b7578ae45e|3.49|2015-02-04 13:49:00|1.4132775322775095|1|82951530124|82|0.6114706929155321|0|58|1256|-80.97058|13|35.03469|WHOLESOME CRACKERS|0.4|1|SENSABLE PITA BITE SEA SALT|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00829515301248|CRACKERS|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|61167633605ee76709b698bcdb41d3b679ff5068|1.13|2015-01-17 17:31:00|1.4132775322775095|1||82|0.6114706929155321|0|58|561|-80.97058|64|35.03469|FR PROD ORGANIC PRODUCE|0.0|4|ORG YELLOW ONIONS BULK|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00294665000004|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|1a0272d276eba72be06f92fc7cce72f6162c3223|1.13|2015-01-15 16:03:00|1.4132775322775095|1||82|0.6114706929155321|0|58|561|-80.97058|64|35.03469|FR PROD ORGANIC PRODUCE|0.0|4|COO ORG RED ONIONS|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00294082000007|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|a11fbc1180378f778dbd927998828f89d26f88a2|3.99|2015-02-28 14:20:00|1.4132775322775095|1|1600043472|82|0.6114706929155321|0|58|81|-80.97058|9|35.03469|RTE CEREAL KIDS|0.0|1|GM CINNAMON TOAST CRUNCH 12.2|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00016000434721|CEREAL|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|3990631ebb9eaa35acc950231b0d34f156ee73c7|4.49|2015-02-20 18:47:00|1.4132775322775095|1|85968600400|82|0.6114706929155321|0|58|46|-80.97058|7|35.03469|PKG CHOC|0.0|1|BARKTHINS DRK ALM W/SEA SALT|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00859686004006|CANDY|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|6b372bfa06f828038d58c671643a18a3e61c93e8|2.5|2014-09-15 15:24:00|1.4132775322775095|1|6414404702|82|0.6114706929155321|0|58|179|-80.97058|27|35.03469|CANNED PASTA|0.0|1|CBRD MW BEEF RAVIOLI|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00064144047093|PREPARED FOODS-RTS|G1 GROCERY|-80.97058|1.4132032182494703|82|2
35.03469|1d4575e8ed6289d77219f26ef660e7e31baf2b2e|3.75|2015-02-01 12:06:00|1.4132775322775095|1|6414404702|82|0.6114706929155321|0|58|179|-80.97058|27|35.03469|CANNED PASTA|0.75|1|CBRD MW BEEF RAVIOLI|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00064144047093|PREPARED FOODS-RTS|G1 GROCERY|-80.97058|1.4132032182494703|82|3
35.03469|2bf40831c3382c84a5aac003b9d0cbc5e990117a|2.5|2014-12-31 12:57:00|1.4132775322775095|1|6414404702|82|0.6114706929155321|0|58|179|-80.97058|27|35.03469|CANNED PASTA|0.5|1|CBRD MW BEEF RAVIOLI|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00064144047093|PREPARED FOODS-RTS|G1 GROCERY|-80.97058|1.4132032182494703|82|2
35.03469|b1eea887170c376703035ee990e3ad5321853b53|2.5|2014-11-28 13:18:00|1.4132775322775095|1|6414404702|82|0.6114706929155321|0|58|179|-80.97058|27|35.03469|CANNED PASTA|0.5|1|CBRD MW BEEF RAVIOLI|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00064144047093|PREPARED FOODS-RTS|G1 GROCERY|-80.97058|1.4132032182494703|82|2
35.03469|b0d5889944c7c170c82242d6977c8da78d351b2d|2.5|2015-01-07 13:38:00|1.4132775322775095|1|6414404702|82|0.6114706929155321|0|58|179|-80.97058|27|35.03469|CANNED PASTA|0.5|1|CBRD MW BEEF RAVIOLI|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00064144047093|PREPARED FOODS-RTS|G1 GROCERY|-80.97058|1.4132032182494703|82|2
35.03469|0c696174ff0f75a333c27f4e784c950a8e870cde|4.29|2014-11-24 14:27:00|1.4132775322775095|1|4400003037|82|0.6114706929155321|0|58|90|-80.97058|13|35.03469|SNACK CRACKERS|2.14|1|WHEAT THIN FIBER GARDEN VEGETA|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00044000030452|CRACKERS|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|310351a3d404ced4d46ca19c5aa2a884e96b562a|3.19|2014-11-30 15:14:00|1.4132775322775095|1|4460001594|82|0.6114706929155321|0|58|399|-80.97058|69|35.03469|NFS-DISINFECTANTS|0.0|1|CLOROX DISINFECT WIPES FRESH|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00044600015934|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|ce62da17ea88f9c8a7e2249257ca492506a0e517|3.99|2014-10-01 13:51:00|1.4132775322775095|1|4400002854|82|0.6114706929155321|1|58|1248|-80.97058|12|35.03469|SANDWICH COOKIES|0.49|1|OREO GOLDEN|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00044000032586|COOKIES|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|9ec182110434287f0a4b3ce20cedba646a45cd62|3.25|2014-10-25 13:12:00|1.4132775322775095|1|4157005617|82|0.6114706929155321|0|58|1265|-80.97058|57|35.03469|ALMOND MILK|0.75|3|ALMOND BREEZE CHOCOLATE|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00041570056257|MILK|DAIRY|-80.97058|1.4132032182494703|82|1
35.03469|88e4c067ccd642a86cd5d9c17d721c2907ef5c3b|4.49|2014-10-04 12:57:00|1.4132775322775095|1|2570071147|82|0.6114706929155321|0|58|442|-80.97058|76|35.03469|NFS-COOKING-STORAGE BAGS|0.99|1|ZIPLOC SANDWICH BAGS|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00025700003915|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|48513111cc5069226dac0fc51490f2797df29d43|2.79|2014-11-08 17:38:00|1.4132775322775095|1|1800000501|82|0.6114706929155321|0|58|327|-80.97058|54|35.03469|DINNER ROLLS-REFRIGERATED|0.0|3|PILLSBURY CINN CREAM CHS ROLLS|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00018000005123|DOUGH PRODUCTS|DAIRY|-80.97058|1.4132032182494703|82|1
35.03469|ae87f35bd06663c7cf56a2c25a0b196adf50bd9b|1.69|2014-11-19 15:33:00|1.4132775322775095|1|2100065897|82|0.6114706929155321|0|58|1441|-80.97058|274|35.03469|MAC AND CHEESE|0.0|1|KRAFT MAC CHEESE NINJA TURTLE|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00021000031542|PREP FOODS DINNERS|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|4f8e1ef7e3da1810b89ac8a6fadca4774529ea7a|2.89|2015-02-19 17:25:00|1.4132775322775095|1|2733100033|82|0.6114706929155321|0|58|495|-80.97058|108|35.03469|NON REFRIGERATED|0.0|19|LA BANDERITA TORTILLA 8 INCH|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00027331000332|TORTILLAS|CASE READY MEATS|-80.97058|1.4132032182494703|82|1
35.03469|dd5c2c5d7aa9c43e0d2601ab2872a733b8d71b71|5.0|2014-10-09 15:46:00|1.4132775322775095|1|8143403117|82|0.6114706929155321|0|58|9935|-80.97058|885|35.03469|NFS POP CAB SAUV|0.0|13|REX GOLIATH CABERNET SAUVIGNON|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00081434031174|POPULAR (4-$7.99)|WINE|-80.97058|1.4132032182494703|82|1
35.03469|0f710f077f14d0aa163e8d6ae046269202f71716|19.99|2015-02-27 14:06:00|1.4132775322775095|1|8143471001|82|0.6114706929155321|0|58|9924|-80.97058|882|35.03469|NFS-PREMIUM BOX|0.0|13|BLACK BOX PINOT NOIR|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00081434710017|PREMIUM BOX|WINE|-80.97058|1.4132032182494703|82|1
35.03469|04c7d4afa88d6087949dd9aad0136e8bb0febf21|0.99|2014-11-14 15:45:00|1.4132775322775095|1||82|0.6114706929155321|0|58|540|-80.97058|64|35.03469|FRESH CELERY|0.0|4|COO CELERY (RPC) 24'S|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00204070000001|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|7540b1ee4a70fff80085db65e0ec13f36c1b87a3|9.59|2015-02-06 07:39:00|1.4132775322775095|1|9955508520|82|0.6114706929155321|0|58|37|-80.97058|10|35.03469|PODS/CUPS/SINGLES|0.0|1|CARIBOU BLEND K-CUPS|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00099555089929|COFFEE|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|d35b7941ac9147f3ad7ed789dff1e9c6c84e7860|8.79|2014-09-29 17:40:00|1.4132775322775095|1|9955508520|82|0.6114706929155321|0|58|37|-80.97058|10|35.03469|PODS/CUPS/SINGLES|0.0|1|CARIBOU BLEND K-CUPS|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00099555089929|COFFEE|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|b7951ae7bb0a9f1a94e7d31e1a248269bc5eddfd|2.99|2014-10-27 14:46:00|1.4132775322775095|1|89000000110|82|0.6114706929155321|0|58|104|-80.97058|16|35.03469|APPLESAUCE-CUPS|0.0|1|GOGO SQUEEZ 4PK APPLE MANGO|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00890000001547|FRUIT-CAN/JAR|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|a285d59ebc13e19f464026ba8b39d643994f8eb0|2.99|2014-12-04 15:52:00|1.4132775322775095|1|89000000110|82|0.6114706929155321|0|58|104|-80.97058|16|35.03469|APPLESAUCE-CUPS|0.0|1|GOGO SQUEEZ 4PK APPLE MANGO|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00890000001547|FRUIT-CAN/JAR|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|771b796f4cd93db70953b42403441ad08e1121ec|5.99|2014-10-15 20:18:00|1.4132775322775095|1|8500001444|82|0.6114706929155321|0|58|9938|-80.97058|885|35.03469|NFS POP PINOT GRS/GRIGIO|0.0|13|CB-BAREFOOT PINOT GRIGIO|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00085000014448|POPULAR (4-$7.99)|WINE|-80.97058|1.4132032182494703|82|1
35.03469|023cdbd66c502bd894b9c5517e47f400956d4954|1.98|2015-02-09 13:43:00|1.4132775322775095|1|7726000266|82|0.6114706929155321|0|58|727|-80.97058|7|35.03469|SEASONAL CANDY-SINGLE FAC|0.5|1|I/O(V15)RS DC MARSH HEART BAR|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00077260002662|CANDY|G1 GROCERY|-80.97058|1.4132032182494703|82|2
35.03469|a5850917fb5c92ca3560604c1b7d65b29cc3e4bd|3.89|2014-12-06 15:31:00|1.4132775322775095|1|7800000117|82|0.6114706929155321|0|58|55|-80.97058|8|35.03469|REGULAR|0.4|23|CANADA DRY GINGERALE|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00078000001174|CARBONATED BEVERAGES|BEVERAGE|-80.97058|1.4132032182494703|82|1
35.03469|46295a1f497c9bc4b9e95d40a25a9b872abca6b6|3.89|2014-10-23 14:25:00|1.4132775322775095|1|7800000117|82|0.6114706929155321|0|58|55|-80.97058|8|35.03469|REGULAR|0.4|23|CANADA DRY GINGERALE|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00078000001174|CARBONATED BEVERAGES|BEVERAGE|-80.97058|1.4132032182494703|82|1
35.03469|3cecef5ed7ad37c97f9acfce369a976ceeec9133|2.29|2014-12-31 16:28:00|1.4132775322775095|1|7800023046|82|0.6114706929155321|0|58|55|-80.97058|8|35.03469|REGULAR|0.79|23|CANADA DRY CBRY G/ALE 2LTR|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00078000156461|CARBONATED BEVERAGES|BEVERAGE|-80.97058|1.4132032182494703|82|1
35.03469|b8f12052342f4ce734143e1aafd79316759b868d|4.85|2014-12-23 19:41:00|1.4132775322775095|1|7790011553|82|0.6114706929155321|0|58|479|-80.97058|105|35.03469|NAT/ORG BREAKFAST SAUSAGE|1.51|19|JIMMY DEAN NATURAL SAUSGE MILD|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00077900306587|BREAKFAST SAUSAGE|CASE READY MEATS|-80.97058|1.4132032182494703|82|1
35.03469|50877b8f1caa7d5c575c340fe3144ce691204a3e|3.74|2014-12-16 18:27:00|1.4132775322775095|1|20542000000|82|0.6114706929155321|0|58|1832|-80.97058|415|35.03469|BH SLICING CHEESE|0.0|6|BOARS HEAD BABY SWISS CHEESE|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00205420000009|SLICING CHEESE|DELI|-80.97058|1.4132032182494703|82|1
35.03469|1e4be84aa907e7d1a7e86395d40db57587e186b5|2.75|2015-01-29 11:44:00|1.4132775322775095|1|20542000000|82|0.6114706929155321|0|58|1832|-80.97058|415|35.03469|BH SLICING CHEESE|0.0|6|BOARS HEAD BABY SWISS CHEESE|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00205420000009|SLICING CHEESE|DELI|-80.97058|1.4132032182494703|82|1
35.03469|72d714c72e77a37b444c3c230565d1ff179e88ea|6.39|2014-10-20 14:46:00|1.4132775322775095|1|3040077377|82|0.6114706929155321|0|58|427|-80.97058|72|35.03469|NFS-TOILET TISSUE|0.0|1|ANGEL SOFT SOFT/STRONG 12DR|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00030400773778|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|950b53e81b1bf11a4816a601e3c3efb714c5e16c|7.75|2014-11-16 17:22:00|1.4132775322775095|1|1258760034|82|0.6114706929155321|0|58|443|-80.97058|76|35.03469|NFS-GARBAGE BAGS|0.4|1|GLAD TALL KTCHN DRAWSTG 13GL|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00012587786284|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|a9acc3bb3295dc7ae07d33aa8cc5ff724ef53170|1.89|2014-11-05 10:57:00|1.4132775322775095|1|2000000065|82|0.6114706929155321|0|58|1275|-80.97058|50|35.03469|BOX VEG|0.0|5|GG EARLY JUNE PEAS BUTTER SAUC|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00020000000909|VEGETABLES-FROZEN|FROZEN|-80.97058|1.4132032182494703|82|1
35.03469|3bb394a4428bd565104d1b51f5e842ca338fac7c|2.99|2015-03-04 08:43:00|1.4132775322775095|1|74447394110|82|0.6114706929155321|0|58|341|-80.97058|57|35.03469|CREAMERS|0.0|3|SO DELICIOUS ALM MLK CRMR-ORIG|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00744473933105|MILK|DAIRY|-80.97058|1.4132032182494703|82|1
35.03469|8a5e480300d6e7e35abbd76e1ec5b09d1e27bf3b|3.29|2014-11-09 14:20:00|1.4132775322775095|1|68896200201|82|0.6114706929155321|0|58|535|-80.97058|64|35.03469|FRESH GREENS|0.0|4|BAG KALE 16 OZ|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00688962002012|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|5c98d16420978f1f81ad27940426c9d229c928f5|7.99|2014-10-19 13:15:00|1.4132775322775095|1|1186311873|82|0.6114706929155321|0|58|2019|-80.97058|505|35.03469|PRESSED COOKED CHEESE|0.0|6|SARTORI BELLAVITANO GOLD|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00011863118733|SPECIALTY CHEESE|DELI|-80.97058|1.4132032182494703|82|1
35.03469|413b3a15a7743b797d42a233e3fe3d7b79f9a8d7|15.99|2014-09-27 16:04:00|1.4132775322775095|1|1820022980|82|0.6114706929155321|0|58|463|-80.97058|84|35.03469|HARD CIDER|0.0|16|JOHNNY APPLESEED 12PK|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00018200229800|SPECIALTY|BEER|-80.97058|1.4132032182494703|82|1
35.03469|ae3026f5b55ed95ae7d28dba5ef9909a8a5850e2|1.81|2014-10-07 17:12:00|1.4132775322775095|1||82|0.6114706929155321|0|58|523|-80.97058|64|35.03469|FRESH POTATOES|0.0|4|"COO RED POTATO ""A""SIZE, BULK"|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00204073000008|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|03ad45cf88dd55050f25e8f43b2a23e509261f20|8.63|2014-09-17 18:14:00|80.970593795509558|1|20898900000|82|35.050189210146748|0|4|1421|-80.994596|201|35.061685|SMART CHICKEN VEGETABLE FED|0.0|2|SMART CHICKEN BONELESS BREAST|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|35.073829668338668|00208989000008|POULTRY|MEAT|-80.97058|80.970583268867514|475|1
35.03469|fca20c9600f5858ba3a70fbbf39fb660f207eac5|6.99|2014-12-11 15:52:00|1.4132775322775095|1|3700087406|82|0.6114706929155321|0|58|427|-80.97058|72|35.03469|NFS-TOILET TISSUE|0.0|1|CHARMIN BATH ULTRA STRONG 4MR|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00037000874393|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|6f435a6d541d8d5cc148bdc46860ec033451392f|8.59|2014-10-05 16:40:00|1.4132775322775095|1|1380014333|82|0.6114706929155321|0|58|1280|-80.97058|48|35.03469|MULTI SERVE MEALS|1.6|5|STOUFFER LASAGNA ITALIANO|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00013800143310|FROZEN MEALS|FROZEN|-80.97058|1.4132032182494703|82|1
35.03469|9bb2a31910fd38a00753c848f85bf4d4d4861108|5.99|2014-10-29 19:37:00|1.4132775322775095|1|8143403128|82|0.6114706929155321|0|58|9938|-80.97058|885|35.03469|NFS POP PINOT GRS/GRIGIO|0.0|13|CB-REX GOLIATH PINOT GRIGIO|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00081434031280|POPULAR (4-$7.99)|WINE|-80.97058|1.4132032182494703|82|1
35.03469|4b74362437c62f8372d248fa024354fb607f6417|1.01|2015-02-18 16:52:00|1.4132775322775095|1||82|0.6114706929155321|0|58|502|-80.97058|64|35.03469|FRESH BANANAS|0.0|4|BANANAS, YELLOW|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00204011000008|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|2985ea6977de689d952950a62dcfadbf2fbd203a|2.95|2014-10-12 18:53:00|1.4132775322775095|1|3800040260|82|0.6114706929155321|0|58|1269|-80.97058|41|35.03469|BREAKFAST SYRUP CARRIER|0.95|5|EGGO BLUEBERRY WAFFLES|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00038000403200|BREAKFAST FOODS FROZEN|FROZEN|-80.97058|1.4132032182494703|82|1
35.03469|23338545bde92d54d4fed7079ce95f61c45bf86e|2.65|2014-09-16 14:29:00|1.4132775322775095|1|1600015110|82|0.6114706929155321|0|58|205|-80.97058|31|35.03469|REMAINING SNACKS|0.0|1|BUGLES ORIGINAL|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00016000283701|SNACKS|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|33668a46ba9b3fc57afb7a772169efccf73dedd9|4.53|2014-09-28 17:10:00|1.4132775322775095|1||82|0.6114706929155321|0|58|529|-80.97058|64|35.03469|FRESH ASPARAGUS|0.5|4|GREEN  ASPARAGUS|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00204080000008|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|a8cac0cd44a449d042dad06557976b35fed5f944|5.99|2015-03-08 10:43:00|80.970593795509558|1|4242122579|82|35.050189210146748|0|4|358|-80.994596|100|35.061685|REGULAR BACON|1.0|19|BOARS HEAD SMOKED BACON 16 OZ|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|35.073829668338668|00042421225792|BACON|CASE READY MEATS|-80.97058|80.970583268867514|475|1
35.03469|06cd043b0e029d74417b027384cc9e2167d9639a|9.69|2014-09-11 17:01:00|1.4132775322775095|1|1780057309|82|0.6114706929155321|0|58|156|-80.97058|24|35.03469|NFS-DOG FOOD-DRY|0.0|1|PURINA ONE SM BITES BEEF &RICE|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00017800464048|PET FOOD/SUPPLIES|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|e65ff8bd39b1643a8f790235d4f0035eabcf1750|9.99|2014-11-22 15:10:00|80.970593795509558|1|8769284102|82|35.050189210146748|0|4|463|-80.994596|84|35.061685|HARD CIDER|0.0|16|ANGRY ORCHARD APPLE GINGER 6PK|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|35.073829668338668|00087692841029|SPECIALTY|BEER|-80.97058|80.970583268867514|475|1
35.03469|40ac256cc603bbed7b91028c4cc57680dd96613a|9.99|2014-11-29 14:29:00|1.4132775322775095|1|8769284102|82|0.6114706929155321|0|58|463|-80.97058|84|35.03469|HARD CIDER|0.0|16|ANGRY ORCHARD APPLE GINGER 6PK|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00087692841029|SPECIALTY|BEER|-80.97058|1.4132032182494703|82|1
35.03469|2de701381abc322896fe262a7db06bca299bfbc6|56.97|2014-09-24 13:59:00|1.4132775322775095|1|3270010875|82|0.6114706929155321|0|58|6893|-80.97058|1582|35.03469|DOG FLEA & TICK|38.160000000000004|18|HARTZ UG DROPS DOG 15LB&UNDR 3|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00032700108748|PET NEEDS|GM|-80.97058|1.4132032182494703|82|3
35.03469|9dea299fd7a19fb75d5c4bfd37fd876deeed6249|4.49|2014-10-10 18:39:00|1.4132775322775095|1|2100000900|82|0.6114706929155321|0|58|317|-80.97058|52|35.03469|CHUNK AND BAR CHEESE|0.0|3|CRACKER BARREL AGED CHUNKS|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00021000009053|CHEESE|DAIRY|-80.97058|1.4132032182494703|82|1
35.03469|b14ee037f10b553cc0ff883a04eea3b96b524948|1.19|2014-12-20 15:51:00|1.4132775322775095|1|7433686394|82|0.6114706929155321|0|58|342|-80.97058|57|35.03469|FRESH MILK|0.2|3|HUNTER 2% MILK 14 OZ|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00074336863950|MILK|DAIRY|-80.97058|1.4132032182494703|82|1
35.03469|e95e55e3e0b99d475a00879f79442fcd0d9bf16e|13.99|2014-10-04 16:04:00|1.4132775322775095|1|1820005990|82|0.6114706929155321|0|58|456|-80.97058|82|35.03469|DOMESTIC SUPER PREM 12PK&>|0.0|16|MICHELOB ULTRA 12PK 12OZ BTL|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00018200059902|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|077ab1cc76cad2f5283a391bfcba55395625a328|8.34|2014-10-26 11:16:00|1.4132775322775095|1|7203624015|82|0.6114706929155321|0|58|149|-80.97058|23|35.03469|WHSE PASTA CORE|2.52|1|HT PASTA SPAGHETTI 16|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00072036240156|PASTA|G1 GROCERY|-80.97058|1.4132032182494703|82|6
35.03469|21dc7d2bc0ef97869f58218319d10b361b42bd72|8.99|2014-10-17 15:55:00|1.4132775322775095|1|7023666033|82|0.6114706929155321|0|58|751|-80.97058|87|35.03469|NFS-BOUQUETS|0.0|9|$9.99  SPRING HOT SPOT|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00070236660330|FLORAL|FLORAL|-80.97058|1.4132032182494703|82|1
35.03469|224a5401db4397ec4d125be0a43900204efa8025|3.34|2014-12-19 12:42:00|1.4132775322775095|1|7203643010|82|0.6114706929155321|0|58|252|-80.97058|45|35.03469|PREMIUM ICE CREAM|0.0|5|HT PREM FUDGE RIPPLE IC|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00072036430168|ICE CREAM|FROZEN|-80.97058|1.4132032182494703|82|1
35.03469|47833d8b5a9c016ba7f989f69e801602ebc76694|12.46|2014-09-27 16:03:00|1.4132775322775095|1|20891800000|82|0.6114706929155321|0|58|657|-80.97058|201|35.03469|STR MDE VALUE ADD POLTRY|1.56|2|HNY/GINGER MRTND CHICKEN KABOB|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00208997000007|POULTRY|MEAT|-80.97058|1.4132032182494703|82|1
35.03469|8f6e715d1bf7a2cc45a26a18967479236524262d|10.99|2015-02-06 18:12:00|1.4132775322775095|1|8224229043|82|0.6114706929155321|0|58|9948|-80.97058|886|35.03469|NFS-PREM-CAB SAUVIGNON|0.0|13|GNARLY HEAD CABERNET SAUV|268b13b72d435151fdf392445abe7e8b27086726|1.0709580078542191|0.61177642288969325|00082242290432|PREMIUM ($8-$10.99)|WINE|-80.97058|1.4132032182494703|82|1
35.297134|f779fe5e321ef9a718ba313bd51b471f2eeea497|4.36|2014-10-20 18:04:00|1.4094857484078087|4||258|0.6160512048176361|0|26|502|-80.737839|64|35.297134|FRESH BANANAS|0.0|4|BANANAS, YELLOW|2e12d05a2593a6e78bf80e96bb228e3cb685ddd3|2.994242260631064|0.61471665291522548|00204011000008|FRESH PRODUCE|PRODUCE|-80.737839|1.409141121495086|258|1
35.297134|68cd3d337590c0bed852eebb231d0e76ce940285|6.85|2014-12-24 15:28:00|80.737901233649083|4|7192147763|258|35.340467527203799|0|46|284|-80.764523|892|35.341927|SUPER PREMIUM PIZZA|0.0|5|12in CAL. P/K TC BBQ CHICKEN|2e12d05a2593a6e78bf80e96bb228e3cb685ddd3|2.994242260631064|35.349871187060224|00071921624910|FROZEN PIZZA|FROZEN|-80.737839|80.737857290208069|220|1
35.297134|93738a6146248fbdd4245d6f484296a6057a042d|6.87|2014-09-25 23:20:00|1.4094857484078087|4|61126999100|258|0.6160512048176361|0|26|97|-80.737839|8|35.297134|ENERGY DRINKS|0.62|23|CB RED BULL ENERGY DRINK|2e12d05a2593a6e78bf80e96bb228e3cb685ddd3|2.994242260631064|0.61471665291522548|00611269991000|CARBONATED BEVERAGES|BEVERAGE|-80.737839|1.409141121495086|258|3
35.297134|799f7701be72205f04bb6e2b614d7a2a4eb2bab9|10.0|2014-10-09 14:27:00|1.4094857484078087|4||258|0.6160512048176361|0|26|512|-80.737839|64|35.297134|FRSH PROD FRSH FRUIT REM|0.0|4|MANGOS|2e12d05a2593a6e78bf80e96bb228e3cb685ddd3|2.994242260631064|0.61471665291522548|00204959000009|FRESH PRODUCE|PRODUCE|-80.737839|1.409141121495086|258|10
35.297134|b29439463ed3648f8a81f058633ae7d408fdada9|1.79|2015-01-06 22:58:00|1.4094857484078087|4|7160300448|258|0.6160512048176361|0|26|3103|-80.737839|1000|35.297134|MPLEMENTS NAIL-TRIM|0.0|17|*** TRIM DLX TOENL CLIP W/FILE|2e12d05a2593a6e78bf80e96bb228e3cb685ddd3|2.994242260631064|0.61471665291522548|00071603004481|COSMETICS|HBC|-80.737839|1.409141121495086|258|1
35.297134|849a476d209f922cf41b7dfa9223e87c5671bfe8|19.99|2014-11-14 17:58:00|1.4094857484078087|4|7203695593|258|0.6160512048176361|0|26|1653|-80.737839|381|35.297134|CELEBRATION CAKES|0.0|14|1/4 DL CHOC CK W WH BUTTRCRM|2e12d05a2593a6e78bf80e96bb228e3cb685ddd3|2.994242260631064|0.61471665291522548|00072036955937|CAKES|BAKERY|-80.737839|1.409141121495086|258|1
34.937113|bfb61f0722fb57c92e2bdb03b88c14e0abd7b6d1|15.99|2015-03-06 17:55:00|80.811922674510953|4|7203661034|372|34.981159183582683|0|12|666|-80.816172|145|35.059823|PACKAGED COOKED|0.0|12|HT COOKED SHRIMP RING 20OZ|304da6c65387d08b4014e5e4b788adba86a7ccd6|3.0434878025527294|35.037868710371079|00072036610348|SHRIMP|SEAFOOD|-80.837892|80.837965995956537|66|1
35.43259|987d41b9bed85e40d9cec769758ef4a0cdafe13a|1.5|2015-03-06 10:55:00|80.606823361882718|3|68954408130|202|35.50838580377652|0|57|685|-80.662946|61|35.412407|GREEK|0.5|3|FAGE TOTAL 2% STRAWBERRY|31bf6bcf965f6cd69782cbfb7814a7fcb3a6be71|5.237307583973766|35.500309569604553|00689544081463|YOGURT|DAIRY|-80.605588|80.605631925590089|68|1
35.43259|336856e3bbdf7befa13b0560b61abb6c457c798f|3.95|2015-02-15 19:12:00|1.4057311447477159|3|1410007467|202|0.6184153580092175|0|52|1025|-80.605588|162|35.43259|WHITE|0.95|7|PEP FH SOURDOUGH WP BRD PP|31bf6bcf965f6cd69782cbfb7814a7fcb3a6be71|5.237307583973766|0.6209993146566879|00014100074670|SLICED BREAD|COMMERCIAL BAKERY|-80.605588|1.406832906106031|202|1
35.43259|14d9686747ca6ad3e10d9cda63f5834ccbdc3563|7.3|2015-03-01 12:09:00|80.606823361882718|3|3010001610|202|35.50838580377652|0|57|1254|-80.662946|12|35.412407|FUDGE ENROBED|1.15|1|FUDGE SHOPPE GRASSHOPPER MINT|31bf6bcf965f6cd69782cbfb7814a7fcb3a6be71|5.237307583973766|35.500309569604553|00030100440574|COOKIES|G1 GROCERY|-80.605588|80.605631925590089|68|2
35.43259|54dad034c133e9eb5ce42831d9c8b37b6a1ea408|2.69|2014-12-23 08:40:00|1.4057311447477159|3|7116904049|202|0.6184153580092175|0|52|18|-80.605588|3|35.43259|CAKE DECORATIONS & ICING|0.0|1|CM CUPCAKE LINERS - WHITE|31bf6bcf965f6cd69782cbfb7814a7fcb3a6be71|5.237307583973766|0.6209993146566879|00071169040497|BAKING SUPPLIES|G1 GROCERY|-80.605588|1.406832906106031|202|1
35.43259|272d72f8afb8829e072771b619d8ddeb7204bd06|2.69|2015-01-26 14:51:00|80.606823361882718|3|7116904049|202|35.50838580377652|0|57|18|-80.662946|3|35.412407|CAKE DECORATIONS & ICING|0.0|1|CM CUPCAKE LINERS - WHITE|31bf6bcf965f6cd69782cbfb7814a7fcb3a6be71|5.237307583973766|35.500309569604553|00071169040497|BAKING SUPPLIES|G1 GROCERY|-80.605588|80.605631925590089|68|1
35.43259|cb2a2db92dd2a31160872c0d38bb372aebb309a1|8.98|2014-09-12 10:50:00|1.4057311447477159|3|2840009217|202|0.6184153580092175|0|52|1981|-80.605588|480|35.43259|CHIPS|0.0|6|STACY'S PITA CHIPS NAKED|31bf6bcf965f6cd69782cbfb7814a7fcb3a6be71|5.237307583973766|0.6209993146566879|00028400092173|DRY GOODS|DELI|-80.605588|1.406832906106031|202|2
35.43259|793f965562455eaaf033527d55066a816daf993b|1.65|2015-01-31 12:53:00|80.606823361882718|3|2920000212|202|35.50838580377652|0|57|1208|-80.662946|23|35.412407|WHSE PASTA VALUE ADD|0.65|1|MUELLER WG ELBOW MAC|31bf6bcf965f6cd69782cbfb7814a7fcb3a6be71|5.237307583973766|35.500309569604553|00029200001709|PASTA|G1 GROCERY|-80.605588|80.605631925590089|68|1
35.43259|7fc42240a018c8ba3f27487fe12dd6a05de9ceb9|3.99|2015-02-25 15:56:00|80.606823361882718|3|2529300122|202|35.50838580377652|0|57|1266|-80.662946|57|35.412407|COCONUT MILK|0.99|3|SILK COCONUT UNSWEET 64 OZ|31bf6bcf965f6cd69782cbfb7814a7fcb3a6be71|5.237307583973766|35.500309569604553|00025293002289|MILK|DAIRY|-80.605588|80.605631925590089|68|1
35.43259|98b6670d53e7bea11a3cc712b33fb3b2fc24f631|23.97|2015-01-08 11:38:00|80.606823361882718|3|7203676196|202|35.50838580377652|0|57|35|-80.662946|10|35.412407|PREMIUM WHOLE BEAN|7.26|1|HT TRADER COFFEE WB FR ROAST|31bf6bcf965f6cd69782cbfb7814a7fcb3a6be71|5.237307583973766|35.500309569604553|00072036762016|COFFEE|G1 GROCERY|-80.605588|80.605631925590089|68|3
35.43259|8fc54de11379a425426950026ff357621476c684|0.99|2014-12-17 16:08:00|1.4057311447477159|3|7203695306|202|0.6184153580092175|0|52|1895|-80.605588|450|35.43259|TEA|0.0|6|FFM LEMONADE|31bf6bcf965f6cd69782cbfb7814a7fcb3a6be71|5.237307583973766|0.6209993146566879|00072036953070|BEVERAGES|DELI|-80.605588|1.406832906106031|202|1
35.43259|2e46cc9d8ae69285abf22c1a80c739b54e157afe|15.98|2015-01-11 14:01:00|1.4057311447477159|3|7203676196|202|0.6184153580092175|0|52|35|-80.605588|10|35.43259|PREMIUM WHOLE BEAN|2.42|1|HT TRADER COFFEE WB COL SUPREM|31bf6bcf965f6cd69782cbfb7814a7fcb3a6be71|5.237307583973766|0.6209993146566879|00072036761989|COFFEE|G1 GROCERY|-80.605588|1.406832906106031|202|2
35.43259|d2f224660395377b9f9564b505cee8c16dbf127a|2.49|2014-12-20 11:10:00|1.4057311447477159|3|7203688048|202|0.6184153580092175|0|52|526|-80.605588|64|35.43259|FRESH MUSHROOMS|0.0|4|HT SLICED BABY BELLAS|31bf6bcf965f6cd69782cbfb7814a7fcb3a6be71|5.237307583973766|0.6209993146566879|00072036880482|FRESH PRODUCE|PRODUCE|-80.605588|1.406832906106031|202|1
35.43259|7dd7e7c6f2b3703979f96216f4db3c9f2caa02a7|4.98|2014-11-09 21:35:00|80.606823361882718|3|7203688048|202|35.50838580377652|0|57|526|-80.662946|64|35.412407|FRESH MUSHROOMS|0.98|4|HT SLICED BABY BELLAS|31bf6bcf965f6cd69782cbfb7814a7fcb3a6be71|5.237307583973766|35.500309569604553|00072036880482|FRESH PRODUCE|PRODUCE|-80.605588|80.605631925590089|68|2
35.43259|fbdf853f4189516007a9b4bdc2d939204364e6c6|3.58|2015-01-15 18:09:00|1.4057311447477159|3|74447390901|202|0.6184153580092175|0|52|687|-80.605588|61|35.43259|BLENDED|0.54|3|SO DELICIOUS ALM MILK CHOCOLAT|31bf6bcf965f6cd69782cbfb7814a7fcb3a6be71|5.237307583973766|0.6209993146566879|00744473909551|YOGURT|DAIRY|-80.605588|1.406832906106031|202|2
35.43259|d3be717ae82813c383503e31f240956e6ee0d5c4|25.9|2014-12-18 15:04:00|80.606823361882718|3|20129900000|202|35.50838580377652|0|57|296|-80.662946|49|35.412407|RANCHER BEEF|10.84|2|VALUE PK BEEF LOIN STRIP STEAK|31bf6bcf965f6cd69782cbfb7814a7fcb3a6be71|5.237307583973766|35.500309569604553|00201299000003|BEEF|MEAT|-80.605588|80.605631925590089|68|1
35.43259|51637467e2dbea90623315fb796f00bb844768bd|1.85|2014-10-07 10:18:00|1.4057311447477159|3|5100002457|202|0.6184153580092175|0|52|212|-80.605588|33|35.43259|CONDENSED SOUP|0.85|1|CAMP COND CREAM OF POTATO|31bf6bcf965f6cd69782cbfb7814a7fcb3a6be71|5.237307583973766|0.6209993146566879|00051000016416|SOUP|G1 GROCERY|-80.605588|1.406832906106031|202|1
35.43259|577f3d34f2592f5053019acfb6d98d3cffeab66b|4.98|2014-09-30 11:08:00|1.4057311447477159|3|7373107000|202|0.6184153580092175|0|52|495|-80.605588|108|35.43259|NON REFRIGERATED|1.49|19|MISSION FAJITA 8 CT|31bf6bcf965f6cd69782cbfb7814a7fcb3a6be71|5.237307583973766|0.6209993146566879|00073731070000|TORTILLAS|CASE READY MEATS|-80.605588|1.406832906106031|202|2
35.603432|4fde3604734e044fad466749c8aac03a7631bed5|5.69|2014-10-31 18:07:00|80.891462859624312|2|7756725423|274|35.634808173632528|0|45|252|-80.860108|45|35.500972|PREMIUM ICE CREAM|2.85|5|BREYERS FRENCH VANILLA I/C|321d19e0f9387bac7d012c77e423ceecea41c4d4|2.1680187109843985|35.636605227883024|00077567254382|ICE CREAM|FROZEN|-80.895009|80.895043849862759|268|1
35.603432|addf4c61eafdaa69649a3e5b2580849938f73844|1.47|2014-10-05 10:36:00|80.891462859624312|2|20575500000|274|35.634808173632528|0|45|1603|-80.860108|371|35.500972|PRIVATE LABEL BREAD|0.0|14|WHEAT BAGUETTE ROUNDS|321d19e0f9387bac7d012c77e423ceecea41c4d4|2.1680187109843985|35.636605227883024|00205760000004|BREAD|BAKERY|-80.895009|80.895043849862759|268|1
35.603432|60638311ef550e4af215fb4b60991b8251969bca|1.76|2015-01-10 14:51:00|80.891462859624312|2|20575500000|274|35.634808173632528|0|45|1603|-80.860108|371|35.500972|PRIVATE LABEL BREAD|0.0|14|WHEAT BAGUETTE ROUNDS|321d19e0f9387bac7d012c77e423ceecea41c4d4|2.1680187109843985|35.636605227883024|00205760000004|BREAD|BAKERY|-80.895009|80.895043849862759|268|1
35.603432|68954617f8881af116b21b21607bd004f4ef9d5c|17.98|2014-10-10 17:14:00|80.891462859624312|2|61278110261|274|35.634808173632528|0|45|265|-80.860108|307|35.500972|FROZEN PIES|4.0|5|M CALLENDER DUTCH APPLE PIE|321d19e0f9387bac7d012c77e423ceecea41c4d4|2.1680187109843985|35.636605227883024|00612781101205|DESSERTS FROZEN|FROZEN|-80.895009|80.895043849862759|268|2
35.603432|9a07a36c258bf0ae1187e879c83bbe4c7b5ab256|3.99|2014-09-20 17:38:00|80.891462859624312|2|64034401028|274|35.634808173632528|0|45|581|-80.860108|136|35.500972|FRESH SALSA|0.0|4|FRESH CUTS MILD SALSA|321d19e0f9387bac7d012c77e423ceecea41c4d4|2.1680187109843985|35.636605227883024|00640344010282|OTHER MERCHANDISE|PRODUCE|-80.895009|80.895043849862759|268|1
35.603432|f74d853fd883df7251cb12c15e158560f0c8f650|2.5|2014-10-04 17:16:00|80.891462859624312|2|78142100610|274|35.634808173632528|0|45|1601|-80.860108|371|35.500972|BRANDED BREAD|0.51|14|LA BREA FRENCH BAGUETTE|321d19e0f9387bac7d012c77e423ceecea41c4d4|2.1680187109843985|35.636605227883024|00781421006108|BREAD|BAKERY|-80.895009|80.895043849862759|268|1
35.603432|210b604b8dcd97a18c7bd455cf0d00926a447d3b|2.99|2015-02-26 16:30:00|80.891462859624312|2|76857303100|274|35.634808173632528|0|45|544|-80.860108|64|35.500972|FRESH PRODUCE FRSH HERBS|0.0|4|ORGANIC LIVING BASIL|321d19e0f9387bac7d012c77e423ceecea41c4d4|2.1680187109843985|35.636605227883024|00768573031004|FRESH PRODUCE|PRODUCE|-80.895009|80.895043849862759|268|1
35.603432|522478532be4697c9f1f88b7d6916e6c3a3e7d53|3.98|2014-09-13 17:12:00|80.891462859624312|2|64420900438|274|35.634808173632528|0|45|24|-80.860108|3|35.500972|FROSTING-READY-TO-SPREAD|0.0|1|DH BUTTERCREME FROSTING|321d19e0f9387bac7d012c77e423ceecea41c4d4|2.1680187109843985|35.636605227883024|00644209471041|BAKING SUPPLIES|G1 GROCERY|-80.895009|80.895043849862759|268|2
35.603432|f33f16289d43c70a989c9381d4ca1e54971b35a6|3.99|2014-09-22 16:27:00|80.891462859624312|2|5783602085|274|35.634808173632528|0|45|522|-80.860108|64|35.500972|FRESH TOMATOES|0.0|4|GOURMET MEDLEY TOMATOES 12 OZ|321d19e0f9387bac7d012c77e423ceecea41c4d4|2.1680187109843985|35.636605227883024|00885773044013|FRESH PRODUCE|PRODUCE|-80.895009|80.895043849862759|268|1
35.603432|9cbcedd0ebb1a01e75bc7dd884161428fbdd32c9|7.99|2015-01-02 17:15:00|80.891462859624312|2|3798212040|274|35.634808186283443|0|45|2016|-80.875654|505|35.585842|SOFT RIPENED|0.0|6|BRIE  7.7 OZ|321d19e0f9387bac7d012c77e423ceecea41c4d4|2.1680187109843985|35.636605227883024|00037982120402|SPECIALTY CHEESE|DELI|-80.895009|80.895012627663064|99|1
35.603432|891dbe38dd00d236ec4f7f0bbc13193b6b870b6b|14.98|2014-11-21 19:14:00|80.891462859624312|2|7203695788|274|35.634808173632528|0|45|1403|-80.860108|389|35.500972|THAW AND SELL PIES|5.0|14|"8"" PECAN PIE"|321d19e0f9387bac7d012c77e423ceecea41c4d4|2.1680187109843985|35.636605227883024|00072036957887|PIES|BAKERY|-80.895009|80.895043849862759|268|2
35.603432|88132c021955c1b2784f661799d26e509636c731|8.99|2014-09-23 17:51:00|80.891462859624312|2|7203695149|274|35.634808173632528|0|45|1937|-80.860108|465|35.500972|COLD PREP FOODS ENTREES|0.0|6|SPINACH & CHEESE QUICHE|321d19e0f9387bac7d012c77e423ceecea41c4d4|2.1680187109843985|35.636605227883024|00072036951465|COLD PREPARED FOODS|DELI|-80.895009|80.895043849862759|268|1
35.603432|cc6932a6528d5e1b481b10147f0ca8df98264456|6.55|2014-12-27 19:04:00|80.891462859624312|2|7570616502|274|35.634808186283443|0|45|254|-80.875654|892|35.585842|PREMIUM PIZZA|2.56|5|PALERMOS PRIMO SPIN/BCN/FETA|321d19e0f9387bac7d012c77e423ceecea41c4d4|2.1680187109843985|35.636605227883024|00075706165193|FROZEN PIZZA|FROZEN|-80.895009|80.895012627663064|99|1
35.603432|fa8aec7163a2610a224e1e4be3d1cf69a5e13f55|2.85|2014-12-09 17:40:00|80.891462859624312|4|4133500053|274|35.623061275341918|0|45|184|-80.861571|28|35.444615|SALAD DRESSINGS-LIQUID|0.0|1|KENS DRS LT VIN BALSMIC BASIL|365551915c3d0ebdf8804d88a2b3498cd03b6467|1.356337036915008|35.636605227883024|00041335329558|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.895009|80.895045074168038|340|1
35.603432|b030849ac779600351645b3b835b024141c98c35|5.41|2014-10-31 09:35:00|1.4102725052409182|4||274|0.6213971134099097|0|1|503|-80.895009|64|35.603432|FRESH GRAPES|0.36|4|GREEN GRAPES, SEEDLESS 12/16|365551915c3d0ebdf8804d88a2b3498cd03b6467|1.356337036915008|0.61833652052202714|00204022000004|FRESH PRODUCE|PRODUCE|-80.895009|1.4118842554804456|274|1
35.603432|88361698505f741108e397e2d610641c6cea1d48|1.37|2015-02-23 20:21:00|1.4102725052409182|4||274|0.6213971134099097|0|1|502|-80.895009|64|35.603432|FRESH BANANAS|0.0|4|BANANAS, YELLOW|365551915c3d0ebdf8804d88a2b3498cd03b6467|1.356337036915008|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.895009|1.4118842554804456|274|1
35.603432|3c9ebc1f3acd8277738e863e4df8962c2f3efd22|11.850000000000001|2014-12-27 16:20:00|1.4102725052409182|4|74816261452|274|0.6213971134099097|0|1|1460|-80.895009|40|35.603432|FROZEN BREAD AND ROLLS|4.35|5|SCHUBERTS PARKERHOUSE ROLLS|365551915c3d0ebdf8804d88a2b3498cd03b6467|1.356337036915008|0.61833652052202714|00748162614528|FROZEN DOUGH|FROZEN|-80.895009|1.4118842554804456|274|3
35.603432|51dd6d6ed81195d368493b8c094f6e4535c09cd5|1.54|2015-01-20 20:15:00|1.4102725052409182|4||274|0.6213971134099097|0|1|502|-80.895009|64|35.603432|FRESH BANANAS|0.0|4|BANANAS, YELLOW|365551915c3d0ebdf8804d88a2b3498cd03b6467|1.356337036915008|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.895009|1.4118842554804456|274|1
35.603432|81e382c54cedcf7a32f7e397f032db89daf92970|2.99|2014-10-06 20:13:00|1.4102725052409182|4|7203688212|274|0.6213971134099097|0|1|555|-80.895009|64|35.603432|PACKAGED SALADS|0.0|4|HT SPRING MIX|365551915c3d0ebdf8804d88a2b3498cd03b6467|1.356337036915008|0.61833652052202714|00072036882127|FRESH PRODUCE|PRODUCE|-80.895009|1.4118842554804456|274|1
35.500972|38b8d6ef732b05c58f11535124a20d9281dbc4a3|4.0|2015-02-12 15:20:00|80.8939826282094|4|66440100015|268|35.528684232767787|0|2|1165|-80.875654|87|35.585842|NFS-FRESH CONSUMER BUNCH|0.0|9|BUNCH- HYPERIUCM ASST.|3850e91bebb5843715171e7728da7fbd46faa94c|1.9148489880663908|35.490689277687849|00664401000153|FLORAL|FLORAL|-80.860108|80.86013553971955|99|1
35.500972|b5af65c7ca07a6e226cf11a4a6a97f978c7da79e|0.95|2015-02-18 21:08:00|80.8939826282094|4|7203663222|268|35.528684232767787|0|2|330|-80.875654|55|35.585842|EGGS|0.0|3|HT GRADE A    LARGE EGGS 6 CT.|3850e91bebb5843715171e7728da7fbd46faa94c|1.9148489880663908|35.490689277687849|00072036632227|EGGS FRESH|DAIRY|-80.860108|80.86013553971955|99|1
35.500972|4d5b29be82bfccf47b75a5aca0c9431c65b6548d|3.49|2015-03-08 17:50:00|80.8939826282094|4|7203670903|268|35.528684232767787|0|2|214|-80.875654|33|35.585842|BROTH|0.49|1|HARRIS TEETER CHICK BROTH 48OZ|3850e91bebb5843715171e7728da7fbd46faa94c|1.9148489880663908|35.490689277687849|00072036709035|SOUP|G1 GROCERY|-80.860108|80.86013553971955|99|1
35.500972|184282340dfe09a1ac1239a3340af57c83fc1ed1|0.89|2015-02-12 20:10:00|80.8939826282094|4|2310001401|268|35.528684232767787|0|2|158|-80.875654|24|35.585842|NFS-DOG FOOD-WET|0.09|1|CESAR PORK TENDERLOIN|3850e91bebb5843715171e7728da7fbd46faa94c|1.9148489880663908|35.490689277687849|00023100056739|PET FOOD/SUPPLIES|G1 GROCERY|-80.860108|80.86013553971955|99|1
35.500972|e1ed62f42b262340030cba2fd81ccb909c959f1b|4.45|2015-03-07 18:45:00|80.8939826282094|4|2310001401|268|35.528684232767787|0|2|158|-80.875654|24|35.585842|NFS-DOG FOOD-WET|0.09|1|CESAR SELECT W/TURKEY|3850e91bebb5843715171e7728da7fbd46faa94c|1.9148489880663908|35.490689277687849|00023100014074|PET FOOD/SUPPLIES|G1 GROCERY|-80.860108|80.86013553971955|99|5
35.667941|45f8a52d27a3d228181bfe1ad9a8c1dc9faad649|6.39|2015-02-21 13:49:00|1.4057311447477159|4|7430500132|178|0.6225230078570788|0|52|82|-80.497332|11|35.667941|VINEGAR|0.0|1|BRAGG ORG VINEGAR APPLE CIDER|3a16ce0183b997ed8d90112e5f8b3387393d14e9|5.633443184298055|0.6209993146566879|00074305001321|CONDIMENTS|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|29248e8c1fee78107c405913670948bb46485cf8|6.38|2014-12-10 13:30:00|1.4057311447477159|4|74759960098|178|0.6225230078570788|0|52|16|-80.497332|3|35.667941|BAKING CHOCOLATE/CHIPS/MORSELS|0.69|1|GHIRADELLI BAR BITTERSWEET 60%|3a16ce0183b997ed8d90112e5f8b3387393d14e9|5.633443184298055|0.6209993146566879|00747599601125|BAKING SUPPLIES|G1 GROCERY|-80.497332|1.4049434824709919|178|2
35.341927|9e1aa7b5947b180ce8858b2e4872d6a59f27402e|2.85|2015-03-05 11:57:00|80.779636304526477|4|3000031186|220|35.378319383012219|0|17|42|-80.860108|6|35.500972|GRANOLA/YOGURT BARS|0.0|1|QUAKER CHEWY LS CHOC CHIP|3c994cb91b3aafa26c5049249b50fd1a277e04ee|2.51462764169963|35.392509581117899|00030000311752|BREAKFAST FOODS|G1 GROCERY|-80.764523|80.764577275849348|268|1
35.341927|ad6ffb4e4fb52b63795c718e0d990bbf7a687e94|5.98|2015-01-17 11:40:00|80.779636304526477|4|3338365583|220|35.378319409358774|0|17|522|-80.66939|64|35.28326|FRESH TOMATOES|0.98|4|SWEET GRAPE TOMATO (PINT)|3c994cb91b3aafa26c5049249b50fd1a277e04ee|2.51462764169963|35.392509581117899|00072036880284|FRESH PRODUCE|PRODUCE|-80.764523|80.764530912447285|46|2
35.341927|3430489d88d256f2fa8823bc691e9ef95c5b93ba|1.49|2015-01-19 15:04:00|80.779636304526477|4|7618316374|220|35.378319408699802|0|17|99|-80.86175|32|35.40953|LIQUID TEA|0.49|1|SNAPPLE ICE TEA|3c994cb91b3aafa26c5049249b50fd1a277e04ee|2.51462764169963|35.392509581117899|00076183163740|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.764523|80.764534606983958|209|1
35.341927|92fb414ab3cc420e11a47c8b860f4dd238b488b5|5.79|2014-09-15 20:25:00|80.779636304526477|4|2100060260|220|35.378319383012219|0|17|315|-80.860108|52|35.500972|CHEESE-PROCESSED-SLICED|0.0|3|KRAFT DELI DELUXE SLICES|3c994cb91b3aafa26c5049249b50fd1a277e04ee|2.51462764169963|35.392509581117899|00021000602605|CHEESE|DAIRY|-80.764523|80.764577275849348|268|1
35.341927|c93cf5563b3223af68a39637ca2c3a13299d08fd|6.19|2014-09-15 21:20:00|80.779636304526477|4|30573016420|220|35.378319383012219|0|17|4347|-80.860108|1205|35.500972|PAIN RELIEVER & SLEEP AID|0.0|17|ADVIL PM CAPLETS|3c994cb91b3aafa26c5049249b50fd1a277e04ee|2.51462764169963|35.392509581117899|00305730164207|PAIN RELIEF|HBC|-80.764523|80.764577275849348|268|1
35.103409|72c9dff56305fc4d77614beaa9202c3ce327b5b9|5.69|2015-02-05 09:05:00|1.4132775322775095|2|2410010523|88|0.6126700657242101|0|58|1252|-80.992182|12|35.103409|LUNCH BOX COOKIES|0.0|1|KBLR VARIETY CHE RAINBW MINI|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00030100940371|COOKIES|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|e2d10c476abff43a8258a86a013f9ae93a9c7cb8|3.69|2015-02-21 17:26:00|1.4132775322775095|2|2500005542|88|0.6126700657242101|0|58|334|-80.992182|56|35.103409|GRAPEFRUIT JUICE-REGRIGERATED|0.0|3|SIMPLY GRAPEFRUIT|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00025000054501|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|6d4c42bbacb18002383920a2b1e89f619c7439b1|4.69|2015-02-19 20:05:00|1.4132775322775095|2|3736300612|88|0.6126700657242101|0|58|1279|-80.992182|48|35.103409|SINGLE SERVE FLAVOR|1.19|5|MICH ANGELO LASAGNA W/MEAT SC|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00037363006127|FROZEN MEALS|FROZEN|-80.992182|1.413580244274486|88|1
35.103409|9bf180be2ea968264d92e1684f7b14c7da453f70|9.4|2014-11-02 17:33:00|1.4132775322775095|2|20220200000|88|0.6126700657242101|0|58|299|-80.992182|49|35.103409|ANGUS BEEF|0.0|2|ANGUS BEEF FILET MIGNON CUSTOM|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00202209000007|BEEF|MEAT|-80.992182|1.413580244274486|88|1
35.103409|ff67d3240149539aaf41f7e98c60bf0200d97072|3.89|2015-03-01 16:21:00|80.992238315890603|2|7457000400|88|35.128336268594701|0|22|275|-80.945176|45|35.323246|SUPER PREMIUM ICE CREAM|0.0|5|H DAZS BUTTER PECAN-|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|35.131650835559327|00074570114009|ICE CREAM|FROZEN|-80.992182|80.99225806093078|166|1
35.103409|1c2a104a3d4a149deca66fa1def915899ccc792a|7.18|2015-01-30 17:13:00|1.4132775322775095|2|7765208254|88|0.6126700657242101|0|58|233|-80.992182|37|35.103409|BLACK TEA|1.18|1|STASH TEA BLACK DOUBLE SPICE|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00077652082654|TEA|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|a1946371f6b7dea2b5327e7464e8fff5a02991bc|7.18|2015-01-30 06:07:00|1.4132775322775095|2|7765208254|88|0.6126700657242101|0|58|233|-80.992182|37|35.103409|BLACK TEA|0.59|1|STASH TEA BLACK DOUBLE SPICE|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00077652082654|TEA|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|ce7f02c09f6469d3e6841816ffd2d6632cf1d0f1|3.59|2014-09-11 16:41:00|1.4132775322775095|2|7765208254|88|0.6126700657242101|0|58|233|-80.992182|37|35.103409|BLACK TEA|0.6|1|STASH TEA BLACK DOUBLE SPICE|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00077652082654|TEA|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|fbe8efc92f5dfb234d5da6b0220d858a7b173c94|4.7|2014-12-22 17:46:00|1.4132775322775095|2|7365121422|88|0.6126700657242101|0|58|160|-80.992182|25|35.103409|OLIVES|1.18|1|MARIO OLIVE RIPE MEDIUM.|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00073651214225|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|386715a991170e85e1cf245698d4a133116c49b5|8.99|2014-12-19 20:56:00|80.992238315890603|2|7203688112|88|35.128336339317826|0|22|583|-80.85753|136|35.116638|NUTS|0.0|4|HT PECAN HALVES TRAY|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|35.131650835559327|00072036881120|OTHER MERCHANDISE|PRODUCE|-80.992182|80.992204710199573|204|1
35.103409|4aa26931f2ca619d4c6e604c66d953f3000389c7|1.69|2015-02-25 21:19:00|1.4132775322775095|2|7203688003|88|0.6126700657242101|0|58|527|-80.992182|64|35.103409|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00072036880031|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|1
35.103409|5b126cf97fb59961cbd5ee41de9d51a5882123a9|1.69|2014-09-17 09:07:00|1.4132775322775095|2|7203688003|88|0.6126700657242101|0|58|527|-80.992182|64|35.103409|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00072036880031|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|1
35.103409|b2719a1b390cbb69fea13213e7fa62cb7809d524|1.69|2015-01-25 19:18:00|1.4132775322775095|2|7203688003|88|0.6126700657242101|0|58|527|-80.992182|64|35.103409|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00072036880031|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|1
35.103409|e15d8742cd5b99dc9767e6f448ce5d327c5bc1dc|12.99|2015-01-13 13:06:00|80.992238315890603|2|7203695587|88|35.128336343430789|0|22|1707|-80.770346|387|35.052812|MESSAGE|3.0|14|12 INCH MESSAGE COOKIE|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|35.131650835559327|00072036955876|COOKIES|BAKERY|-80.992182|80.992196467209283|40|1
35.103409|ff9573a7d8ac9a8abfe00682144c1f8b39b27aa6|6.95|2014-11-27 13:43:00|1.4132775322775095|2|3760048620|88|0.6126700657242101|0|58|358|-80.992182|100|35.103409|REGULAR BACON|0.0|19|HORMEL BLACK LABEL LOW SALT|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00037600486200|BACON|CASE READY MEATS|-80.992182|1.413580244274486|88|1
35.103409|a7fffa671b16f53cfe274d4820c7b53fe8a93f62|9.97|2015-01-27 19:39:00|1.4132775322775095|2|3700086514|88|0.6126700657242101|0|58|427|-80.992182|72|35.103409|NFS-TOILET TISSUE|0.0|1|CHARMIN BATH ULTRA SOFT 24DR|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00037000851233|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|0375dd71253842c037ff8789a80c0b5be230a822|0.64|2015-02-06 06:11:00|1.4132775322775095|2||88|0.6126700657242101|0|58|502|-80.992182|64|35.103409|FRESH BANANAS|0.0|4|BANANAS, YELLOW|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00204011000008|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|1
35.103409|213dd4cda1f482a2d33c8556471ccb50e9a5a4ce|3.58|2014-10-16 12:07:00|1.4132775322775095|2|1500007430|88|0.6126700657242101|0|58|1257|-80.992182|1|35.103409|POUCH BABY FOOD|0.58|1|GERBER 2ND ORG BAN ACIA GRANOL|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00015000074456|BABY FOOD|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|212a384908174d9fddc17df201fdad9ac40bae67|1.79|2014-09-18 08:16:00|1.4132775322775095|2|1500007430|88|0.6126700657242101|0|58|1257|-80.992182|1|35.103409|POUCH BABY FOOD|0.45|1|GERBER 2ND ORGANC APPLE BLKBRY|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00015000074357|BABY FOOD|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|15f7a6fe31cfac5577791f70045c9057d2629707|4.99|2015-02-08 16:11:00|1.4132775322775095|2|7430000070|88|0.6126700657242101|0|58|5188|-80.992182|1305|35.103409|BABY OINTMENTS|0.0|17|DESITIN OINTMENT   -00070|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00074300000701|BABY HBC|HBC|-80.992182|1.413580244274486|88|1
35.103409|c339ed6776f1190ecd876f357125349996111190|6.98|2015-01-16 11:05:00|1.4132775322775095|2|2840023981|88|0.6126700657242101|0|58|203|-80.992182|31|35.103409|CHEESE SNACKS|1.74|1|CHEETOS JUMBO PUFFS|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00028400239875|SNACKS|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|3fded03e04f0d1cb3d3e82f04f941c005fd7ef84|11.3|2015-02-21 18:26:00|1.4132775322775095|2|4470007502|88|0.6126700657242101|0|58|484|-80.992182|101|35.103409|BEEF WIENERS|2.83|19|OSCAR MAYER JUMBO BEEF FRANK|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00044700073377|WIENERS|CASE READY MEATS|-80.992182|1.413580244274486|88|2
35.103409|66d6cfa9ff706bff6886ecbf8c6b7e88c20bd66c|2.69|2015-01-30 19:24:00|1.4132775322775095|2||88|0.6126700657242101|0|58|528|-80.992182|64|35.103409|FRESH BROCCOLI|0.0|4|COO BROCCOLI, BUN 25# (RPC)|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00204060000004|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|1
35.103409|b875791bbe2394e74a2fc2371c6d5a181493a008|12.99|2014-12-24 10:06:00|80.992238315890603|2|8210073851|88|35.128336344793674|0|22|9948|-80.816172|886|35.059823|NFS-PREM-CAB SAUVIGNON|0.0|13|THE DREAMING TREE CABERNET|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|35.131650835559327|00082100738519|PREMIUM ($8-$10.99)|WINE|-80.992182|80.992192380416611|66|1
35.103409|eee7931c9fa7cd4253a381e753dc1103bd905f51|8.530000000000001|2015-03-07 12:23:00|1.4132775322775095|2|20165700000|88|0.6126700657242101|0|58|297|-80.992182|49|35.103409|GROUND BEEF|1.0|2|HT GROUND BEEF CHUCK 80% LEAN|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00201657000003|BEEF|MEAT|-80.992182|1.413580244274486|88|2
35.103409|d1eb93fa8a7462da7eb20031c59fc2b42bb38837|6.87|2015-03-08 13:07:00|1.4132775322775095|2|1450001098|88|0.6126700657242101|0|58|1275|-80.992182|50|35.103409|BOX VEG|0.95|5|BE STEAMFRESH MIXED VEGES|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00014500011282|VEGETABLES-FROZEN|FROZEN|-80.992182|1.413580244274486|88|3
35.103409|7f520895233fca91cf01602a276483ec2c62445b|2.29|2015-02-16 17:42:00|1.4132775322775095|2|2670012915|88|0.6126700657242101|0|58|1267|-80.992182|53|35.103409|DIPS AND SPREADS|0.79|3|DEAN'S LITE FRENCH ONION DIP|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00026700322006|CULTURES|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|a00e13764720cbae181a04d50c009b39ad8c3fdb|2.85|2015-03-04 11:45:00|1.4132775322775095|2|1380010321|88|0.6126700657242101|0|58|1279|-80.992182|48|35.103409|SINGLE SERVE FLAVOR|0.0|5|STOUF MAC&BEEF W/TOMATOES|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00013800447845|FROZEN MEALS|FROZEN|-80.992182|1.413580244274486|88|1
35.103409|3a004de3d99b8b074197cc248319e5591756c244|7.16|2014-09-20 19:05:00|1.4132775322775095|2|1500007430|88|0.6126700657242101|0|58|1257|-80.992182|1|35.103409|POUCH BABY FOOD|0.46|1|GERBER 2ND ORG AP MAG RICE VAN|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00015000074463|BABY FOOD|G1 GROCERY|-80.992182|1.413580244274486|88|4
35.103409|dec64c807b20832a52d0ca4ff2a33ad7eeb65197|4.19|2014-10-11 15:41:00|1.4132775322775095|2|2100062503|88|0.6126700657242101|0|58|318|-80.992182|52|35.103409|SHREDDED/GRATED CHEESE|1.69|3|KRAFT 2% SHARP SHRED|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00021000024605|CHEESE|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|4f9305fb187420ce0f4d2f801e168f1cda5ff8f1|4.25|2015-02-01 13:24:00|1.4132775322775095|2|2840023186|88|0.6126700657242101|0|58|199|-80.992182|31|35.103409|DIPS & SALSAS|0.0|1|RUFFLES CREAMY BUF RNCH DIP|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00028400231862|SNACKS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|3e738b3eda818c2d5715d0020ec7c7ee0ec929b4|4.25|2014-12-10 20:24:00|1.4132775322775095|2|2840023186|88|0.6126700657242101|0|58|199|-80.992182|31|35.103409|DIPS & SALSAS|0.0|1|RUFFLES CREAMY BUF RNCH DIP|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00028400231862|SNACKS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|30bc6509a8107faa063a75285fb0ac9e8f106ffc|4.25|2015-01-19 20:27:00|1.4132775322775095|2|2840023186|88|0.6126700657242101|0|58|199|-80.992182|31|35.103409|DIPS & SALSAS|0.0|1|RUFFLES CREAMY BUF RNCH DIP|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00028400231862|SNACKS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|78e89055145069f8f5a7b646613f67ea5d6f5bf5|7.79|2015-03-04 20:40:00|80.992238315890603|2|30045027125|88|35.128336268594701|0|22|4236|-80.945176|1200|35.323246|DEX ADULT/CHILDREN|0.0|17|TYL SEVERE COLD/FLU CAPLETS|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|35.131650835559327|00300450270269|COUGH/COLD/SINUS|HBC|-80.992182|80.99225806093078|166|1
35.103409|e10bd6b2c6a52f108eb04f27d986062d281bf4b1|5.99|2015-02-15 13:13:00|1.4132775322775095|2|2100002492|88|0.6126700657242101|0|58|315|-80.992182|52|35.103409|CHEESE-PROCESSED-SLICED|2.0|3|KRAFT 2% AMERICAN SINGLE|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00021000024926|CHEESE|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|0fe2d551638fa911cdcdd997f91e8583758fb720|4.99|2014-12-20 17:31:00|1.4132775322775095|2|2840008313|88|0.6126700657242101|0|58|204|-80.992182|31|35.103409|TORTILLA CHIPS|1.0|1|TOSTITOS RSTC FAMILY SIZE|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00028400083133|SNACKS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|c5172f5db88529c1b1874426bed8106d6ef1380e|7.55|2015-03-02 21:34:00|1.4132775322775095|2|3100067010|88|0.6126700657242101|0|58|1280|-80.992182|48|35.103409|MULTI SERVE MEALS|0.56|5|PF CHANG SHANGHAI BEEF|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00031000670009|FROZEN MEALS|FROZEN|-80.992182|1.413580244274486|88|1
35.103409|e927193940fa24a455c297d89fa04cec727b88af|5.38|2014-10-05 19:46:00|1.4132775322775095|2|20597100000|88|0.6126700657242101|0|58|1821|-80.992182|410|35.103409|BH TURKEY|0.0|6|BOARS HEAD LOW SODIUM TURKEY|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00205971000008|BH MEAT|DELI|-80.992182|1.413580244274486|88|1
35.103409|9e282c3da05a2343481f8294de5df649c2d72c35|3.98|2014-10-04 15:57:00|80.992238315890603|2|7203648011|88|35.128336343430789|0|22|274|-80.770346|44|35.052812|ICE|0.0|5|HT BAGGED ICE 10LB (456)|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|35.131650835559327|00000000004560|ICE|FROZEN|-80.992182|80.992196467209283|40|2
35.103409|7f6e1ebc6d1de9109e08b90340fde9a41d1ca661|10.99|2014-10-18 19:09:00|1.4132775322775095|2|1338590127|88|0.6126700657242101|0|58|9958|-80.992182|886|35.103409|NFS-PREM-OTHER WHITE|0.0|13|BILTMORE SEASONAL|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00013385901275|PREMIUM ($8-$10.99)|WINE|-80.992182|1.413580244274486|88|1
35.103409|b292f6eac43455944f958cd0c952f89c409e10d5|4.99|2015-01-31 08:14:00|1.4132775322775095|2|1111018700|88|0.6126700657242101|0|58|1647|-80.992182|379|35.103409|PACKAGED MUFFINS|1.02|14|FFM 4 CT BLUEBERRY MUFFIN|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00011110187000|MUFFINS|BAKERY|-80.992182|1.413580244274486|88|1
35.103409|e003d1082b87774532c899e8caf41f9f342bccfe|1.69|2014-11-21 11:17:00|1.4132775322775095|2|1200000129|88|0.6126700657242101|0|58|55|-80.992182|8|35.103409|REGULAR|0.0|23|CB PEPSI COLA 20 0Z|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00012000001291|CARBONATED BEVERAGES|BEVERAGE|-80.992182|1.413580244274486|88|1
35.103409|fd9f86517e779d0726c7920ca5bc5641058bcb7c|3.58|2014-10-20 17:16:00|1.4132775322775095|2|1500007430|88|0.6126700657242101|0|58|1257|-80.992182|1|35.103409|POUCH BABY FOOD|0.29|1|GERBER 2ND ORG BAN BLUE BLACKB|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00015000074449|BABY FOOD|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|8b66367eee6e8d898890e62de9ffd9ee81ad642a|1.79|2015-01-10 20:41:00|1.4132775322775095|2|85686200311|88|0.6126700657242101|0|58|3939|-80.992182|1075|35.103409|SHAVING CREAM MEN-CREAM|0.0|17|BRUT CLASSIC SHAVE FOAM|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00856862003112|SHAVING NEEDS/MEN HAIR|HBC|-80.992182|1.413580244274486|88|1
35.103409|0860601c7655610bc5addadf5ca19acf9cb1c8a5|2.99|2015-01-31 18:21:00|1.4132775322775095|2|1340008242|88|0.6126700657242101|0|58|239|-80.992182|38|35.103409|RICE-PACKAGED & BULK|0.0|1|COMET RICE WHITE|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00013400082422|RICE GRAINS AND BEANS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|c5be62e4a85bf99ddea87254678b1acea134b4bb|8.99|2014-10-28 18:07:00|1.4132775322775095|2|8769230050|88|0.6126700657242101|0|58|458|-80.992182|82|35.103409|CRAFT BEER|0.0|16|SAM ADAMS SEASONAL 6PK|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00087692300502|DOMESTIC BEER|BEER|-80.992182|1.413580244274486|88|1
35.103409|6edbf409ea59c61696dcee2a7ccd40ba5f62530b|5.49|2015-02-09 19:17:00|1.4132775322775095|2|3680022087|88|0.6126700657242101|0|58|4338|-80.992182|1205|35.103409|PAIN RELIEVER-CHILDREN|0.0|17|TC IBU SUSP BERRY|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00036800220874|PAIN RELIEF|HBC|-80.992182|1.413580244274486|88|1
35.103409|e160ff29e53694fb6ff41ca80baf6bdc736f47fc|5.09|2015-01-21 20:27:00|1.4132775322775095|2|3680013444|88|0.6126700657242101|0|58|4189|-80.992182|1200|35.103409|ALLERGY REMEDY-CHILDREN|0.0|17|TC CHILDREN  ALLERGY-CHERRY|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00036800134447|COUGH/COLD/SINUS|HBC|-80.992182|1.413580244274486|88|1
35.103409|dc507330406d935fc5f8196af32bbd9f35f5053f|19.99|2014-12-11 08:55:00|80.992238315890603|2|7203695893|88|35.128336344793674|0|22|1653|-80.816172|381|35.059823|CELEBRATION CAKES|0.0|14|1/4 DL WHT CAKE / WHT BUTCREAM|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|35.131650835559327|00072036958938|CAKES|BAKERY|-80.992182|80.992192380416611|66|1
35.103409|19eb8ff1e5c130822166a6b35d59db02d8daee82|5.99|2015-02-04 22:11:00|1.4132775322775095|2|7203695041|88|0.6126700657242101|0|58|1654|-80.992182|381|35.103409|DESSERT CAKES|0.0|14|2 CT. CHOC OVERLOAD TORTE|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00072036950413|CAKES|BAKERY|-80.992182|1.413580244274486|88|1
35.103409|f07ffa73c7f08a0e2e9b8a7ec0463da227647e1c|5.99|2015-01-16 20:03:00|1.4132775322775095|2|7203695041|88|0.6126700657242101|0|58|1654|-80.992182|381|35.103409|DESSERT CAKES|0.0|14|2 CT. CHOC OVERLOAD TORTE|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00072036950413|CAKES|BAKERY|-80.992182|1.413580244274486|88|1
35.103409|9abec9c7771989c928982df65748d12a33904ade|34.99|2014-12-17 07:42:00|80.992238315890603|2|7203695496|88|35.128336344793674|0|22|1653|-80.816172|381|35.059823|CELEBRATION CAKES|0.0|14|1/2 SHT DL WHITE CAKE W/BUTCR|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|35.131650835559327|00072036954961|CAKES|BAKERY|-80.992182|80.992192380416611|66|1
35.103409|cd5e2576b77f3efae4c3ae2da8b2605d2b05b5c0|0.97|2014-12-16 11:16:00|80.992238315890603|2|7203698758|88|35.128335951326136|0|22|31|-80.895009|4|35.603432|NON CARBONATED WATER|0.0|1|HT SPRING WATER|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|35.131650835559327|00072036987587|BOTTLED WATER|G1 GROCERY|-80.992182|80.99235353557772|274|1
35.103409|30b74f9317193c804073e9c6bf599f18283a4564|1.79|2014-09-22 21:11:00|1.4132775322775095|2|85686200311|88|0.6126700657242101|0|58|3939|-80.992182|1075|35.103409|SHAVING CREAM MEN-CREAM|0.0|17|BRUT REVOLUTION SHAVE FOAM|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00856862003105|SHAVING NEEDS/MEN HAIR|HBC|-80.992182|1.413580244274486|88|1
35.103409|8cab2fe0140a5d579ab8cb15d0f1089d0746cbda|2.99|2014-12-27 19:45:00|1.4132775322775095|2|61300873513|88|0.6126700657242101|0|58|99|-80.992182|32|35.103409|LIQUID TEA|0.0|1|ARNOLD PALMER LITE TEA|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00613008720858|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|7f6f4eaf5079fed9ef9dc01285f0edcf3d91b458|6.87|2014-10-04 19:14:00|80.992238315890603|2|61126999100|88|35.128336345633599|0|22|97|-80.760919|8|35.024332|ENERGY DRINKS|0.62|23|CB RED BULL ENERGY DRINK|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|35.131650835559327|00611269991000|CARBONATED BEVERAGES|BEVERAGE|-80.992182|80.992188720954516|343|3
35.103409|c4ed4c8ff2e00ef18784075fb65c5454f65ae37d|2.69|2014-09-26 18:59:00|1.4132775322775095|2|61300873513|88|0.6126700657242101|0|58|99|-80.992182|32|35.103409|LIQUID TEA|0.0|1|ARNOLD PALMER LITE TEA|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00613008720858|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|a2868490ea0f99d7d7f9e113ae3e34857b73ca95|2.69|2014-10-01 20:40:00|1.4132775322775095|2|61300873513|88|0.6126700657242101|0|58|99|-80.992182|32|35.103409|LIQUID TEA|0.0|1|ARNOLD PALMER LITE TEA|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00613008720858|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|6533b91faff3458c2e6e1016b05cf849a4f0293b|2.69|2014-10-21 21:40:00|1.4132775322775095|2|61300873513|88|0.6126700657242101|0|58|99|-80.992182|32|35.103409|LIQUID TEA|0.0|1|ARNOLD PALMER LITE TEA|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00613008720858|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|62cb4bf5a86bf1ea6d6f1c99171c5f4d18166f42|2.99|2014-11-15 16:45:00|1.4132775322775095|2|61300873513|88|0.6126700657242101|0|58|99|-80.992182|32|35.103409|LIQUID TEA|0.0|1|ARNOLD PALMER LITE TEA|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00613008720858|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|5d32cf57ea8cce71e69089e6ec298b4a79481243|2.69|2014-09-20 17:02:00|1.4132775322775095|2|61300873513|88|0.6126700657242101|0|58|99|-80.992182|32|35.103409|LIQUID TEA|0.0|1|ARNOLD PALMER LITE TEA|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00613008720858|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|2ed1e7677af8d82f609cb513b1e0476b2203ea7a|2.69|2014-10-13 20:39:00|1.4132775322775095|2|61300873513|88|0.6126700657242101|0|58|99|-80.992182|32|35.103409|LIQUID TEA|0.0|1|ARNOLD PALMER LITE TEA|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00613008720858|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|614960d74548a77d931c6d6d47e2e27bfc49dc97|11.68|2015-02-22 17:28:00|1.4132775322775095|2|20165900000|88|0.6126700657242101|0|58|297|-80.992182|49|35.103409|GROUND BEEF|1.95|2|GROUND BEEF 93% LEAN|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00201659000001|BEEF|MEAT|-80.992182|1.413580244274486|88|2
35.103409|52f575f0591f9e12662e2540cc6f7cf9a5685cec|9.78|2014-09-10 08:47:00|1.4132775322775095|2|7261346022|88|0.6126700657242101|0|58|417|-80.992182|71|35.103409|NFS-FABRIC SOFTENERS|1.89|1|ALL FABRIC SOFTENER SHEET 80CT|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00072613460229|LAUNDRY SUPPLIES|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|70be2e9d1ff48771d36d31a20ffe9e46642170b6|2.99|2015-02-14 17:27:00|1.4132775322775095|2|7726009248|88|0.6126700657242101|0|58|727|-80.992182|7|35.103409|SEASONAL CANDY-SINGLE FAC|0.49|1|I/O(V15)RS TWEEN HEART|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00077260092489|CANDY|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|c5c4ab1d9450a4eec3fd2d4c212f418d8c8480c4|19.99|2014-12-06 19:49:00|80.992238315890603|2|85516500507|88|35.128336268594701|0|22|9981|-80.945176|888|35.323246|NFS-U/PREM-OTHER RED|0.0|13|MEIOMI SONOMA PINOT NOIR|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|35.131650835559327|00855165005076|ULTRA PREMIUM ($15-$19.99)|WINE|-80.992182|80.99225806093078|166|1
35.103409|6e59eff08e62249f1345be47b984670cde11067b|2.79|2014-11-18 06:24:00|1.4132775322775095|2|5000092917|88|0.6126700657242101|0|58|341|-80.992182|57|35.103409|CREAMERS|0.79|3|I/OCOFFEEMATE RUM CAKE|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00050000929177|MILK|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|7de8c0e59656cd88cc4fe995eccafd1c6e17a553|6.99|2015-01-29 20:04:00|1.4132775322775095|2|4900002890|88|0.6126700657242101|0|58|55|-80.992182|8|35.103409|REGULAR|6.99|23|CHERRY COKE 12OZ 12PK FP CAN|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00049000031034|CARBONATED BEVERAGES|BEVERAGE|-80.992182|1.413580244274486|88|1
35.103409|5e2b5abab8605a7c6d24621b2b19a9eecafbdda8|5.99|2015-03-06 15:19:00|1.4132775322775095|2|7756725423|88|0.6126700657242101|0|58|252|-80.992182|45|35.103409|PREMIUM ICE CREAM|1.41|5|BREYERS S&D VANILLA I/C|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00077567281302|ICE CREAM|FROZEN|-80.992182|1.413580244274486|88|1
35.103409|ad2f4694bc80f4c0da651c6cc30fc157f86c2009|1.29|2014-12-14 12:12:00|80.992238315890603|2|8379152001|88|35.128336309919597|0|22|1981|-80.826724|480|35.195689|CHIPS|0.0|6|DIRTY POT CHIP LIGHTLY SALTED|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|35.131650835559327|00083791520018|DRY GOODS|DELI|-80.992182|80.992234021046201|412|1
35.103409|f8d68f47edb4310f45617b3cdf9a680e0d1346c3|3.99|2014-10-15 11:31:00|1.4132775322775095|2|7203695939|88|0.6126700657242101|0|58|1641|-80.992182|377|35.103409|PACKAGED DONUTS|0.5|14|PUMPKIN DONUT HOLES|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00072036959393|DONUTS|BAKERY|-80.992182|1.413580244274486|88|1
35.103409|f75a04d533f2df210ffb228655eedff380767c88|3.89|2014-10-12 07:51:00|1.4132775322775095|2|61126954601|88|0.6126700657242101|0|58|97|-80.992182|8|35.103409|ENERGY DRINKS|0.0|23|CB RED BULL SUPER SLEEK 16 OZ|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00611269546019|CARBONATED BEVERAGES|BEVERAGE|-80.992182|1.413580244274486|88|1
35.103409|237e09e8afb58c151a74182a8d150f9a9688ddd6|2.99|2014-11-18 15:36:00|1.4132775322775095|2|1380016610|88|0.6126700657242101|0|58|1278|-80.992182|48|35.103409|SINGLE SERVE NUTRITIONAL|0.0|5|LC ASPARAGUS CHS RAVIOLI|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00013800557292|FROZEN MEALS|FROZEN|-80.992182|1.413580244274486|88|1
35.103409|9f4ab347f0799173e2618581dd175d934a432abd|13.99|2014-11-12 17:47:00|1.4132775322775095|2|8500001773|88|0.6126700657242101|0|58|9983|-80.992182|889|35.103409|NFS-SPARKLING|0.0|13|CB-LA MARCA PROSECCO|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00085000017739|SPARKLING|WINE|-80.992182|1.413580244274486|88|1
35.103409|b4197412fba74ca6c7c7e84239aa58267a39d2f7|1.59|2015-01-20 11:14:00|1.4132775322775095|2|7800005240|88|0.6126700657242101|0|58|55|-80.992182|8|35.103409|REGULAR|0.25|23|A&W ROOTBEER 20OZ|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00078000052404|CARBONATED BEVERAGES|BEVERAGE|-80.992182|1.413580244274486|88|1
35.103409|8e72a3008c819c53dd62df934c332709339661d7|6.99|2015-01-05 06:16:00|1.4132775322775095|2|5000025117|88|0.6126700657242101|0|58|341|-80.992182|57|35.103409|CREAMERS|0.81|3|COFFEE-MATE ITAL SWT CREAM LIQ|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00050000605354|MILK|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|3761be75242ef934251fb16c0cba0172264fc99f|3.97|2015-03-02 20:51:00|1.4132775322775095|2|7203640052|88|0.6126700657242101|0|58|231|-80.992182|37|35.103409|INSTANT TEA|0.0|1|HT ICED TEA MIX|40862e6f39847af7ac20e16f57d87ae819667111|1.7224194277868072|0.61177642288969325|00072036400529|TEA|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.43259|14c12f8e8856be10ea29b3310df277acaea776f7|3.49|2015-01-09 12:41:00|80.606823361882718|2|7800000117|202|35.50077063756757|0|57|55|-80.875654|8|35.585842|REGULAR|0.0|23|CANADA DRY GINGERALE|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00078000001174|CARBONATED BEVERAGES|BEVERAGE|-80.605588|80.605617967200075|99|1
35.43259|45b0ccd6cca190da86d8609de19e80c444cd9782|0.99|2014-12-26 15:41:00|80.606823361882718|2|7339000780|202|35.500770634342871|0|57|48|-80.662946|7|35.412407|REGISTER GUM|0.0|1|(FE)MENTOS ROLLS SPEARMINT|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00073390007805|CANDY|G1 GROCERY|-80.605588|80.605627508662138|68|1
35.43259|93e2f688adea89ebbfd3d4ef7bfc7f11e35acdf5|0.99|2015-01-31 11:53:00|80.606823361882718|2|7339000780|202|35.500770634342871|0|57|48|-80.662946|7|35.412407|REGISTER GUM|0.0|1|(FE)MENTOS ROLLS SPEARMINT|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00073390007805|CANDY|G1 GROCERY|-80.605588|80.605627508662138|68|1
35.43259|5101a40e1bf69c70836b786658b5ccb1ee0ff866|19.98|2014-11-21 14:46:00|80.606823361882718|2|8158401310|202|35.50077063756757|0|57|9959|-80.875654|887|35.585842|NFS-S/PREM-CHARDONNAY|0.0|13|CB-K. JACKSON V.R. CHARDONNAY|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00081584013105|SUPER PREMIUM ($11-$14.99)|WINE|-80.605588|80.605617967200075|99|2
35.43259|3e04cb67fca430aef29e41c35b7f02d7c6013e40|0.99|2014-10-05 18:19:00|80.606823361882718|2|7339000780|202|35.50077063756757|0|57|48|-80.875654|7|35.585842|REGISTER GUM|0.0|1|(FE)MENTOS ROLLS SPEARMINT|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00073390007805|CANDY|G1 GROCERY|-80.605588|80.605617967200075|99|1
35.43259|65995779983c72e4d2f29119ebc76f3df8b59b50|1.15|2014-12-04 09:33:00|80.606823361882718|2|20401100000|202|35.50077063756757|0|57|502|-80.875654|64|35.585842|FRESH BANANAS|0.0|4|CHIQUITA BANANAS, YELLOW|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00074904040110|FRESH PRODUCE|PRODUCE|-80.605588|80.605617967200075|99|1
35.43259|6755afa5960545097946d38abbad8bbfc267bd38|1.67|2014-12-11 12:07:00|80.606823361882718|2||202|35.50077063756757|0|57|501|-80.875654|64|35.585842|FRESH PEARS|0.0|4|RED PEARS|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00204417000008|FRESH PRODUCE|PRODUCE|-80.605588|80.605617967200075|99|1
35.43259|2c1e2413ff09bd2b009fca67486b106c13808a41|1.45|2014-12-06 15:59:00|80.606823361882718|2||202|35.50077063756757|0|57|501|-80.875654|64|35.585842|FRESH PEARS|0.0|4|ANJOU PEARS|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00204416000009|FRESH PRODUCE|PRODUCE|-80.605588|80.605617967200075|99|1
35.43259|30ece7fc6577d94a4110da1a3a67e0a95a56672b|0.98|2014-11-25 12:17:00|80.606823361882718|2||202|35.50077063756757|0|57|501|-80.875654|64|35.585842|FRESH PEARS|0.0|4|ANJOU PEARS|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00204416000009|FRESH PRODUCE|PRODUCE|-80.605588|80.605617967200075|99|1
35.43259|2ff446ea64e8e1480841bebd5f51e04bce2fecc7|14.95|2014-10-30 10:09:00|80.606823361882718|2|20136900000|202|35.50077063756757|0|57|296|-80.875654|49|35.585842|RANCHER BEEF|6.8|2|BEEF LOIN T-BONE STEAK|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00201369000001|BEEF|MEAT|-80.605588|80.605617967200075|99|1
35.43259|cbc0aa33170fbfd53723c0f0bdbce60e094feae8|1.33|2014-09-12 13:13:00|80.606823361882718|2|89470001004|202|35.50077063756757|0|57|685|-80.875654|61|35.585842|GREEK|0.33|3|CHOBANI NF POMEGRANATE|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00894700010151|YOGURT|DAIRY|-80.605588|80.605617967200075|99|1
35.43259|405b624200d2f5e1fff475da8bcfa7601e4172fd|10.99|2014-11-15 12:10:00|80.606823361882718|2|1813820102|202|35.50077063756757|0|57|9959|-80.875654|887|35.585842|NFS-S/PREM-CHARDONNAY|2.02|13|CB-EDNA VALLEY CHARDONNAY|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00018138201022|SUPER PREMIUM ($11-$14.99)|WINE|-80.605588|80.605617967200075|99|1
35.43259|332a70e0f8e847344703beea832321e1f1f77ddc|1.89|2015-02-27 10:12:00|80.606823361882718|2|31254662380|202|35.50077063756757|0|57|4207|-80.875654|1200|35.585842|COUGH DROP-ADULT|0.39|17|HALLS STRAWBERRY     -62380|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00312546623804|COUGH/COLD/SINUS|HBC|-80.605588|80.605617967200075|99|1
35.43259|f692483ec484d1c6eb3eebe4f5d5cad1c2d434da|3.49|2015-02-07 14:03:00|80.606823361882718|2|8912522000|202|35.50077063756757|0|57|151|-80.875654|23|35.585842|DSD PASTA CORE|0.5|1|ANCIENT HRVST ORG QN LINGUINI.|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00089125230004|PASTA|G1 GROCERY|-80.605588|80.605617967200075|99|1
35.43259|050282f40bc651a595dc9d27ceeff49b06cd9fac|3.49|2015-01-28 17:28:00|80.606823361882718|2|8912522000|202|35.50077063756757|0|57|151|-80.875654|23|35.585842|DSD PASTA CORE|0.5|1|ANCIENT HRVST ORG QUIN SPAGHT|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00089125250002|PASTA|G1 GROCERY|-80.605588|80.605617967200075|99|1
35.43259|9fc1a27ea87175b81640f0e5aac349afd36041df|1.99|2015-03-07 11:21:00|80.606823361882718|2|60322422423|202|35.50077063756757|0|57|533|-80.875654|64|35.585842|FRESH PEPPERS|0.0|4|MINI SWEET PEPPERS 1LB|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00603224224230|FRESH PRODUCE|PRODUCE|-80.605588|80.605617967200075|99|1
35.43259|e88589e8a29aa4b12c3f6ad625f5fa55c8ec864e|2.99|2015-01-10 11:32:00|80.606823361882718|2|7203670574|202|35.500770634342871|0|57|46|-80.662946|7|35.412407|PKG CHOC|0.49|1|HTT CHOC COVERED RAISINS|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00072036705754|CANDY|G1 GROCERY|-80.605588|80.605627508662138|68|1
35.43259|046b4dff8e6e154a0530cd958a109e8f8c61ca13|6.99|2015-02-13 08:48:00|80.606823361882718|2|7203670967|202|35.50077063756757|0|57|37|-80.875654|10|35.585842|PODS/CUPS/SINGLES|1.99|1|HT HOUSE BLEND K-CUP|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00072036709684|COFFEE|G1 GROCERY|-80.605588|80.605617967200075|99|1
35.43259|f29618093cf8bc5934c969546d3d93a56f8b2ab4|4.99|2014-10-23 10:05:00|80.606823361882718|2|8265750406|202|35.50077063756757|0|57|31|-80.875654|4|35.585842|NON CARBONATED WATER|1.0|1|(U)DEER PARK WATER 24PK .5LT|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00082657504063|BOTTLED WATER|G1 GROCERY|-80.605588|80.605617967200075|99|1
35.43259|a46acc47378a46f0df0dcf79cb9d011786b584f1|8.49|2014-09-27 10:50:00|80.606823361882718|2|78260516150|202|35.50077063756757|0|57|37|-80.875654|10|35.585842|PODS/CUPS/SINGLES|2.5|1|CHOCK FON K-CUP SOHO MORNING|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00071038012181|COFFEE|G1 GROCERY|-80.605588|80.605617967200075|99|1
35.43259|624b72e884f741b6a2fab4d6b32fc61ba189e9b6|1.57|2014-09-25 13:24:00|80.606823361882718|2|7203601075|202|35.50077063756757|0|57|1267|-80.875654|53|35.585842|DIPS AND SPREADS|0.0|3|HT FRENCH ONION DIP 16 OZ|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00072036010759|CULTURES|DAIRY|-80.605588|80.605617967200075|99|1
35.43259|670eefdc5be9359c3185087f95f75409f4387a75|3.49|2015-03-03 14:46:00|80.606823361882718|2|3010000133|202|35.50077063756757|0|57|88|-80.875654|13|35.585842|FLAKED SODA CRACKERS|0.99|1|ZESTA ORIGINAL|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00030100001331|CRACKERS|G1 GROCERY|-80.605588|80.605617967200075|99|1
35.43259|d762ae63840edf3cbd5dc97d94fd9ed8a582ea5d|9.99|2014-11-02 13:33:00|80.606823361882718|2|7050109220|202|35.500770620614382|0|57|3527|-80.746334|1045|35.41832|HAIR CARE SHPOO-MED|0.0|17|NEUTROGENA T/GEL SHAMPOO|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00070501092200|HAIR & SCALP CARE|HBC|-80.605588|80.60565420495395|190|1
35.43259|95fb323caea405e7346486e00baa20d1448a76f9|1.49|2014-11-06 15:25:00|80.606823361882718|2||202|35.50077063756757|0|57|501|-80.875654|64|35.585842|FRESH PEARS|0.0|4|RED PEARS|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00233118000000|FRESH PRODUCE|PRODUCE|-80.605588|80.605617967200075|99|1
35.43259|230dd3b7d30667f77cba223b2dc7811eb1087a31|17.58|2014-10-28 15:47:00|80.606823361882718|2|9955508520|202|35.50077063756757|0|57|37|-80.875654|10|35.585842|PODS/CUPS/SINGLES|4.39|1|GRN MTN DONUT SHOP DECAF KCUPS|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00099555085273|COFFEE|G1 GROCERY|-80.605588|80.605617967200075|99|2
35.43259|afd0d1a44a1d1188bc3c205d50e63de8fea31c7e|17.98|2014-10-31 15:28:00|80.606823361882718|2|8500001819|202|35.50077063756757|0|57|9955|-80.875654|886|35.585842|NFS-PREM-MALBEC|1.02|13|ALAMOS MENDOZA MALBEC|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00085000018194|PREMIUM ($8-$10.99)|WINE|-80.605588|80.605617967200075|99|2
35.43259|d87eac3e97d74a4245ec085e23d84cb8afcde49e|8.99|2014-10-31 15:29:00|80.606823361882718|2|8500001819|202|35.50077063756757|0|57|9955|-80.875654|886|35.585842|NFS-PREM-MALBEC|0.0|13|ALAMOS MENDOZA MALBEC|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00085000018194|PREMIUM ($8-$10.99)|WINE|-80.605588|80.605617967200075|99|1
35.43259|bb89be373d716d6eee04ba825f931a1fbe958f21|39.74|2014-11-24 11:39:00|80.606823361882718|2|20000800000|202|35.50077063756757|0|57|974|-80.875654|201|35.585842|FRESH TURKEY|11.98|2|HT FRESH TOM TURKEY 16-20 LB|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00200008000006|POULTRY|MEAT|-80.605588|80.605617967200075|99|1
35.43259|acc5de81787fc210a8d604bab02ab01825084e24|9.98|2014-12-20 17:27:00|80.606823361882718|2|3993800645|202|35.50077063497185|0|57|7407|-80.895009|1600|35.603432|CHRISTMAS PARTY GOODS/DECOR|1.98|18|PLASTIC TABLECOVER|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00039938006532|SEASONAL MERCHANDISE|GM|-80.605588|80.605625836955667|274|2
35.43259|a83afa019916b88f04c0d0d5d4dcb8ef3dd3c753|0.99|2014-12-01 16:41:00|80.606823361882718|2|7339000780|202|35.500770634342871|0|57|48|-80.662946|7|35.412407|REGISTER GUM|0.1|1|MENTOS MINT ROLL 15CT|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00073390000110|CANDY|G1 GROCERY|-80.605588|80.605627508662138|68|1
35.43259|4c6c473791a5c6dc7c7fd0291329799232b59591|6.99|2014-12-20 16:44:00|80.606823361882718|2|3770032228|202|35.50077063756757|0|57|423|-80.875654|72|35.585842|NFS-DISPOSE PLATES/BOWLS|2.0|1|CHINET PLATTER|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00037700322286|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.605588|80.605617967200075|99|1
35.43259|75198c0dfae66830d4fb64c71560b2b43c26808e|1.17|2014-12-19 16:00:00|80.606823361882718|2|7203690021|202|35.50077063756757|0|57|1033|-80.875654|163|35.585842|HAMBURGER|0.0|7|H T HAMBURGER BUNS|43166d9b1bc69df7e60a9afb900e55c512d04a79|4.711117707427967|35.500309569604553|00072036900210|BUNS/ROLLS|COMMERCIAL BAKERY|-80.605588|80.605617967200075|99|1
35.17739|99ebc2457265c88f28be6cc6568970452986bacf|7.99|2015-02-25 17:52:00|80.801203185414451|1|3077109653|208|35.181623388901841|0|24|499|-80.861571|110|35.444615|MEATBALLS|1.0|19|ALFRESCO MEATBALL ITALIAN|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00030771096544|FROZEN CASE MEAT|CASE READY MEATS|-80.80146|80.801472966259681|340|1
35.17739|d478519c38a3ad4d731aaf172ac2528e0f7b09e4|1.79|2015-01-09 07:34:00|1.4094857484078087|1|2000011274|208|0.613961277758128|0|26|245|-80.80146|39|35.17739|VEGETABLES-CORE|0.79|1|GREEN GIANT CORN S SWT YEL/WH|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00020000112749|VEGETABLES-CAN/JAR|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|4a0ecb5aaa98cf3b834c4edcee267e284d069321|4.19|2014-10-12 18:00:00|1.4094857484078087|1|1800000159|208|0.613961277758128|0|26|328|-80.80146|54|35.17739|SWEET ROLLS-REFRIGERATED|0.0|3|GRANDS CINNAMON ROLLS|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00018000001590|DOUGH PRODUCTS|DAIRY|-80.80146|1.4102515174184975|208|1
35.17739|4b0f2f2070264ff442ad3d9e26b8a2fa45d90d37|1.8|2015-01-27 08:18:00|1.4094857484078087|1|4667500010|208|0.613961277758128|0|26|682|-80.80146|61|35.17739|KIDS|0.6|3|YOCRUNCH VANILLA WITH M&M'S|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00046675000792|YOGURT|DAIRY|-80.80146|1.4102515174184975|208|2
35.17739|49f2dbf3c2356d4f5f6662857ffd924ebd74beab|3.19|2014-11-16 17:00:00|1.4094857484078087|1|4667501350|208|0.613961277758128|0|26|682|-80.80146|61|35.17739|KIDS|0.0|3|YOCRUNCH STRAW/SPRINKLINS 4 PK|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00046675013365|YOGURT|DAIRY|-80.80146|1.4102515174184975|208|1
35.17739|512e499b1737ab2972084a3964195a3f893a1d81|7.98|2015-03-02 15:28:00|1.4094857484078087|1|4610000012|208|0.613961277758128|0|26|318|-80.80146|52|35.17739|SHREDDED/GRATED CHEESE|1.99|3|SARGENTO OTB TRAD 4 CHS MEX|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00046100011072|CHEESE|DAIRY|-80.80146|1.4102515174184975|208|2
35.17739|ccd96c12da9a39a9ef8e3ffacbde9ae4278bb5fd|1.8|2014-10-06 14:43:00|1.4094857484078087|1|4667500010|208|0.613961277758128|0|26|682|-80.80146|61|35.17739|KIDS|0.8|3|YOCRUNCH VANILLA WITH M&M'S|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00046675000792|YOGURT|DAIRY|-80.80146|1.4102515174184975|208|2
35.17739|6a88ad5a9c132d8be8c6c3cd83a0ca9bae7d2d5f|3.19|2014-11-25 08:37:00|1.4094857484078087|1|4667501350|208|0.613961277758128|0|26|682|-80.80146|61|35.17739|KIDS|0.0|3|YOCRUNCH STRAW/DOVE CHOC 4 PK|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00046675013310|YOGURT|DAIRY|-80.80146|1.4102515174184975|208|1
35.17739|3fbcccfbe3e74179cd0146528fb8af1775b76940|1.8|2014-12-11 09:08:00|80.801203185414451|1|4667500010|208|35.181623400933425|0|24|682|-80.78468|61|35.096737|KIDS|0.0|3|YOCRUNCH VANILLA WITH M&M'S|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00046675000792|YOGURT|DAIRY|-80.80146|80.801463954731219|30|2
35.17739|08af2d324136e99240d403716cd0db13e5644c79|2.85|2014-09-21 12:28:00|1.4094857484078087|1|4600028869|208|0.613961277758128|0|26|77|-80.80146|272|35.17739|HISP SAUCES/SEASONINGS|0.0|1|OEP SEASONING TACO MILD|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00046000288765|HISPANIC PREP. FOODS|G1 GROCERY|-80.80146|1.4102515174184975|208|3
35.17739|12a01aa83ea176cfc110458011d35fd12ad35ae4|1.8|2015-01-06 08:29:00|1.4094857484078087|1|4667500010|208|0.613961277758128|0|26|682|-80.80146|61|35.17739|KIDS|0.0|3|YOCRUNCH VANILLA WITH M&M'S|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00046675000792|YOGURT|DAIRY|-80.80146|1.4102515174184975|208|2
35.17739|eea8f7fa3ec81db9383625ed86f3c67bbfe78906|1.19|2014-09-23 17:06:00|1.4094857484078087|1|3940001747|208|0.613961277758128|0|26|242|-80.80146|39|35.17739|CANNED BEANS|0.19|1|BUSH BEAN BLACK|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00039400018803|VEGETABLES-CAN/JAR|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|fff4cf1f8766ee31b96f3777b07fe725caffb559|5.99|2014-12-19 21:19:00|1.4094857484078087|1|3993803438|208|0.613961277758128|0|26|7407|-80.80146|1600|35.17739|CHRISTMAS PARTY GOODS/DECOR|0.99|18|GLITZ BEV NAP GREEN FOIL|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00039938034399|SEASONAL MERCHANDISE|GM|-80.80146|1.4102515174184975|208|1
35.17739|fecc56efe9ee76670980d4e94fd05c7c0601d6bb|13.29|2014-12-05 17:50:00|80.801203185414451|1|3700013882|208|35.181623401886974|0|24|389|-80.825175|66|35.152722|NFS-LAUNDRY DETERGENTS|0.0|1|TIDE FREE & GENTLE 64 LD|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00037000138907|DETERGENTS|G1 GROCERY|-80.80146|80.801461885435899|160|1
35.17739|67a751c757e66eb0827a96c11e7d8fefe087de25|10.21|2014-12-05 21:56:00|1.4094857484078087|1||208|0.613961277758128|0|26|503|-80.80146|64|35.17739|FRESH GRAPES|0.0|4|GREEN GRAPES, SEEDLESS 12/16|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00204022000004|FRESH PRODUCE|PRODUCE|-80.80146|1.4102515174184975|208|1
35.17739|69cc747d77d93780277b47ace9bbaf7a5129c24b|12.38|2015-01-01 11:33:00|1.4094857484078087|1|20331300000|208|0.613961277758128|0|26|641|-80.80146|137|35.17739|PREMIUM PORK|0.0|2|PORK LOIN CHOPS BONE-IN CUSTOM|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00203314000005|PORK|MEAT|-80.80146|1.4102515174184975|208|1
35.17739|80b5e15d1300c4b20b263c619a7d771b7d153045|3.99|2014-09-10 18:04:00|80.801203185414451|1|64339250026|208|35.181623368345569|0|24|62|-80.895009|7|35.603432|SPECIALTY BAR/BOX CHOCOLATE|0.0|1|SCHARF BERG MILK ALMOND BAR|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00643392500774|CANDY|G1 GROCERY|-80.80146|80.801480703762195|274|1
35.17739|45c2e64d2c20de50b53b8aa850a0775310b0a627|13.98|2015-02-16 09:10:00|1.4094857484078087|1|82476000205|208|0.613961277758128|0|26|561|-80.80146|64|35.17739|FR PROD ORGANIC PRODUCE|0.0|4|ORG STRAWBERRIES 1 LB|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00769197404144|FRESH PRODUCE|PRODUCE|-80.80146|1.4102515174184975|208|2
35.17739|d62a40a5d6e312bd86c4b993b5478464bd3210dc|2.29|2014-12-30 16:49:00|80.801203185414451|1|7800023046|208|35.181623401886974|0|24|54|-80.825175|8|35.152722|DIET|1.29|23|CANADA DRY DT G/ALE 2 LITER|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00078000148466|CARBONATED BEVERAGES|BEVERAGE|-80.80146|80.801461885435899|160|1
35.17739|69dd5b0ca779ea2d0dea842a18996901768c0c29|4.85|2014-10-23 09:02:00|80.801203185414451|1|7790011553|208|35.181623400933425|0|24|361|-80.78468|105|35.096737|BREAKFAST SAUSAGE|0.0|19|JIMMY DEAN MILD SAUSAGE|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00077900115530|BREAKFAST SAUSAGE|CASE READY MEATS|-80.80146|80.801463954731219|30|1
35.17739|a126c39fde70951a1c958c1b83c48170868598a3|18.16|2014-09-15 18:00:00|1.4094857484078087|1|20242200000|208|0.613961277758128|0|26|299|-80.80146|49|35.17739|ANGUS BEEF|0.0|2|ANGUS BEEF SKIRT STEAK FAJITAS|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00202422000006|BEEF|MEAT|-80.80146|1.4102515174184975|208|2
35.17739|4783d16330955c1dd3fe73f552d7f8ecb4e35b22|7.99|2015-02-09 07:48:00|1.4094857484078087|1|2840000288|208|0.613961277758128|0|26|205|-80.80146|31|35.17739|REMAINING SNACKS|1.0|1|FRITOLAY CLASSIC 20 CTN|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00028400002882|SNACKS|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|8c98709da87d597b3878cc41e6d8fed033818776|7.99|2015-02-22 20:06:00|1.4094857484078087|1|2840000288|208|0.613961277758128|0|26|205|-80.80146|31|35.17739|REMAINING SNACKS|1.0|1|FRITOLAY CLASSIC 20 CTN|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00028400002882|SNACKS|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|b64f00d54ff9ab3efba41dfec283d18fda6259f2|8.07|2014-12-11 18:04:00|80.801203185414451|1|7008506010|208|35.181623368345569|0|24|1277|-80.895009|279|35.603432|FROZEN SNACKS|2.07|5|BAGEL BITES CHEESE/SAUS/PEP|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00070085060138|FROZEN SANDWICH AND SNACKS|FROZEN|-80.80146|80.801480703762195|274|3
35.17739|9d8ac9443c540e5d9063ea7081893e4c5828a432|4.69|2014-11-23 14:08:00|1.4094857484078087|1|2700042063|208|0.613961277758128|0|26|242|-80.80146|39|35.17739|CANNED BEANS|1.19|1|HUNTS CHILI KIT|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00027000420638|VEGETABLES-CAN/JAR|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|beb7dedc2fbb9fccde1ffe10568d36d8adfa9e91|0.85|2014-10-31 15:10:00|1.4094857484078087|1||208|0.613961277758128|0|26|524|-80.80146|64|35.17739|FRESH PROD FRESH ONIONS|0.0|4|COO YELLOW ONIONS, LRG|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00204665000003|FRESH PRODUCE|PRODUCE|-80.80146|1.4102515174184975|208|1
35.17739|9823af0293b5f071682693dabda2223b81ca3e19|3.99|2014-09-21 17:04:00|1.4094857484078087|1|7020050025|208|0.613961277758128|0|26|580|-80.80146|136|35.17739|OTHER MERCH DRESSINGS|0.0|4|MARZ CHUNKY BLUE CHEESE DRESS|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00070200500211|OTHER MERCHANDISE|PRODUCE|-80.80146|1.4102515174184975|208|1
35.17739|d0a1963c7f919f54ae98b9706f5429a3ec50769f|2.85|2014-11-09 17:11:00|80.801203185414451|1|7203604237|208|35.181623368345569|0|24|41|-80.895009|6|35.603432|BREAKFAST BARS|0.88|1|HT BAR CEREAL BLUEBERRY|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00072036042392|BREAKFAST FOODS|G1 GROCERY|-80.80146|80.801480703762195|274|1
35.17739|ba16486de706b98f9ce6da14f3153e69e43a85c8|3.99|2014-12-31 14:27:00|1.4094857484078087|1|7020050025|208|0.613961277758128|0|26|580|-80.80146|136|35.17739|OTHER MERCH DRESSINGS|0.0|4|MARZ CHUNKY BLUE CHEESE DRESS|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00070200500211|OTHER MERCHANDISE|PRODUCE|-80.80146|1.4102515174184975|208|1
35.17739|58b5115ca1a45abed0256ce365242634f80cb06d|3.99|2015-01-02 19:09:00|1.4094857484078087|1|7020050025|208|0.613961277758128|0|26|580|-80.80146|136|35.17739|OTHER MERCH DRESSINGS|0.0|4|MARZ CHUNKY BLUE CHEESE DRESS|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00070200500211|OTHER MERCHANDISE|PRODUCE|-80.80146|1.4102515174184975|208|1
35.17739|5c852b5873a564911a06da15eb07342628e9f25c|4.99|2014-11-03 16:47:00|1.4094857484078087|1|7447029089|208|0.613961277758128|0|26|6789|-80.80146|1568|35.17739|MAGAZINES QUARTERLY|0.0|18|BOURBON REVIEW|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00074470290896|MAGAZINES|GM|-80.80146|1.4102515174184975|208|1
35.17739|2fd36238308dae1a2c2200e59f15f0503658de31|1.99|2014-11-04 17:58:00|80.801203185414451|1|7962597178|208|35.181623368345569|0|24|3303|-80.895009|1025|35.603432|BATH ACCESSORIES|0.0|17|BODY BENEFITS LUX BATH SPONGE|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00079625971781|BATH PRODUCTS|HBC|-80.80146|80.801480703762195|274|1
35.17739|413125945451716f2f649ab5e3d3d0ffea4ad06c|2.99|2014-12-23 09:06:00|1.4094857484078087|1|7172000611|208|0.613961277758128|0|26|52|-80.80146|7|35.17739|PKG NON CHOC|0.0|1|TOOTSIE ROLL MIDGEES|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00071720006115|CANDY|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|0083ef2ac5bb5c3ad6c0b8f9d89f9b286902a61e|2.0|2014-11-27 11:43:00|1.4094857484078087|1|7203663118|208|0.613961277758128|0|26|1262|-80.80146|57|35.17739|HALF N HALF WHIPPING CREAM|0.0|3|HT HALF & HALF|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00072036632043|MILK|DAIRY|-80.80146|1.4102515174184975|208|1
35.17739|ec74d6b405ca9f5bac2ab1a0fdeb812b7c067590|3.99|2015-03-02 08:05:00|80.801203185414451|1|7203670342|208|35.181623401886974|0|24|443|-80.825175|76|35.152722|NFS-GARBAGE BAGS|0.0|1|YH KTCHN BAG HANDLE TIE|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00072036703422|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.80146|80.801461885435899|160|1
35.17739|222bb3a842ab35270a8eac6e8eb9f5b39404ccc9|4.98|2015-02-14 16:17:00|80.801203185414451|1|4150880012|208|35.181623368345569|0|24|30|-80.895009|4|35.603432|CARBONATED WATER|0.49|1|SAN PELLEGRINO 750ML|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00041508800129|BOTTLED WATER|G1 GROCERY|-80.80146|80.801480703762195|274|2
35.17739|1c6162a6c770f32d3b010ae3114a662ee51bf642|2.49|2015-02-01 12:39:00|1.4094857484078087|1||208|0.613961277758128|0|26|561|-80.80146|64|35.17739|FR PROD ORGANIC PRODUCE|0.0|4|ORG ICEBERG LETTUCE|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00294061000004|FRESH PRODUCE|PRODUCE|-80.80146|1.4102515174184975|208|1
35.17739|8b64f119f9cb92cc0befa05cae5e9a2619c23bbf|4.49|2015-01-07 19:08:00|80.801203185414451|1|74759930652|208|35.181623368345569|0|24|62|-80.895009|7|35.603432|SPECIALTY BAR/BOX CHOCOLATE|0.0|1|GHIRARDELLI SEASALT SOIREE|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00747599313059|CANDY|G1 GROCERY|-80.80146|80.801480703762195|274|1
35.17739|63e07456682d6bc39f360ee7315f9d7176afa08a|1.99|2014-09-20 14:24:00|80.801203185414451|1|7203648011|208|35.181623401019287|0|24|274|-80.824767|44|35.116751|ICE|0.0|5|HT BAGGED ICE 10LB (456)|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00000000004560|ICE|FROZEN|-80.80146|80.801463814662625|294|1
35.17739|c987551936e0751c12163a64054107a47225fd6a|9.99|2014-10-24 19:19:00|1.4094857484078087|1|3410057509|208|0.613961277758128|0|26|455|-80.80146|82|35.17739|DOMESTIC PREMIUM 12PK&>|0.0|16|MILLER LITE 12PK 12OZ BTL|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00034100575090|DOMESTIC BEER|BEER|-80.80146|1.4102515174184975|208|1
35.17739|8e2503571708e8da50a358541aaf92a9a0d6fea6|2.49|2014-09-28 16:17:00|1.4094857484078087|1|1410008550|208|0.613961277758128|0|26|89|-80.80146|12|35.17739|GRAHAM CRACKERS|0.0|1|PF GF SWEET GRAHAM COOK CREAM|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00014100098317|COOKIES|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|1aa7bdcdf6f9365c09204c525c784ca73e009842|4.7700000000000005|2015-03-04 19:38:00|80.801203185414451|1|18473900016|208|35.181623368345569|0|24|31|-80.895009|4|35.603432|NON CARBONATED WATER|1.77|1|HINT BLACKBERRY ESS WATER|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00184739000309|BOTTLED WATER|G1 GROCERY|-80.80146|80.801480703762195|274|3
35.17739|4549d337d80f3a56e35b17a4ee788c2af078da86|3.18|2015-02-27 16:10:00|1.4094857484078087|1|18473900016|208|0.613961277758128|0|26|31|-80.80146|4|35.17739|NON CARBONATED WATER|0.0|1|HINT BLACKBERRY ESS WATER|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00184739000309|BOTTLED WATER|G1 GROCERY|-80.80146|1.4102515174184975|208|2
35.17739|b051542c597f53953dcfbd78988ab0b7ac86b3c3|3.18|2015-02-14 13:29:00|80.801203185414451|1|18473900016|208|35.181623402155267|0|24|31|-80.826724|4|35.195689|NON CARBONATED WATER|0.0|1|HINT BLACKBERRY ESS WATER|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00184739000309|BOTTLED WATER|G1 GROCERY|-80.80146|80.801460393259035|412|2
35.17739|d9ea6fc3dfa8728dd878716ea9a33113e2b6d48c|3.18|2015-02-10 20:21:00|1.4094857484078087|1|7684020027|208|0.613961277758128|0|26|275|-80.80146|45|35.17739|SUPER PREMIUM ICE CREAM|0.0|5|BEN & JERRY COOKIE DOUGH INDV|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00076840200276|ICE CREAM|FROZEN|-80.80146|1.4102515174184975|208|2
35.17739|8639cc2d4b346ab8e3e485e558152aa00fdc9021|5.99|2015-02-20 18:41:00|1.4094857484078087|1|7336108798|208|0.613961277758128|0|26|6787|-80.80146|1568|35.17739|MAGAZINES MONTHLY|0.0|18|CLEAN EATING|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00073361087980|MAGAZINES|GM|-80.80146|1.4102515174184975|208|1
35.17739|bfbe55903b72385291ceb248a20c1290f38c4628|3.99|2014-11-10 07:32:00|1.4094857484078087|1|8390000649|208|0.613961277758128|0|26|365|-80.80146|56|35.17739|REFRIGERATED TEAS|0.0|3|GOLD PEAK SWEET BLACK TEA|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00083900006495|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.80146|1.4102515174184975|208|1
35.17739|06d942c359f114a9bc7511c7ca7097ff2a668e5d|1.2|2015-01-22 14:21:00|80.801203185414451|1|7047000100|208|35.181623402155267|0|24|687|-80.826724|61|35.195689|BLENDED|0.0|3|YOPLAIT STRAWBERRY YOGURT|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00070470003009|YOGURT|DAIRY|-80.80146|80.801460393259035|412|2
35.17739|4e1bd3fc6cd5e4bc0dc263551223587ee6ab812c|1.39|2015-02-11 20:03:00|1.4094857484078087|1|1330054701|208|0.613961277758128|0|26|11|-80.80146|2|35.17739|MUFFIN MIXES|0.39|1|M WHITE BANANA NUT MUFFIN|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00013300579022|BAKING MIXES|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|84b999db72cd6ffbdcdfe65df5a7cdc557c99755|6.27|2015-02-08 15:58:00|1.4094857484078087|1|7203676359|208|0.613961277758128|0|26|345|-80.80146|57|35.17739|ORGANIC MILK|0.0|3|HTO ORGANIC 2% MILK GAL|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00072036763600|MILK|DAIRY|-80.80146|1.4102515174184975|208|1
35.17739|44939fe6fd58f168a00a52c13edd6ffb4eee9775|1.29|2015-01-16 12:26:00|1.4094857484078087|1|8379152001|208|0.613961277758128|0|26|1981|-80.80146|480|35.17739|CHIPS|0.0|6|DIRTY POTATO CHIP BBQ|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00083791520049|DRY GOODS|DELI|-80.80146|1.4102515174184975|208|1
35.17739|591de04e465543d26692448097c0bb25b4a6550e|2.58|2014-12-15 14:36:00|1.4094857484078087|1|8379152001|208|0.613961277758128|0|26|1981|-80.80146|480|35.17739|CHIPS|0.0|6|DIRTY POTATO CHIP BBQ|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00083791520049|DRY GOODS|DELI|-80.80146|1.4102515174184975|208|2
35.17739|58ff312688d59b04feb50feba3a4bcb55acd4d85|5.38|2014-11-19 18:19:00|80.801203185414451|1|73434100030|208|35.181623368345569|0|24|31|-80.895009|4|35.603432|NON CARBONATED WATER|0.4|1|LE BLEU ULT PURE CLR WATER 6PK|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00734341000305|BOTTLED WATER|G1 GROCERY|-80.80146|80.801480703762195|274|2
35.17739|793f7f5870ac1ac157cf11aa46f35c8e195bca24|3.29|2014-11-09 17:22:00|80.801203185414451|1|1410008786|208|35.181623402155267|0|24|1033|-80.826724|163|35.195689|HAMBURGER|0.0|7|PEP GOLDEN POTATO HAMS PP|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00014100091417|BUNS/ROLLS|COMMERCIAL BAKERY|-80.80146|80.801460393259035|412|1
35.17739|c085c0b84d2f0c8ef0f6b8ba956601366d733634|4.99|2014-11-12 17:54:00|80.801203185414451|1|88852610227|208|35.181623368345569|0|24|6785|-80.895009|1568|35.603432|MAGAZINES WEEKLY|0.0|18|PEOPLE|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00888526102275|MAGAZINES|GM|-80.80146|80.801480703762195|274|1
35.17739|e49e78a9161acfa37f4418ce5c63e8dab56ed42b|7.49|2015-02-09 15:10:00|1.4094857484078087|1|3770032228|208|0.613961277758128|0|26|423|-80.80146|72|35.17739|NFS-DISPOSE PLATES/BOWLS|0.0|1|CHINET DINNER PLATE 10 3/8IN|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00037700322262|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|db4e53be58fd1941dafb7af3abfb653e7f8f87cf|9.870000000000001|2014-10-17 14:46:00|80.801203185414451|1|1410008786|208|35.18162340182883|0|24|1035|-80.810056|163|35.219587|SANDWICH ROLL|0.0|7|PEP SLIDER BUNS  PP|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00014100093404|BUNS/ROLLS|COMMERCIAL BAKERY|-80.80146|80.801462071682707|401|3
35.17739|4909c8be2f52e1485d89ded0cae7ff5f308b2028|25.98|2015-01-16 12:29:00|1.4094857484078087|1|7203695587|208|0.613961277758128|0|26|1707|-80.80146|387|35.17739|MESSAGE|6.0|14|12 INCH MESSAGE COOKIE|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00072036955876|COOKIES|BAKERY|-80.80146|1.4102515174184975|208|2
35.17739|d6099e5c4a41608ac434c064f38c60f2b8de9d2d|5.99|2014-12-04 19:08:00|1.4094857484078087|1|89477300101|208|0.613961277758128|0|26|55|-80.80146|8|35.17739|REGULAR|0.0|23|ZEVIA GINGER ALE|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00894773001117|CARBONATED BEVERAGES|BEVERAGE|-80.80146|1.4102515174184975|208|1
35.17739|244bfdf8b1eaef443c2393683f10375bd82d8d6d|2.99|2014-10-15 15:31:00|1.4094857484078087|1|1600040175|208|0.613961277758128|0|26|15|-80.80146|2|35.17739|REMAINING BAKING MIXES|0.0|1|BC HRSHY CHOC CHUNK COOKIE MIX|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00016000401761|BAKING MIXES|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|1985fdf9fa0d3faa680f0d15de6bd8c713cbf839|10.99|2014-12-18 07:37:00|1.4094857484078087|1|74759931930|208|0.613961277758128|0|26|727|-80.80146|7|35.17739|SEASONAL CANDY-SINGLE FAC|1.5|1|I/O(C14)GHIR XL PEPP BARK|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00747599319303|CANDY|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|a9ef77d01acebe152a8cc558d1c48af92453acb0|13.47|2015-02-11 13:00:00|1.4094857484078087|1|70897191772|208|0.613961277758128|0|26|1703|-80.80146|387|35.17739|SEASONAL COOKIES|4.5|14|VALENTINE PINK FRSTD SGR COOK|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00708971917722|COOKIES|BAKERY|-80.80146|1.4102515174184975|208|3
35.17739|910391380fd4cfdc87410c34f67e1c94932683f0|6.99|2014-10-25 15:23:00|80.801203185414451|1|7480802477|208|35.181623400506673|0|24|6788|-80.85753|1568|35.116638|MAGAZINES BI-MONTHLY|0.0|18|SMARTPHONE & PCKT|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00074808024773|MAGAZINES|GM|-80.80146|80.801464587856344|204|1
35.17739|e1a1ab46f09bad006ef3447be02f1a061410bb7c|3.99|2014-12-24 09:18:00|80.801203185414451|1|7203676038|208|35.181623402155267|0|24|160|-80.826724|25|35.195689|OLIVES|0.99|1|HT TRADER OLIVES KALAMATA PTD|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00072036760364|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.80146|80.801460393259035|412|1
35.17739|fd1885664fc8873b2dc08b00b6c267e63a889113|11.97|2014-09-19 12:40:00|80.801203185414451|1|7203697777|208|35.181623369917077|0|24|31|-80.875654|4|35.585842|NON CARBONATED WATER|3.16|1|(U) HT PURIFIED WATER 24 PK|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00072036977779|BOTTLED WATER|G1 GROCERY|-80.80146|80.801480217051378|99|3
35.17739|9f134a6bb57cb36497fc17d8836c4f9391533a8f|11.97|2014-09-19 12:40:00|80.801203185414451|1|7203697777|208|35.181623369917077|0|24|31|-80.875654|4|35.585842|NON CARBONATED WATER|3.1599999999999997|1|(U) HT PURIFIED WATER 24 PK|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00072036977779|BOTTLED WATER|G1 GROCERY|-80.80146|80.801480217051378|99|3
35.17739|7e22bda679994ad3179065abb0624e3072e7a50c|15.96|2014-09-19 12:42:00|80.801203185414451|1|7203697777|208|35.181623369917077|0|24|31|-80.875654|4|35.585842|NON CARBONATED WATER|4.65|1|(U) HT PURIFIED WATER 24 PK|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00072036977779|BOTTLED WATER|G1 GROCERY|-80.80146|80.801480217051378|99|4
35.17739|4ff0a74e38a45b929ad3aa0ae5ed16b7d0c5d485|2.99|2015-02-13 17:46:00|80.801203185414451|1|7203698611|208|35.181623401886974|0|24|55|-80.825175|8|35.152722|REGULAR|0.0|23|HT CLUB SODA 6PK GLASS|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00072036986139|CARBONATED BEVERAGES|BEVERAGE|-80.80146|80.801461885435899|160|1
35.17739|584776fcfe32e1e049872e596b7a9e85219947ff|11.97|2014-09-19 12:41:00|80.801203185414451|1|7203697777|208|35.181623369917077|0|24|31|-80.875654|4|35.585842|NON CARBONATED WATER|3.16|1|(U) HT PURIFIED WATER 24 PK|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00072036977779|BOTTLED WATER|G1 GROCERY|-80.80146|80.801480217051378|99|3
35.17739|521bb40231cbdf3533a888fae953b77af26baecf|11.97|2014-09-19 12:41:00|80.801203185414451|1|7203697777|208|35.181623369917077|0|24|31|-80.875654|4|35.585842|NON CARBONATED WATER|3.16|1|(U) HT PURIFIED WATER 24 PK|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00072036977779|BOTTLED WATER|G1 GROCERY|-80.80146|80.801480217051378|99|3
35.17739|c0b0cf6a9ae6fed96e56dfde91477fe063e03bdc|5.39|2014-11-26 08:02:00|80.801203185414451|1|3450015193|208|35.181623401886974|0|24|312|-80.825175|51|35.152722|BUTTER|0.0|3|LOL BUTTER HALF STICKS|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00034500151818|BUTTER & MARGARINE|DAIRY|-80.80146|80.801461885435899|160|1
35.17739|9ce120b05b526907a22bc7e831b750c94861f93d|16.15|2014-10-07 10:45:00|80.801203185414451|1|31254720436|208|35.181623402155267|0|24|4189|-80.826724|1200|35.195689|ALLERGY REMEDY-CHILDREN|0.0|17|ZYRTEC CHILDREN DISSOLVE TABS|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00300450242259|COUGH/COLD/SINUS|HBC|-80.80146|80.801460393259035|412|1
35.17739|7bdf2ea9d1f6da751e96cb00ed0c8073678619f8|2.47|2015-03-09 19:23:00|80.801203185414451|1||208|35.181623400933425|0|24|561|-80.78468|64|35.096737|FR PROD ORGANIC PRODUCE|0.28|4|ORG BANANAS|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00294011000009|FRESH PRODUCE|PRODUCE|-80.80146|80.801463954731219|30|1
35.17739|23601f9711c57b75d14f9c6de586b0996cde21aa|1.0|2014-11-22 12:11:00|80.801203185414451|1|3400000031|208|35.181623401019287|0|24|47|-80.824767|7|35.116751|REGISTER BARS|0.25|1|YORK PEPPERMINT PATTIES|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|35.194272495053255|00034000003303|CANDY|G1 GROCERY|-80.80146|80.801463814662625|294|1
35.17739|91b728a4aee2d1b31f9922399bf423e6741c24a3|18.99|2014-09-29 16:39:00|1.4094857484078087|1|20941200000|208|0.613961277758128|0|26|672|-80.80146|147|35.17739|SCALLOPS|2.0|12|WC FRESH SEA SCALLOPS  (US)|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00209412000008|MOLLUSK|SEAFOOD|-80.80146|1.4102515174184975|208|1
35.17739|a58631dbdb2f9c337fd808e1c2adef7add45c13c|3.0|2015-02-17 18:16:00|1.4094857484078087|1|7457008202|208|0.613961277758128|0|26|275|-80.80146|45|35.17739|SUPER PREMIUM ICE CREAM|0.5|5|HAAGEN DAZ VANILLA CUP|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00074570082025|ICE CREAM|FROZEN|-80.80146|1.4102515174184975|208|2
35.17739|22a79b7ee9f44e4e81e1409d6af809078bd64b30|1.79|2015-03-01 15:32:00|1.4094857484078087|1||208|0.613961277758128|0|26|561|-80.80146|64|35.17739|FR PROD ORGANIC PRODUCE|0.0|4|ORG GREEN BELL PEPPERS|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00294065000000|FRESH PRODUCE|PRODUCE|-80.80146|1.4102515174184975|208|1
35.17739|7131a444f148d6a8396969704c4b78d4459b0a68|1.49|2014-12-24 16:17:00|1.4094857484078087|1|7203653022|208|0.613961277758128|0|26|1273|-80.80146|50|35.17739|BAG VEG NON STEAM|0.0|5|HT WHITE SHOEPEG CORN|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00072036530288|VEGETABLES-FROZEN|FROZEN|-80.80146|1.4102515174184975|208|1
35.17739|7967a2e0b3569f54a14b1c6f5d5b93a87aecd4e6|1.98|2014-12-12 14:00:00|1.4094857484078087|1|2880000057|208|0.613961277758128|0|26|242|-80.80146|39|35.17739|CANNED BEANS|0.0|1|HANOVER EZO CHICK PEAS|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00028800000570|VEGETABLES-CAN/JAR|G1 GROCERY|-80.80146|1.4102515174184975|208|2
35.17739|b6bed27017c53f8023e4f6e58364ab63200d6161|2.49|2014-09-21 12:34:00|1.4094857484078087|1|5040073942|208|0.613961277758128|0|26|1033|-80.80146|163|35.17739|HAMBURGER|0.2|7|BALL PARK WHITE HAMS 8PK PP|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00050400739420|BUNS/ROLLS|COMMERCIAL BAKERY|-80.80146|1.4102515174184975|208|1
35.17739|cbb86660f6e05eb2ee357e421e3b9c4100816b92|10.99|2015-02-02 16:18:00|1.4094857484078087|1|5210000467|208|0.613961277758128|0|26|217|-80.80146|34|35.17739|EXTRACTS FOOD COLORING|0.0|1|MC GOURMET ORG PURE VAN.EXTRAT|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00052100004679|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|7bc9e5b983e3b67d58209830de100f508f9a0963|4.99|2015-01-16 12:23:00|1.4094857484078087|1|3680013440|208|0.613961277758128|0|26|4235|-80.80146|1200|35.17739|PSE SOLID SINGLE INDGREDIENT|0.0|17|(PP) PSE TC M/S NASAL DEC TAB|43bf72ec0995d99287bf4a31b3c69e68ebe31909|0.2925178664717518|0.61471665291522548|00036800134409|COUGH/COLD/SINUS|HBC|-80.80146|1.4102515174184975|208|1
35.140781|609fc43865ddd11cec6a2729cc284a43896f6fad|2.99|2015-02-21 14:43:00|80.632521683083056|4|85598300265|39|35.184527846975918|0|39|583|-80.70901|136|35.17335|NUTS|0.0|4|CREATIVE SNACK WASABI PEAS|444071edb93ae1ec5d33aa15e4d8b507e2a89f06|3.0228014849361657|35.177497916598789|00855983002653|OTHER MERCHANDISE|PRODUCE|-80.62331|80.623312666567841|174|1
35.140781|29ef2f1c742f65250436119c429e173d016e1faa|2.99|2014-09-14 14:08:00|80.632521683083056|4|85598300265|39|35.184527846464213|0|39|583|-80.661096|136|35.172688|NUTS|0.0|4|CREATIVE SNACK WASABI PEAS|444071edb93ae1ec5d33aa15e4d8b507e2a89f06|3.0228014849361657|35.177497916598789|00855983002653|OTHER MERCHANDISE|PRODUCE|-80.62331|80.623318608100064|474|1
35.140781|8ee4ccae79b8386a4c047329f276cf4f258cb852|8.98|2014-12-18 16:01:00|80.632521683083056|4|4470003050|39|35.184527846464213|0|39|840|-80.661096|102|35.172688|TUBS|2.24|19|OM DELI FRESH ROTISSERE CHCKEN|444071edb93ae1ec5d33aa15e4d8b507e2a89f06|3.0228014849361657|35.177497916598789|00044700030998|LUNCHMEATS|CASE READY MEATS|-80.62331|80.623318608100064|474|2
35.140781|591f553035b8a1110112625950b59f0092a99065|4.79|2014-10-12 12:08:00|80.632521683083056|4|4470003050|39|35.184527846464213|0|39|840|-80.661096|102|35.172688|TUBS|1.79|19|OM DELI FRESH BLACK FOREST HAM|444071edb93ae1ec5d33aa15e4d8b507e2a89f06|3.0228014849361657|35.177497916598789|00044700032527|LUNCHMEATS|CASE READY MEATS|-80.62331|80.623318608100064|474|1
35.140781|8dad8c8b1b3df5cb53eb89f74a5d8d9dd03161c2|6.98|2014-11-30 11:11:00|80.632521683083056|4|4812127620|39|35.184527846464213|0|39|1037|-80.661096|164|35.172688|ENGLISH MUFFINS|1.74|7|THOMAS 100% WHEAT ENG MUFN PP|444071edb93ae1ec5d33aa15e4d8b507e2a89f06|3.0228014849361657|35.177497916598789|00048121184070|BREAKFAST|COMMERCIAL BAKERY|-80.62331|80.623318608100064|474|2
35.140781|c5ae5dbe198a946a6b2b20de6231b3583d1c9609|3.01|2015-02-22 13:10:00|80.632521683083056|4|20037600000|39|35.184527846464213|0|39|1801|-80.661096|400|35.172688|FFM TURKEY|0.0|6|TURKEY BREAST|444071edb93ae1ec5d33aa15e4d8b507e2a89f06|3.0228014849361657|35.177497916598789|00200376000004|FFM MEAT|DELI|-80.62331|80.623318608100064|474|1
35.140781|1ea33e14b26bee706f6cd5571265edb2e40d53ca|12.450000000000001|2014-12-07 14:30:00|80.632521683083056|4|4369505631|39|35.184527846464213|0|39|1276|-80.661096|279|35.172688|FROZEN SANDWICHES|2.45|5|LEAN POCKETS BACON, EGG & CHS|444071edb93ae1ec5d33aa15e4d8b507e2a89f06|3.0228014849361657|35.177497916598789|00043695062502|FROZEN SANDWICH AND SNACKS|FROZEN|-80.62331|80.623318608100064|474|5
35.140781|f7ebd37b92944812ecb30d02fa4075c03c45a135|9.99|2015-01-04 13:27:00|80.632521683083056|4|3410057636|39|35.184527846464213|0|39|455|-80.661096|82|35.172688|DOMESTIC PREMIUM 12PK&>|0.0|16|MILLER LITE 12PK CAN|444071edb93ae1ec5d33aa15e4d8b507e2a89f06|3.0228014849361657|35.177497916598789|00034100576363|DOMESTIC BEER|BEER|-80.62331|80.623318608100064|474|1
35.140781|1820a2a4bf767ca061b42db427b00ed6e5905d5a|8.63|2014-10-08 17:08:00|80.632521683083056|4|20701800000|39|35.184527846464213|0|39|1935|-80.661096|465|35.172688|CHEF CASE|2.16|6|FRUIT & NUT CHICKEN SALAD|444071edb93ae1ec5d33aa15e4d8b507e2a89f06|3.0228014849361657|35.177497916598789|00207018000002|COLD PREPARED FOODS|DELI|-80.62331|80.623318608100064|474|1
35.43259|22b571d94c01c826816bf935d8e1ed618eac0e1d|2.49|2014-09-27 11:02:00|80.607132136635443|2|7156766109|202|35.477427483181714|0|9|52|-80.770346|7|35.052812|PKG NON CHOC|0.0|1|JBELLY SOURS|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00071567950589|CANDY|G1 GROCERY|-80.605588|80.605846872738738|40|1
35.43259|a8ef9f6cdfa34dd86a28799942689419b2b66971|3.79|2014-09-28 01:44:00|1.4057311447477159|2|7020055600|202|0.6184153580092175|0|52|582|-80.605588|136|35.43259|DIPS-REFRIG. & DRY|0.0|4|MARZ CARAMEL APPLE DIP|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|0.6209993146566879|00070200556003|OTHER MERCHANDISE|PRODUCE|-80.605588|1.406832906106031|202|1
35.43259|c2afa293282956a0e4dbc275bda3c2ec620f9674|23.96|2015-01-03 16:57:00|80.607132136635443|2|74759931696|202|35.477427483181714|0|9|727|-80.770346|7|35.052812|SEASONAL CANDY-SINGLE FAC|2.99|1|I/O(C14)GHIR IMPRESSIONS SUB|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00747599316968|CANDY|G1 GROCERY|-80.605588|80.605846872738738|40|4
35.43259|b2292006635020beb7d6d35f46a1c85cf746283b|3.39|2014-10-26 13:36:00|80.607132136635443|2|3700007100|202|35.477427483181714|0|9|393|-80.770346|68|35.052812|NFS-AIR FRESHENERS|0.4|1|FEBREZE AIR AFFECT GREEK SEASD|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00037000905981|FRESHENERS/DEODORIZERS|G1 GROCERY|-80.605588|80.605846872738738|40|1
35.43259|e2649e8cf5c1dc28f6b3c0b4c2457b704d43a550|19.99|2015-01-30 19:17:00|80.607132136635443|2|1780013476|202|35.477427412135583|0|9|156|-80.8062|24|35.037115|NFS-DOG FOOD-DRY|5.0|1|BENEFUL HEALTHY FIESTA|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00017800141970|PET FOOD/SUPPLIES|G1 GROCERY|-80.605588|80.605864797593071|27|1
35.43259|2b26bb2d89e9880bbf18b4c2afe07123deb558c4|1.29|2015-01-26 13:06:00|80.607132136635443|2|2100002322|202|35.477427483181714|0|9|714|-80.770346|274|35.052812|MICROWAVE MEALS|0.29|1|VELVEETA CUP ORIGINAL|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00021000023226|PREP FOODS DINNERS|G1 GROCERY|-80.605588|80.605846872738738|40|1
35.43259|136091527d8d34625b40402f03fa03f23e15e0f9|19.99|2015-03-09 17:43:00|80.607132136635443|2|1780013476|202|35.477427483181714|0|9|156|-80.770346|24|35.052812|NFS-DOG FOOD-DRY|4.51|1|BENEFUL HEALTHY FIESTA|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00017800141970|PET FOOD/SUPPLIES|G1 GROCERY|-80.605588|80.605846872738738|40|1
35.43259|30651502f80ae8ef86cd3c1390f053518705198b|1.29|2015-02-16 14:12:00|80.607132136635443|2|2100002322|202|35.477427483181714|0|9|714|-80.770346|274|35.052812|MICROWAVE MEALS|0.0|1|VELVEETA CUP ORIGINAL|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00021000023226|PREP FOODS DINNERS|G1 GROCERY|-80.605588|80.605846872738738|40|1
35.43259|2357fd537930d503fe89678d9749215410a0d045|19.99|2015-01-04 12:26:00|80.607132136635443|2|1780013476|202|35.477427483181714|0|9|156|-80.770346|24|35.052812|NFS-DOG FOOD-DRY|4.51|1|BENEFUL HEALTHY FIESTA|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00017800141970|PET FOOD/SUPPLIES|G1 GROCERY|-80.605588|80.605846872738738|40|1
35.43259|5a5ae44ec2b478cbfd5d06c69d0b9007808ef695|19.99|2014-12-16 19:26:00|80.607132136635443|2|1780013476|202|35.477427483181714|0|9|156|-80.770346|24|35.052812|NFS-DOG FOOD-DRY|4.51|1|BENEFUL HEALTHY FIESTA|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00017800141970|PET FOOD/SUPPLIES|G1 GROCERY|-80.605588|80.605846872738738|40|1
35.43259|5235e5641dddbd31b514b04540b9dde4b05fe685|2.29|2014-09-25 12:55:00|80.607132136635443|2|4132100541|202|35.477427483181714|0|9|184|-80.770346|28|35.052812|SALAD DRESSINGS-LIQUID|0.0|1|D WISHBONE DRS FF VIN ITALIAN|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00041000005411|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.605588|80.605846872738738|40|1
35.43259|8213681055cfb9a5a072087d33cb6ba45d2a16ab|1.89|2014-10-19 17:33:00|80.607132136635443|2|4000000432|202|35.477427412135583|0|9|47|-80.8062|7|35.037115|REGISTER BARS|0.0|1|E  SNICKERS KING SIZE BAR|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00040000002635|CANDY|G1 GROCERY|-80.605588|80.605864797593071|27|1
35.43259|4c3dc0637e33acc3ff3ce4861518baa4e974876d|21.99|2015-01-08 14:42:00|80.607132136635443|2|8985402092|202|35.477427483181714|0|9|9972|-80.770346|888|35.052812|NFS-U/PREM-CAB SAUVIGNON|0.0|13|WILDHORSE CABERNET|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00089854020921|ULTRA PREMIUM ($15-$19.99)|WINE|-80.605588|80.605846872738738|40|1
35.43259|53b8b76794f3e02d0dbd07c5cd5e132ac1aa9613|0.79|2014-11-16 16:05:00|80.607132136635443|2||202|35.477427412135583|0|9|532|-80.8062|64|35.037115|FRESH CUCUMBERS|0.0|4|COO CUCUMBERS S/S|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00204062000002|FRESH PRODUCE|PRODUCE|-80.605588|80.605864797593071|27|1
35.43259|36b555acb81dd62fc98f428b004673b19847fec5|9.99|2014-11-17 20:35:00|80.607132136635443|2|61262020112|202|35.477427483181714|0|9|458|-80.770346|82|35.052812|CRAFT BEER|0.0|16|FOOTHILLS HOPPYUM IPA 6PK|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00612620201127|DOMESTIC BEER|BEER|-80.605588|80.605846872738738|40|1
35.43259|0bb6c8f4a95105031db977d8cbff7d5a1a50e094|1.38|2014-09-24 14:16:00|80.607132136635443|2|71070842249|202|35.477427412135583|0|9|580|-80.8062|136|35.037115|OTHER MERCH DRESSINGS|0.0|4|ORGANIC FF ITALIAN DRESSING|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00710708422492|OTHER MERCHANDISE|PRODUCE|-80.605588|80.605864797593071|27|2
35.43259|f712643a5655b159eb69bcf984d612cf4551e9f5|5.97|2015-01-25 15:16:00|80.607132136635443|2|7203688096|202|35.477427483181714|0|9|526|-80.770346|64|35.052812|FRESH MUSHROOMS|0.0|4|HT SLICED WHITE MUSHROOMS|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00072036880963|FRESH PRODUCE|PRODUCE|-80.605588|80.605846872738738|40|3
35.43259|46fb93df68051c55420e637ccb9af73e41dcddb2|9.99|2014-11-03 21:01:00|80.607132136635443|2|8500000843|202|35.477427483181714|0|9|9951|-80.770346|886|35.052812|NFS-PREM-PINOT GRIS/GRIG|0.0|13|CB-ECCO DOMANI PINOT GRIGIO|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00085000008430|PREMIUM ($8-$10.99)|WINE|-80.605588|80.605846872738738|40|1
35.43259|6078b976510d69cea7367982967f06db594b2d8a|10.99|2014-12-29 20:49:00|80.607132136635443|2|8600387388|202|35.477427483181714|0|9|9934|-80.770346|885|35.052812|NFS POP CHARDONNAY|0.0|13|CB-WOODBRIDGE CHARDONNAY 1.5L|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00086003873889|POPULAR (4-$7.99)|WINE|-80.605588|80.605846872738738|40|1
35.43259|b6c63b812e157543589407cbdce674822d6c84dc|4.97|2015-03-08 10:46:00|80.607132136635443|2|7229000227|202|35.477427483181714|0|9|1271|-80.770346|41|35.052812|PROTEIN BREAKFAST|0.0|5|TENN PRIDE CHKN&BTTRMLK BISC|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00072290022406|BREAKFAST FOODS FROZEN|FROZEN|-80.605588|80.605846872738738|40|1
35.43259|7310e3e593ccba99bfabb7bfc82bad596a45502c|4.98|2014-09-20 10:42:00|80.607132136635443|2|7878350610|202|35.477427483181714|0|9|527|-80.770346|64|35.052812|FRESH CARROTS|0.0|4|MATCHSTICK CARROTS, PKG|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00078783506101|FRESH PRODUCE|PRODUCE|-80.605588|80.605846872738738|40|2
35.43259|749ecaa6af34300352b2191c9abaf8e26a80f39f|3.49|2015-03-03 16:15:00|80.607132136635443|2|7203670327|202|35.477427483181714|0|9|440|-80.770346|76|35.052812|NFS-ALUMINUM FOIL|0.0|1|YH ALUM FOIL HD 50 FT|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00072036703279|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.605588|80.605846872738738|40|1
35.43259|e6d0e70e070823a8508feb346cbc8de13410e1cb|1.99|2015-01-19 14:37:00|80.607132136635443|2|3600039408|202|35.477427483181714|0|9|426|-80.770346|72|35.052812|NFS-PAPER TOWELS|0.0|1|VIVA VANTAGE SINGLE ROLL 59CT|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00036000394085|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.605588|80.605846872738738|40|1
35.43259|2e5851f9b24e13d418977da9baf15365dd01a90f|8.99|2014-11-25 17:57:00|80.607132136635443|2|2484218211|202|35.477427412135583|0|9|1886|-80.8062|440|35.037115|FILLED PASTA|0.0|6|BUITONI SPINACH RICOTTA TORT|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00024842751319|PASTA|DELI|-80.605588|80.605864797593071|27|1
35.43259|576e72d11558165fdf85e464f25366b9af875932|8.99|2014-10-01 22:28:00|80.607132136635443|2|8130859207|202|35.477427483181714|0|9|9947|-80.770346|886|35.052812|NFS-PREM-CHARDONNAY|0.0|13|CB-CUPCAKE CHARDONNAY|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00081308592077|PREMIUM ($8-$10.99)|WINE|-80.605588|80.605846872738738|40|1
35.43259|ba3a10ab377a64f0f8aad4efd14cd08c09289ceb|8.99|2014-09-18 21:07:00|80.607132136635443|2|8130859207|202|35.477427483181714|0|9|9947|-80.770346|886|35.052812|NFS-PREM-CHARDONNAY|0.0|13|CB-CUPCAKE CHARDONNAY|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00081308592077|PREMIUM ($8-$10.99)|WINE|-80.605588|80.605846872738738|40|1
35.43259|359d945ace6ac30638b3be6ce54e74852e098a96|1.69|2014-10-07 21:01:00|80.607132136635443|2|4900000044|202|35.477427483181714|0|9|54|-80.770346|8|35.052812|DIET|0.0|23|CB COKE ZERO 20 OZ|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00049000040869|CARBONATED BEVERAGES|BEVERAGE|-80.605588|80.605846872738738|40|1
35.43259|8444666a24cc0b35bd4dc058b1b582154ea248a6|1.39|2014-10-12 15:30:00|80.607132136635443|2|1254661959|202|35.477427412135583|0|9|48|-80.8062|7|35.037115|REGISTER GUM|0.39|1|TRIDENT SUGARLESS GUM|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00012546612296|CANDY|G1 GROCERY|-80.605588|80.605864797593071|27|1
35.43259|0a7148f796ff7a96a563d825cee272a0497c2173|2.29|2015-01-31 10:54:00|80.607132136635443|2|4000040145|202|35.477427483181714|0|9|62|-80.770346|7|35.052812|SPECIALTY BAR/BOX CHOCOLATE|0.0|1|DOVE DARK CHOCOLATE BAR|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00040000401896|CANDY|G1 GROCERY|-80.605588|80.605846872738738|40|1
35.43259|bc0cb2a87d94e840349f8ed4ffda4632952139cb|1.99|2015-02-01 11:00:00|80.607132136635443|2|7203688083|202|35.477427483181714|0|9|526|-80.770346|64|35.052812|FRESH MUSHROOMS|0.2|4|HT WHITE MUSHROOMS, 8 OZ WHOLE|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00072036880833|FRESH PRODUCE|PRODUCE|-80.605588|80.605846872738738|40|1
35.43259|a58d78c2c6e6590387bc41aafa26a90b9dc986bf|2.29|2014-11-23 15:42:00|80.607132136635443|2|1200000649|202|35.477427483181714|0|9|854|-80.770346|32|35.052812|LIQUID ICED COFFEES|0.0|1|STARBUCK'S FRAPPUCCINO MOCHA|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00012000006494|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.605588|80.605846872738738|40|1
35.43259|293b54ef76e28cfd8aee6e7fb6f629e883fe624f|10.49|2014-11-05 10:10:00|80.607132136635443|2|9484130014|202|35.477427412135583|0|9|4922|-80.8062|1245|35.037115|EAR DROP-HOMEOPATHIC|0.0|17|SIMILASAN EAR RELIEF|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00094841255149|EYE & EAR CARE|HBC|-80.605588|80.605864797593071|27|1
35.43259|a6511a9470923a20ed12fdec2be92055f4ab019f|1.5|2014-10-03 10:41:00|80.607132136635443|2|3663203732|202|35.477427483181714|0|9|685|-80.770346|61|35.052812|GREEK|0.5|3|DANNON LNF GREEK PINEAPPLE|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00036632037343|YOGURT|DAIRY|-80.605588|80.605846872738738|40|1
35.43259|088e17e09203443e0e46c46c98991855804fa8b5|1.17|2014-11-03 21:54:00|80.607132136635443|2|7203669099|202|35.477427483181714|0|9|4834|-80.770346|1235|35.052812|COTTON/SWABS|0.0|17|HT PAPER STICK SWABS  -69099|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00072036690999|FIRST AID|HBC|-80.605588|80.605846872738738|40|1
35.43259|d53d9ce03fdf7e829c69f6175a243991979ffc14|1.79|2014-11-17 20:39:00|80.607132136635443|2|5200033875|202|35.477427483181714|0|9|171|-80.770346|20|35.052812|ISOTONIC DRINKS|0.9|1|GATORADE G2 FRUIT PUNCH|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00052000321982|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.605588|80.605846872738738|40|1
35.43259|6bc6734a5b47f3f293b9498b908c54bfa986ca3d|4.79|2015-01-10 22:17:00|80.607132136635443|2|7214001565|202|35.477427412135583|0|9|3204|-80.8062|1015|35.037115|ST LIP CARE|0.0|17|NIVEA LIP CARE & COLOR CORAL|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00072140015657|HAND & BODY LOTION/SUN CARE|HBC|-80.605588|80.605864797593071|27|1
35.43259|de0b6ccda718713b536019c673faa79fc35ef25a|2.77|2014-09-20 10:42:00|80.607132136635443|2||202|35.477427483181714|0|9|500|-80.770346|64|35.052812|FRESH APPLES|0.0|4|FUJI APPLES|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00204131000001|FRESH PRODUCE|PRODUCE|-80.605588|80.605846872738738|40|1
35.43259|a1044a35a97109bd0f73ba7b4511d11cf96df2f4|4.49|2015-01-31 10:53:00|80.607132136635443|2|7203670428|202|35.477427483181714|0|9|685|-80.770346|61|35.052812|GREEK|0.1|3|HT NF PLAIN GREEK YOGURT|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00072036704283|YOGURT|DAIRY|-80.605588|80.605846872738738|40|1
35.43259|06f7e16c1b2c50ec9a0eeca5b95b9cc3fac255f4|2.99|2014-11-25 18:01:00|80.607132136635443|2|3485602884|202|35.477427412135583|0|9|1200|-80.8062|6|35.037115|FRUIT SNACKS|0.0|1|WELCH'S FRUIT SNACKS MIX FRUIT|47709a3c6339d0069aa9b842fc910e8b478e2730|3.0981960717856984|35.47365851958088|00034856028888|BREAKFAST FOODS|G1 GROCERY|-80.605588|80.605864797593071|27|1
35.297134|d7dabd1d5fd0708afa5ebbbe377d81f0186f3829|6.99|2015-02-26 17:16:00|1.4094857484078087|4|7580587490|258|0.6160512048176361|0|26|2018|-80.737839|505|35.297134|PRESSED CHEESE|2.0|6|STELLA FONTINELLA WEDGE|49a8a26c8571553cd14258abc3ec67e8de18b8d7|2.002221782459263|0.61471665291522548|00075805874903|SPECIALTY CHEESE|DELI|-80.737839|1.409141121495086|258|1
35.297134|b91e61f1aae58b3c67cf61969e4bbb14388488d8|4.0|2014-12-04 17:40:00|1.4094857484078087|4||258|0.6160512048176361|0|26|511|-80.737839|64|35.297134|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|49a8a26c8571553cd14258abc3ec67e8de18b8d7|2.002221782459263|0.61471665291522548|00204770000004|FRESH PRODUCE|PRODUCE|-80.737839|1.409141121495086|258|2
35.297134|319fc32494987fbd293ef155863c8f5d093f0fb8|4.0|2015-01-22 16:59:00|1.4094857484078087|4||258|0.6160512048176361|0|26|511|-80.737839|64|35.297134|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|49a8a26c8571553cd14258abc3ec67e8de18b8d7|2.002221782459263|0.61471665291522548|00204770000004|FRESH PRODUCE|PRODUCE|-80.737839|1.409141121495086|258|2
35.297134|838e5d59328f4cd34d0b459d701e1bdeff82af23|3.05|2015-01-04 18:20:00|1.4094857484078087|4|20666000000|258|0.6160512048176361|0|26|2019|-80.737839|505|35.297134|PRESSED COOKED CHEESE|0.0|6|JARLSBERG WHEEL (FC)|49a8a26c8571553cd14258abc3ec67e8de18b8d7|2.002221782459263|0.61471665291522548|00206660000002|SPECIALTY CHEESE|DELI|-80.737839|1.409141121495086|258|1
35.323246|16352f9afd888b58221bdd249ff30312bbdf3385|1.99|2015-01-02 15:13:00|1.4102725052409182|4|68396988515|166|0.6165069451919168|0|1|8481|-80.945176|1769|35.323246|BATTERY-WATCH & CALC|0.0|18|AC DELCO CR 2032|4d6fe536dad8f9a55dba158da86a4d4bab11b814|1.3823929949234939|0.61833652052202714|00683969885156|BATTERY & FLASHLIGHT|GM|-80.945176|1.4127598348062935|166|1
35.323246|756c1dce464e31836427fa114a1dca79a69f50cf|4.99|2014-12-24 18:39:00|80.945255278477163|4|2840008313|166|35.343252384360525|0|13|204|-80.810056|31|35.219587|TORTILLA CHIPS|1.0|1|TOSTITOS RSTC FAMILY SIZE|4d6fe536dad8f9a55dba158da86a4d4bab11b814|1.3823929949234939|35.37387923947206|00028400083133|SNACKS|G1 GROCERY|-80.945176|80.945187397551479|401|1
35.323246|ecca3d60fbe39000b10948f57468adb1007acbb6|3.99|2014-11-07 18:37:00|1.4102725052409182|4|7203695676|166|0.6165069451919168|0|1|1656|-80.945176|381|35.323246|CUP CAKES|0.0|14|FFM MINI VANILLA CUPCAKES|4d6fe536dad8f9a55dba158da86a4d4bab11b814|1.3823929949234939|0.61833652052202714|00072036956767|CAKES|BAKERY|-80.945176|1.4127598348062935|166|1
35.323246|dcba6945e7d6e73584e8214330714d5694145173|7.98|2014-09-13 19:17:00|1.4102725052409182|4|7184509830|166|0.6165069451919168|0|1|207|-80.945176|32|35.323246|COCKTAIL MIXES|0.0|1|COCO LOPEZ CREAM OF COCONUT|4d6fe536dad8f9a55dba158da86a4d4bab11b814|1.3823929949234939|0.61833652052202714|00071845098309|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.945176|1.4127598348062935|166|2
35.323246|c1a92b35ac83fdfb4c0decf3adb016c3d159bba5|11.97|2014-11-15 16:29:00|1.4102725052409182|4|7184509830|166|0.6165069451919168|0|1|207|-80.945176|32|35.323246|COCKTAIL MIXES|1.2000000000000002|1|COCO LOPEZ CREAM OF COCONUT|4d6fe536dad8f9a55dba158da86a4d4bab11b814|1.3823929949234939|0.61833652052202714|00071845098309|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.945176|1.4127598348062935|166|3
35.323246|0c6b15c91b1d60e34e39f170d13bd84dc3557a66|11.07|2014-11-22 15:50:00|1.4102725052409182|4|2100062503|166|0.6165069451919168|0|1|318|-80.945176|52|35.323246|SHREDDED/GRATED CHEESE|1.84|3|KRAFT 2%  MILD CHEDDAR SHRED|4d6fe536dad8f9a55dba158da86a4d4bab11b814|1.3823929949234939|0.61833652052202714|00021000024667|CHEESE|DAIRY|-80.945176|1.4127598348062935|166|3
35.323246|b70b2fe8a74707daec222261ab5a975e6639b6fc|3.39|2014-11-15 16:28:00|1.4102725052409182|4|1312000286|166|0.6165069451919168|0|1|1469|-80.945176|278|35.323246|REGULAR CUT FRIES|1.7|5|ORE-IDA GOLDEN FRIES|4d6fe536dad8f9a55dba158da86a4d4bab11b814|1.3823929949234939|0.61833652052202714|00013120002588|FROZEN POTATO|FROZEN|-80.945176|1.4127598348062935|166|1
35.323246|2bbe4c645da4e0b867870d9957039a10f5ec21a0|2.99|2015-02-01 15:01:00|1.4102725052409182|4|7044650000|166|0.6165069451919168|0|1|498|-80.945176|111|35.323246|PICKLES & SAUERKRAUT|0.9|19|BOARS HEAD SAUERKRAUT 32 OZ|4d6fe536dad8f9a55dba158da86a4d4bab11b814|1.3823929949234939|0.61833652052202714|00070446500006|MISC. PACKAGED MEATS|CASE READY MEATS|-80.945176|1.4127598348062935|166|1
35.323246|b625c295379fffb32006947a5f9f008b39aeeefc|12.870000000000001|2015-02-24 13:33:00|1.4102725052409182|4|1380010067|166|0.6165069451919168|0|1|1279|-80.945176|48|35.323246|SINGLE SERVE FLAVOR|0.95|5|STOUFFER MACARONI & CHEESE|4d6fe536dad8f9a55dba158da86a4d4bab11b814|1.3823929949234939|0.61833652052202714|00013800103420|FROZEN MEALS|FROZEN|-80.945176|1.4127598348062935|166|3
35.323246|8a0b11bc2cbf0d2df4d19299db91dfab662703ad|6.0|2015-02-23 11:58:00|1.4102725052409182|4||166|0.6165069451919168|0|1|1617|-80.945176|373|35.323246|ROLLS BULK|0.0|14|BULK ROLLS|4d6fe536dad8f9a55dba158da86a4d4bab11b814|1.3823929949234939|0.61833652052202714|00072036955555|ROLLS|BAKERY|-80.945176|1.4127598348062935|166|8
35.323246|63b08301b34be818010069bfa2d5aefc58515152|2.25|2014-10-18 19:04:00|1.4102725052409182|4||166|0.6165069451919168|0|1|1617|-80.945176|373|35.323246|ROLLS BULK|0.0|14|BULK ROLLS|4d6fe536dad8f9a55dba158da86a4d4bab11b814|1.3823929949234939|0.61833652052202714|00072036955555|ROLLS|BAKERY|-80.945176|1.4127598348062935|166|3
35.323246|9127cb2d4f321369e0a7e1070131e87ac95e1e74|6.99|2015-02-24 13:34:00|1.4102725052409182|4|71921814141|166|0.6165069451919168|0|1|6204|-80.945176|1548|35.323246|HIGH END|0.0|18|PURAFILTER 2000 14/14/1|4d6fe536dad8f9a55dba158da86a4d4bab11b814|1.3823929949234939|0.61833652052202714|00719218141411|FURNACE FILTERS|GM|-80.945176|1.4127598348062935|166|1
35.323246|eed5596d328d79fb79a103ea5e7194b9335f2ccf|24.99|2015-02-13 20:49:00|1.4102725052409182|4|7203696866|166|0.6165069451919168|0|1|740|-80.945176|87|35.323246|NFS-ROSE BQT|5.0|9|15 STEM ROSE BOUQUET|4d6fe536dad8f9a55dba158da86a4d4bab11b814|1.3823929949234939|0.61833652052202714|00072036968661|FLORAL|FLORAL|-80.945176|1.4127598348062935|166|1
35.323246|16e7b092472e34b59fe2cc9899628ebcd895c3d7|3.59|2014-12-26 20:12:00|1.4102725052409182|4|7225002096|166|0.6165069451919168|0|1|1033|-80.945176|163|35.323246|HAMBURGER|0.6|7|CBC WHITE GRINDER SUB ROLL 6PK|4d6fe536dad8f9a55dba158da86a4d4bab11b814|1.3823929949234939|0.61833652052202714|00072250020961|BUNS/ROLLS|COMMERCIAL BAKERY|-80.945176|1.4127598348062935|166|1
35.297134|262aed0b8ebdf37569fefbbc1f539703aa876699|6.49|2015-02-06 18:52:00|80.737901233649083|4|7203676033|258|35.358252619956154|0|46|194|-80.844274|30|35.204336|OLIVE OIL|0.0|1|HT TRADER EV OLV OIL TRAD 17|506a6fdfb21d1e2beaeadfc6c26bf49646f91b72|4.2231534722856425|35.349871187060224|00072036760333|SHORTENING/OIL|G1 GROCERY|-80.737839|80.737947500836285|61|1
35.297134|0c18a0e8cf158507b860dca7adc43ec9153d85d4|2.65|2014-12-22 20:03:00|80.737901233649083|4|4119601000|258|35.35825257386837|0|46|1201|-80.825175|33|35.152722|RTS CANNED|1.33|1|PROG TRAD CHICKEN ROTINI|506a6fdfb21d1e2beaeadfc6c26bf49646f91b72|4.2231534722856425|35.349871187060224|00041196911169|SOUP|G1 GROCERY|-80.737839|80.737981253740671|160|1
35.297134|d684256369dccfcae6cfb989dc4a5160a3e65816|5.99|2015-01-22 20:12:00|80.737901233649083|4|79285001444|258|35.358252644719229|0|46|3272|-80.810056|1023|35.219587|NATURAL/ORGANIC PRODUCT|0.0|17|BURTS B TOWELETTES SENS|506a6fdfb21d1e2beaeadfc6c26bf49646f91b72|4.2231534722856425|35.349871187060224|00792850016774|NATURAL PERSONAL CARE|HBC|-80.737839|80.73792399921274|401|1
35.297134|de31b4d3ce80f7546aee4be93e4514f703e25d5e|4.49|2014-09-30 13:10:00|80.737901233649083|4|81857000790|258|35.35825257386837|0|46|725|-80.825175|66|35.152722|NFS-DISHWASHING LIQUID|0.7|1|WATKINS LIQ DISH LAVENDAR|506a6fdfb21d1e2beaeadfc6c26bf49646f91b72|4.2231534722856425|35.349871187060224|00818570007905|DETERGENTS|G1 GROCERY|-80.737839|80.737981253740671|160|1
35.297134|6e1d7d736b98435d4ffcc470c37889ec084c4eed|5.99|2015-02-26 10:47:00|80.737901233649083|4|73800400036|258|35.358252612079141|0|46|1699|-80.80146|387|35.17739|EVERYDAY (COOKIES)|0.0|14|BLACK & WHITE MINI COOKIE|506a6fdfb21d1e2beaeadfc6c26bf49646f91b72|4.2231534722856425|35.349871187060224|00738004000367|COOKIES|BAKERY|-80.737839|80.737953973863668|208|1
35.297134|64dcb1a597305e9eebc1769e00cb346f6cb36634|6.19|2014-09-11 12:45:00|80.737901233649083|4|8010000365|258|35.35825257386837|0|46|3045|-80.825175|1000|35.152722|BRAND-REVLON|1.0|17|REV XTRA LFE TOP COAT 216500|506a6fdfb21d1e2beaeadfc6c26bf49646f91b72|4.2231534722856425|35.349871187060224|00080100003651|COSMETICS|HBC|-80.737839|80.737981253740671|160|1
35.297134|43a7f08121fc6dd8429e6b6887c112209a8b3985|9.99|2014-11-11 07:44:00|80.737901233649083|4|3774114020|258|35.358252644719229|0|46|6965|-80.810056|1586|35.219587|GM READING GLASSES|0.0|18|JUST READERS DESIGNER|506a6fdfb21d1e2beaeadfc6c26bf49646f91b72|4.2231534722856425|35.349871187060224|00037741140245|READING GLASSES|GM|-80.737839|80.73792399921274|401|1
35.037115|65695b8c99ddbb936fa3abb61c0963c27c66d4e7|4.0|2014-09-18 09:51:00|80.805842308733688|4|84115200734|27|35.054353186293675|0|49|1165|-80.848528|87|35.053394|NFS-FRESH CONSUMER BUNCH|0.0|9|BUNCH- 3/$12 NOVELTY POMS|5231d2da48d0ffcf21e80fb567791b3612086f90|1.1911170444411914|35.053350220983141|00841152007345|FLORAL|FLORAL|-80.8062|80.80620045475446|11|1
35.037115|55659ab2ecc9f914c456e8ca24753e54f0b2ddad|3.29|2014-10-08 18:57:00|80.805842308733688|4|3000005040|27|35.054353185384002|0|49|12|-80.770346|2|35.052812|PANCAKE MIXES|0.0|1|AJEMIMA COMPLETE PANCAKE M|5231d2da48d0ffcf21e80fb567791b3612086f90|1.1911170444411914|35.053350220983141|00030000050705|BAKING MIXES|G1 GROCERY|-80.8062|80.806206855491965|40|1
35.037115|013334c8cec0ce85cdf363ed292830052eec6230|1.24|2014-09-30 18:19:00|80.805842308733688|4||27|35.054353185384002|0|49|502|-80.770346|64|35.052812|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5231d2da48d0ffcf21e80fb567791b3612086f90|1.1911170444411914|35.053350220983141|00204011000008|FRESH PRODUCE|PRODUCE|-80.8062|80.806206855491965|40|1
35.037115|891af6b98665bb9873efa3862a1d505b5ac858df|2.49|2014-11-11 10:40:00|80.805842308733688|4||27|35.054353185427679|0|49|512|-80.847383|64|35.024464|FRSH PROD FRSH FRUIT REM|0.0|4|COCONUTS|5231d2da48d0ffcf21e80fb567791b3612086f90|1.1911170444411914|35.053350220983141|00204262000000|FRESH PRODUCE|PRODUCE|-80.8062|80.806206689619628|317|1
35.037115|3bd8af6c0570bf37e2947075ee9200f95838d3e5|11.99|2015-03-01 16:06:00|80.805842308733688|4|8678511073|27|35.054353185384002|0|49|9969|-80.770346|887|35.052812|NFS-S/PREM-OTHER RED|0.0|13|ROSCATO ROSSO DOLCE|5231d2da48d0ffcf21e80fb567791b3612086f90|1.1911170444411914|35.053350220983141|00086785110738|SUPER PREMIUM ($11-$14.99)|WINE|-80.8062|80.806206855491965|40|1
35.037115|86c189133dd48555cc2828849f7fc637991f644f|1.29|2014-09-22 19:38:00|80.805842308733688|4|980000761|27|35.054353185384002|0|49|48|-80.770346|7|35.052812|REGISTER GUM|0.0|1|TIC TAC ORANGE BIG PACK|5231d2da48d0ffcf21e80fb567791b3612086f90|1.1911170444411914|35.053350220983141|00009800007639|CANDY|G1 GROCERY|-80.8062|80.806206855491965|40|1
35.037115|bbd1701e1a7e9c96ab0ece8b3dbe9e04e8e23df0|3.49|2014-10-27 19:14:00|80.805842308733688|4|2840024018|27|35.054353185384002|0|49|205|-80.770346|31|35.052812|REMAINING SNACKS|0.0|1|FUNYUNS|5231d2da48d0ffcf21e80fb567791b3612086f90|1.1911170444411914|35.053350220983141|00028400240185|SNACKS|G1 GROCERY|-80.8062|80.806206855491965|40|1
35.037115|0e530b9b5290016b6dec06b17345a63b18ffb499|3.19|2014-11-12 18:53:00|80.805842308733688|4|2100000028|27|35.054353185384002|0|49|316|-80.770346|52|35.052812|CREAM CHEESE|0.69|3|PHILLY FREE SOFT CREAM CHEESE|5231d2da48d0ffcf21e80fb567791b3612086f90|1.1911170444411914|35.053350220983141|00021000001545|CHEESE|DAIRY|-80.8062|80.806206855491965|40|1
35.037115|4f28b9dc01106b0f39c924b516bd9542976c99ea|1.23|2014-10-13 18:54:00|80.805842308733688|4||27|35.054353185384002|0|49|505|-80.770346|64|35.052812|FRESH SOFT FRUIT|0.13|4|BLACK PLUMS|5231d2da48d0ffcf21e80fb567791b3612086f90|1.1911170444411914|35.053350220983141|00204040000000|FRESH PRODUCE|PRODUCE|-80.8062|80.806206855491965|40|1
35.037115|f55a842218afc45c805ffb7f366438dde07a7607|4.0|2015-01-05 09:50:00|80.805842308733688|4|84115200700|27|35.054353185384002|0|49|1165|-80.770346|87|35.052812|NFS-FRESH CONSUMER BUNCH|0.0|9|BUNCH- MIXED DYED DAISIES|5231d2da48d0ffcf21e80fb567791b3612086f90|1.1911170444411914|35.053350220983141|00841152007000|FLORAL|FLORAL|-80.8062|80.806206855491965|40|1
35.037115|56164e6ff99df1fc3b4d2710eac784c251b47ebe|3.59|2014-10-15 19:11:00|80.805842308733688|4|7433610102|27|35.054353185384002|0|49|342|-80.770346|57|35.052812|FRESH MILK|0.0|3|HIGHLAND CREST WHOLE MILK|5231d2da48d0ffcf21e80fb567791b3612086f90|1.1911170444411914|35.053350220983141|00074336879203|MILK|DAIRY|-80.8062|80.806206855491965|40|1
35.037115|8143148e060891c8e0bd54a8a9d54289f066415c|1.29|2015-03-02 19:21:00|80.805842308733688|4|1254661959|27|35.054353185384002|0|49|48|-80.770346|7|35.052812|REGISTER GUM|0.0|1|TRIDENT SPEARMINT|5231d2da48d0ffcf21e80fb567791b3612086f90|1.1911170444411914|35.053350220983141|00012546615310|CANDY|G1 GROCERY|-80.8062|80.806206855491965|40|1
35.037115|32ad4f1cb834e4a2076a3d607e6e5e3d786681ac|2.99|2015-01-27 18:54:00|80.805842308733688|4|2100000028|27|35.054353185384002|0|49|316|-80.770346|52|35.052812|CREAM CHEESE|0.99|3|PHILLY LIGHT SOFT CRM CHEESE|5231d2da48d0ffcf21e80fb567791b3612086f90|1.1911170444411914|35.053350220983141|00021000000289|CHEESE|DAIRY|-80.8062|80.806206855491965|40|1
35.037115|3ae68150327989fad98f6ef411298453da968c42|2.99|2014-12-21 13:26:00|80.805842308733688|4|7027223202|27|35.054353185384002|0|49|323|-80.770346|57|35.052812|TOPPINGS-REFRIGERATED|0.0|3|REDDI WIP EXTRA CREAMY|5231d2da48d0ffcf21e80fb567791b3612086f90|1.1911170444411914|35.053350220983141|00070272232034|MILK|DAIRY|-80.8062|80.806206855491965|40|1
35.037115|ac427d0499697c0af8eff446b95861d1dd5c7dae|15.98|2015-01-19 19:20:00|80.805842308733688|4|3338314604|27|35.054353185384002|0|49|509|-80.770346|64|35.052812|FRESH CITRUS-REMAINING|6.0|4|CLEMENTINES 5LB BOX|5231d2da48d0ffcf21e80fb567791b3612086f90|1.1911170444411914|35.053350220983141|00033383146041|FRESH PRODUCE|PRODUCE|-80.8062|80.806206855491965|40|2
35.037115|40bccc44a747c6726e424a836cb3089c234c97d8|7.99|2015-01-14 18:45:00|80.805842308733688|4|3338314604|27|35.054353185384002|0|49|509|-80.770346|64|35.052812|FRESH CITRUS-REMAINING|3.0|4|CLEMENTINES 5LB BOX|5231d2da48d0ffcf21e80fb567791b3612086f90|1.1911170444411914|35.053350220983141|00033383146041|FRESH PRODUCE|PRODUCE|-80.8062|80.806206855491965|40|1
35.037115|b352e6cf0432296b7206d68b6cbd21dc5d628659|2.29|2015-01-09 18:14:00|80.805842308733688|4||27|35.054353185384002|0|49|561|-80.770346|64|35.052812|FR PROD ORGANIC PRODUCE|0.0|4|ORG BANANAS|5231d2da48d0ffcf21e80fb567791b3612086f90|1.1911170444411914|35.053350220983141|00294011000009|FRESH PRODUCE|PRODUCE|-80.8062|80.806206855491965|40|1
35.037115|756f912323ad9bf171d617e29f269dca05fb81b6|7.99|2014-10-05 17:51:00|80.805842308733688|4|7527890970|27|35.054353186253742|0|49|291|-80.760919|48|35.024332|FROZEN POUTLRY|0.0|5|FOSTER FARMS HOT N SPICY WINGS|5231d2da48d0ffcf21e80fb567791b3612086f90|1.1911170444411914|35.053350220983141|00075278909706|FROZEN MEALS|FROZEN|-80.8062|80.806201503526196|343|1
35.037115|aa89b61ea4c07eac6248f50aace5d7ec7ef84229|1.99|2014-12-24 09:21:00|1.4091206135396188|4||27|0.611513017149893|0|47|274|-80.8062|44|35.037115|ICE|0.0|5|HT BAGGED ICE|5231d2da48d0ffcf21e80fb567791b3612086f90|1.1911170444411914|0.61242566243833529|00072036480118|ICE|FROZEN|-80.8062|1.4103342460250419|27|1
35.037115|83272d5a2870ec51f2e9412ece961a4c5568a4ba|5.99|2014-09-18 09:57:00|80.805842308733688|4|902135050|27|35.054353186293675|0|49|480|-80.848528|87|35.053394|NFS-FLORAL,GARDENING-MIS|0.0|9|"10"" HARDY MUM"|5231d2da48d0ffcf21e80fb567791b3612086f90|1.1911170444411914|35.053350220983141|00009021350507|FLORAL|FLORAL|-80.8062|80.80620045475446|11|1
35.037115|de10964ae7ed27f7873b999e8f7125d63449df17|5.99|2014-09-18 10:07:00|80.805842308733688|4|902135050|27|35.054353186293675|0|49|480|-80.848528|87|35.053394|NFS-FLORAL,GARDENING-MIS|0.0|9|"10"" HARDY MUM"|5231d2da48d0ffcf21e80fb567791b3612086f90|1.1911170444411914|35.053350220983141|00009021350507|FLORAL|FLORAL|-80.8062|80.80620045475446|11|1
35.037115|9d4d237b88b6fa23dc1258a0c407e5ea403ef47a|4.29|2015-02-11 18:44:00|80.805842308733688|4|2840016014|27|35.054353185384002|0|49|201|-80.770346|31|35.052812|POTATO CHIPS|0.29|1|LAYS CLASSIC|5231d2da48d0ffcf21e80fb567791b3612086f90|1.1911170444411914|35.053350220983141|00028400160148|SNACKS|G1 GROCERY|-80.8062|80.806206855491965|40|1
35.037115|b21a7d4ca2c7181ae302fee65fcb32a34cc5a495|9.99|2015-01-17 19:09:00|1.4091206135396188|4|2370001118|27|0.611513017149893|0|47|291|-80.8062|48|35.037115|FROZEN POUTLRY|2.0|5|TYSON ANYTZR BUFFALO HOT WINGS|5231d2da48d0ffcf21e80fb567791b3612086f90|1.1911170444411914|0.61242566243833529|00023700011183|FROZEN MEALS|FROZEN|-80.8062|1.4103342460250419|27|1
35.444615|0d4fda5b5db2047331b08b09ee4c46003433a011|7.96|2015-01-25 13:51:00|1.4102725052409182|2|8660040320|340|0.6186252338517699|0|1|173|-80.861571|27|35.444615|CANNED POULTRY|2.96|1|B BEE PREM CHICKEN BRST|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00086600403205|PREPARED FOODS-RTS|G1 GROCERY|-80.861571|1.4113006522851637|340|4
35.444615|290f6b85c80471afdf69c6bff16e75c7af519980|2.0|2014-12-26 18:52:00|1.4102725052409182|2|7203605067|340|0.6186252338517699|0|1|60|-80.861571|9|35.444615|HOT CEREAL|0.33|1|HT OATS 18 QUCIK|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00072036050649|CEREAL|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.444615|5dbb01f08ec33b187a27c5449c7b79295ffe56e9|1.36|2014-10-23 13:58:00|1.4102725052409182|2||340|0.6186252338517699|0|1|502|-80.861571|64|35.444615|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|5731e0e3664e9f1e13c14a7534f3050f9c60a454|1.27|2015-02-21 20:25:00|1.4102725052409182|2||340|0.6186252338517699|0|1|502|-80.861571|64|35.444615|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|9b934bb09a984e7658b7e5db2dc0c89a51fc9d04|0.94|2015-01-24 16:28:00|80.86161257435397|2||340|35.477261455978947|0|36|502|-80.762919|64|35.442529|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|35.472272108304431|00204011000008|FRESH PRODUCE|PRODUCE|-80.861571|80.861588133595376|471|1
35.444615|fd57cf85c72ae3e0b1b4ce56e03f8a86f8c55545|1.47|2015-01-31 09:39:00|1.4102725052409182|2||340|0.6186252338517699|0|1|502|-80.861571|64|35.444615|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|97a2f3b4fdaf2d09625198c86ba0a3a575a9a507|1.48|2014-10-11 21:13:00|1.4102725052409182|2||340|0.6186252338517699|0|1|502|-80.861571|64|35.444615|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|f79f9bc17a17157f3459558d60ed4de4bad0efca|1.76|2014-10-16 15:20:00|1.4102725052409182|2||340|0.6186252338517699|0|1|502|-80.861571|64|35.444615|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|8c8e71a03d134aca4823a17d172caf9fd45bf161|0.83|2014-11-16 14:20:00|1.4102725052409182|2||340|0.6186252338517699|0|1|502|-80.861571|64|35.444615|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|659ea013111603297ab1c62e1f7827b662ad9a52|9.99|2014-12-29 16:08:00|1.4102725052409182|2|7203661016|340|0.6186252338517699|0|1|297|-80.861571|49|35.444615|GROUND BEEF|1.52|2|GROUND CHUCK 80% LEAN 2 LB|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00072036610164|BEEF|MEAT|-80.861571|1.4113006522851637|340|1
35.444615|223daa7ddb168de58d10b41fa4e48a96dacf00a4|2.59|2014-10-04 14:36:00|1.4102725052409182|2|7203655029|340|0.6186252338517699|0|1|331|-80.861571|52|35.444615|NATURAL SLICED|0.0|3|HT PROVOLONE SLICES|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00072036550170|CHEESE|DAIRY|-80.861571|1.4113006522851637|340|1
35.444615|ade5aa1bcad1dc2aca5d9099cc6170c76fb04802|2.89|2015-03-07 14:23:00|1.4102725052409182|2|7203655029|340|0.6186252338517699|0|1|331|-80.861571|52|35.444615|NATURAL SLICED|0.92|3|HT PROVOLONE SLICES|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00072036550170|CHEESE|DAIRY|-80.861571|1.4113006522851637|340|1
35.444615|f7c16bd3e7258adeacd4214061692f3ebb09fcc6|7.88|2014-12-13 21:20:00|1.4102725052409182|2|7203656065|340|0.6186252338517699|0|1|315|-80.861571|52|35.444615|CHEESE-PROCESSED-SLICED|0.0|3|HT 2% SINGLE WRAP CHEESE|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00072036600844|CHEESE|DAIRY|-80.861571|1.4113006522851637|340|4
35.444615|89ae0bd0036b6bbe590ba8842ce9b53ba7f62152|2.27|2015-01-11 13:51:00|1.4102725052409182|2|7203656065|340|0.6186252338517699|0|1|315|-80.861571|52|35.444615|CHEESE-PROCESSED-SLICED|0.0|3|HT 2% SINGLE WRAP CHEESE|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00072036600844|CHEESE|DAIRY|-80.861571|1.4113006522851637|340|1
35.444615|6d329f2f535025ed1293a85e4ea6f0f480737dcc|4.54|2015-01-27 20:13:00|80.86161257435397|2|7203656065|340|35.477261456422909|0|36|315|-80.782849|52|35.372142|CHEESE-PROCESSED-SLICED|0.0|3|HT 2% SINGLE WRAP CHEESE|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|35.472272108304431|00072036600844|CHEESE|DAIRY|-80.861571|80.861586807149422|122|2
35.444615|94f10d831c895a37239f31d57e1efb33fcde51be|5.9|2015-02-26 13:03:00|80.86161257435397|2|7203663125|340|35.477261444606086|0|36|1262|-80.780702|57|35.318911|HALF N HALF WHIPPING CREAM|0.0|3|HT LIGHT WHIPPING CREAM|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|35.472272108304431|00072036630995|MILK|DAIRY|-80.861571|80.861608587849247|167|2
35.444615|7863f0a4e7d90390fbaf5645d87a0f4da839b5df|0.5|2014-11-14 18:13:00|1.4102725052409182|2||340|0.6186252338517699|0|1|543|-80.861571|64|35.444615|FRESH GARLIC|0.0|4|COO GARLIC, WHITE, BULK|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00204608000008|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|d190c970a1088156542459d8b7f5a612cf3d074d|2.49|2014-12-23 14:09:00|1.4102725052409182|2|4369505631|340|0.6186252338517699|0|1|1276|-80.861571|279|35.444615|FROZEN SANDWICHES|0.49|5|HOT PKT CHEESEBURGER SANDWICH|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00043695071238|FROZEN SANDWICH AND SNACKS|FROZEN|-80.861571|1.4113006522851637|340|1
35.444615|cadcc3095c6aa1e8db4090c9d0131e37353bcf26|9.38|2014-12-16 21:43:00|1.4102725052409182|2|4900002468|340|0.6186252338517699|0|1|54|-80.861571|8|35.444615|DIET|4.69|23|DIET COKE .5 LITER/6 PK.|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.861571|1.4113006522851637|340|2
35.444615|1344d9862c66c78e2003a642aec0b182fbeaf368|4.99|2015-02-11 20:44:00|80.86161257435397|2|4900002468|340|35.477261455978947|0|36|54|-80.762919|8|35.442529|DIET|0.65|23|DIET COKE .5 LITER/6 PK.|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|35.472272108304431|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.861571|80.861588133595376|471|1
35.444615|69857af73752972a0780f8bf213425146578869c|1.99|2014-11-09 16:40:00|1.4102725052409182|2|5100017520|340|0.6186252338517699|0|1|1201|-80.861571|33|35.444615|RTS CANNED|0.49|1|CAM HOMESTYLE CREOLE CHICKEN|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00051000195647|SOUP|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.444615|7afcd4784b3ecb4c2702199fec5e03bc7479be17|1.72|2014-09-21 18:13:00|1.4102725052409182|2||340|0.6186252338517699|0|1|502|-80.861571|64|35.444615|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|5f83e44e0e0389ff2bc68a7925cdfe1da06bfe32|1.32|2015-02-06 19:29:00|80.86161257435397|2||340|35.477261455978947|0|36|502|-80.762919|64|35.442529|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|35.472272108304431|00204011000008|FRESH PRODUCE|PRODUCE|-80.861571|80.861588133595376|471|1
35.444615|7225d541c51c0c002ec99f54f78f3ff4ee9a5f10|1.58|2014-09-15 22:53:00|80.86161257435397|2||340|35.477261456788234|0|36|502|-80.86175|64|35.40953|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|35.472272108304431|00204011000008|FRESH PRODUCE|PRODUCE|-80.861571|80.861585625746713|209|1
35.444615|e2b22b6eb7b40474c553005cd21493a98c34735d|2.07|2014-09-27 14:08:00|1.4102725052409182|2||340|0.6186252338517699|0|1|502|-80.861571|64|35.444615|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|92ccbdf71e92021ecf9edd3ba82c4985ace39bf0|11.38|2014-09-13 15:00:00|1.4102725052409182|2|1450000711|340|0.6186252338517699|0|1|1274|-80.861571|50|35.444615|BAG VEG PROTEIN|2.84|5|BE VOILA TERIYAKI CHICKEN|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00014500007148|VEGETABLES-FROZEN|FROZEN|-80.861571|1.4113006522851637|340|2
35.444615|6faf0cb5d9b8935355834def3fe36bfca2993613|3.79|2014-12-27 08:50:00|1.4102725052409182|2|7203603030|340|0.6186252338517699|0|1|4296|-80.861571|1205|35.444615|ACETAMINOPHEN|0.0|17|HT ACETAMINOPHEN CAPS 24CT|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00072036030306|PAIN RELIEF|HBC|-80.861571|1.4113006522851637|340|1
35.444615|e447a28fd0e5387168f1176e40d3d228fa499fbd|2.69|2015-01-03 11:41:00|1.4102725052409182|2|7203608053|340|0.6186252338517699|0|1|78|-80.861571|11|35.444615|MUSTARD|0.8|1|HT MUSTARD DIJON CLASSIC|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00072036080554|CONDIMENTS|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.444615|0553baf8b0732b93b551a7f74b68ac8258813041|20.950000000000003|2014-10-20 20:14:00|80.86161257435397|2|2000012636|340|35.477261455978947|0|36|1275|-80.762919|50|35.442529|BOX VEG|12.0|5|GG ASPARAGUS CUTS NO SAUCE|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|35.472272108304431|00020000126364|VEGETABLES-FROZEN|FROZEN|-80.861571|80.861588133595376|471|5
35.444615|0ab90784cd78c76668e88d44f77db3e5759c9943|5.49|2015-02-28 17:12:00|1.4102725052409182|2|7597116682|340|0.6186252338517699|0|1|1837|-80.861571|420|35.444615|FFM PRESLICED MEATS|5.49|6|FRESH FOOD ROASTED TURKEY BRST|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00072036959867|PRESLICED MEAT|DELI|-80.861571|1.4113006522851637|340|1
35.444615|768d1d48539307d84f501de111bc9c6fd8d6a063|1.0|2015-01-27 14:41:00|1.4102725052409182|2|4000000435|340|0.6186252338517699|0|1|47|-80.861571|7|35.444615|REGISTER BARS|0.5|1|(FE)TWIX CARAMEL COOKIE BAR|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00040000004356|CANDY|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.444615|f1c9fef2db4d8c5a4e6689f80211a7b7f656cd63|3.19|2014-10-24 20:23:00|80.86161257435397|2|20139200000|340|35.477261455978947|0|36|296|-80.762919|49|35.442529|RANCHER BEEF|0.0|2|BEEF TENDERLOIN TIPS|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|35.472272108304431|00201392000009|BEEF|MEAT|-80.861571|80.861588133595376|471|1
35.444615|3cb63285e546b0e4d48da4243699d1e43a298baa|3.99|2015-02-06 19:25:00|80.86161257435397|2|7073405372|340|35.477261455978947|0|36|232|-80.762919|37|35.442529|WELLNESS TEA|0.0|1|CELESTIAL WELL SLPY THROAT TMR|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|35.472272108304431|00070734513701|TEA|G1 GROCERY|-80.861571|80.861588133595376|471|1
35.444615|e2090efec3a5eedd329ad42e82e517f9aa3f7c88|3.99|2015-02-25 19:50:00|80.86161257435397|2|4610000094|340|35.477261455978947|0|36|318|-80.762919|52|35.442529|SHREDDED/GRATED CHEESE|2.0|3|SARGENTO CB 6 CHEESE ITALIAN|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|35.472272108304431|00046100000915|CHEESE|DAIRY|-80.861571|80.861588133595376|471|1
35.444615|375299ab71dd53744843c82e63906e5b8f887322|3.25|2014-11-14 16:35:00|1.4102725052409182|2|7203656080|340|0.6186252338517699|0|1|318|-80.861571|52|35.444615|SHREDDED/GRATED CHEESE|0.0|3|HT SHRED SHARP CHED CHEESE 2%|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00072036590466|CHEESE|DAIRY|-80.861571|1.4113006522851637|340|1
35.444615|788917f07e5c37d4f397e8a6e200463ae9011daf|6.5|2015-02-10 14:29:00|80.86161257435397|2|7203656080|340|35.477261455978947|0|36|318|-80.762919|52|35.442529|SHREDDED/GRATED CHEESE|0.0|3|HT SHRED SHARP CHED CHEESE 2%|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|35.472272108304431|00072036590466|CHEESE|DAIRY|-80.861571|80.861588133595376|471|2
35.444615|2aa0aaee4552b407be1a2c5b31c319cc2b0c79cb|4.99|2014-12-17 17:43:00|1.4102725052409182|2|3338307764|340|0.6186252338517699|0|1|500|-80.861571|64|35.444615|FRESH APPLES|0.0|4|GALA APPLES 3LB BAG|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00072036880314|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|f0945f61c90b0ad302253c607ef6064d3451ad2e|3.99|2015-01-20 15:19:00|1.4102725052409182|2|7203659054|340|0.6186252338517699|0|1|499|-80.861571|110|35.444615|MEATBALLS|1.32|19|HT HOMESTYLE MEATBALLS|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00072036590541|FROZEN CASE MEAT|CASE READY MEATS|-80.861571|1.4113006522851637|340|1
35.444615|4e378a720b405d66002113f293a61dc43711f504|3.29|2014-12-01 20:32:00|80.86161257435397|2|85591900302|340|35.477261455978947|0|36|41|-80.762919|6|35.442529|BREAKFAST BARS|1.65|1|S BCH CEREAL BAR PROT FIT PB|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|35.472272108304431|00855919003013|BREAKFAST FOODS|G1 GROCERY|-80.861571|80.861588133595376|471|1
35.444615|55d6ee8f113fec976d712ebeec3dbb9ed7428c13|3.99|2015-02-09 20:27:00|80.86161257435397|2|7203670859|340|35.477261455978947|0|36|1280|-80.762919|48|35.442529|MULTI SERVE MEALS|0.99|5|HTT CHICKEN STIR FRY|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|35.472272108304431|00072036708595|FROZEN MEALS|FROZEN|-80.861571|80.861588133595376|471|1
35.444615|89839c1f371a843159a0f0dc656b54a7cc6bfe32|3.25|2015-03-02 13:22:00|1.4102725052409182|2|7203656080|340|0.6186252338517699|0|1|318|-80.861571|52|35.444615|SHREDDED/GRATED CHEESE|0.0|3|HT SHREDDED MOZZ/PROVLONE|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00072036705174|CHEESE|DAIRY|-80.861571|1.4113006522851637|340|1
35.444615|29a83555d323a12fbf1d89c62376bf40f3d427ef|3.79|2014-11-18 21:35:00|1.4102725052409182|2|5565364600|340|0.6186252338517699|0|1|92|-80.861571|13|35.444615|REMAINING CRACKERS|0.79|1|BRETON MINI ORIG CRACKERS|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00055653646006|CRACKERS|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.444615|8751dcd3582c070fc6518df91ccd020d34597ae3|5.39|2014-10-02 15:31:00|1.4102725052409182|2|7192167217|340|0.6186252338517699|0|1|254|-80.861571|892|35.444615|PREMIUM PIZZA|2.7|5|TOMBSTONE 12IN ORG SAUS&PEPP|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00071921561970|FROZEN PIZZA|FROZEN|-80.861571|1.4113006522851637|340|1
35.444615|440721dfffd70377be95827bf96d659e838fe781|9.99|2015-02-15 16:47:00|80.86161257435397|2|84560401578|340|35.477261444606086|0|36|6984|-80.780702|1600|35.318911|VALENTINE NOVELTY-IMPORT|7.49|18|I/O VAL RAZOR CHILLER 18OZ|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|35.472272108304431|00845604015780|SEASONAL MERCHANDISE|GM|-80.861571|80.861608587849247|167|1
35.444615|d278377b1838d2cabfedcc2be56ef1b9babf86da|5.69|2014-12-03 19:33:00|80.86161257435397|2|5190001602|340|35.477261455978947|0|36|839|-80.762919|102|35.442529|STACK PACKS|0.0|19|LOF PREMIUM SMOKED HAM|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|35.472272108304431|00051900016011|LUNCHMEATS|CASE READY MEATS|-80.861571|80.861588133595376|471|1
35.444615|1901a335f11b1aafb31a7a85df0e70945ce59ac3|3.94|2014-09-12 19:46:00|80.86161257435397|2|7203629075|340|35.477261455978947|0|36|1211|-80.762919|272|35.442529|HISP SALSA/DIPS|0.0|1|HT SALSA MEDIUM|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|35.472272108304431|00072036290755|HISPANIC PREP. FOODS|G1 GROCERY|-80.861571|80.861588133595376|471|2
35.444615|6784492583741e41c95d3a9f4cd64c019547f119|4.29|2014-10-12 21:41:00|1.4102725052409182|2|70897141855|340|0.6186252338517699|0|1|1703|-80.861571|387|35.444615|SEASONAL COOKIES|0.8|14|BOO PURPLE FRSTD SUGAR COOKIES|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00708971418557|COOKIES|BAKERY|-80.861571|1.4113006522851637|340|1
35.444615|e60dd60b312fbdf83d5a61513dad3cc67d011523|2.85|2014-11-03 11:05:00|1.4102725052409182|2|4133500053|340|0.6186252338517699|0|1|184|-80.861571|28|35.444615|SALAD DRESSINGS-LIQUID|0.0|1|KENS DRS LT HONEY MUSTARD|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|0.61833652052202714|00041335335177|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.444615|1729c9c94a84bbd2d84df55dffe95dda58f46fd7|2.19|2014-09-16 22:10:00|80.86161257435397|2|4900005010|340|35.477261444674177|0|36|55|-80.814133|8|35.333742|REGULAR|0.2|23|CLASSIC COKE 2 LT CONTOUR|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|35.472272108304431|00049000050103|CARBONATED BEVERAGES|BEVERAGE|-80.861571|80.861608498598827|472|1
35.444615|76402da88712dd8d4313bfa0d746a49f1bffeab5|2.19|2014-11-07 20:15:00|80.86161257435397|2|4900005010|340|35.477261455978947|0|36|55|-80.762919|8|35.442529|REGULAR|0.2|23|SPRITE  2 LITER|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|35.472272108304431|00049000050158|CARBONATED BEVERAGES|BEVERAGE|-80.861571|80.861588133595376|471|1
35.444615|b1791c10b3b3b7ab873d11261c1b69e0c4ebf0ef|10.3|2014-10-08 20:06:00|80.86161257435397|2|7218063473|340|35.477261455978947|0|36|284|-80.762919|892|35.442529|SUPER PREMIUM PIZZA|4.3|5|RED BARON RISING SAU&PEPP PZZA|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|35.472272108304431|00072180567345|FROZEN PIZZA|FROZEN|-80.861571|80.861588133595376|471|2
35.444615|2e1a5b7e06569606a797eac7fccc42983c4c352b|7.98|2015-03-02 21:54:00|80.86161257435397|2|4610000012|340|35.477261455978947|0|36|318|-80.762919|52|35.442529|SHREDDED/GRATED CHEESE|1.99|3|SARGENTO OTB MOZZA FINE CUT|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|35.472272108304431|00046100000557|CHEESE|DAIRY|-80.861571|80.861588133595376|471|2
35.444615|019872ac0df2c6585e6af0dcfeca9ddf7159ffc1|5.78|2014-11-05 20:22:00|80.86161257435397|2|7203655029|340|35.477261455978947|0|36|331|-80.762919|52|35.442529|NATURAL SLICED|1.45|3|HT PROVOLONE 2% SLICES|5333d453cd602e6a66918ffa21dc58cded5d618b|2.255791475881002|35.472272108304431|00072036983978|CHEESE|DAIRY|-80.861571|80.861588133595376|471|2
35.219587|1e82915e97d149a9e9235cdec874e0d563b919bd|3.49|2014-10-01 20:09:00|80.810069425230125|3|4000024947|401|35.24504930456466|0|23|52|-80.85013|7|35.175855|PKG NON CHOC|0.0|1|STARBURST FAVEREDS LAYDWN BAG|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00040000329688|CANDY|G1 GROCERY|-80.810056|80.810075837400746|218|1
35.219587|9040c5ae6b394a0b994b6a62845683c6d4fd4e9a|4.49|2014-12-02 20:44:00|80.810069425230125|3|4000031532|401|35.24504930456466|0|23|727|-80.85013|7|35.175855|SEASONAL CANDY-SINGLE FAC|0.8|1|I/O(C14)M&M PLAIN CHRISTMAS|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00040000315322|CANDY|G1 GROCERY|-80.810056|80.810075837400746|218|1
35.219587|b12dffd0e76677b7a3535ba118ccfc46d87b8e05|0.79|2014-10-30 16:29:00|80.810069425230125|3||401|35.24504930456466|0|23|532|-80.85013|64|35.175855|FRESH CUCUMBERS|0.0|4|COO CUCUMBERS S/S|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00204062000002|FRESH PRODUCE|PRODUCE|-80.810056|80.810075837400746|218|1
35.219587|212901f4f7eac07eff39e938cbd7df7e526d2dad|4.0|2014-11-22 13:48:00|80.810069425230125|3|66440100015|401|35.24504930456466|0|23|1165|-80.85013|87|35.175855|NFS-FRESH CONSUMER BUNCH|0.0|9|BUNCH- HYPERIUCM ASST.|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00664401000153|FLORAL|FLORAL|-80.810056|80.810075837400746|218|1
35.219587|e905f20f1756de32c93ce61ad13c5f343a648c0b|7.96|2015-01-11 18:33:00|80.810069425230125|3|78616233800|401|35.24504930456466|0|23|31|-80.85013|4|35.175855|NON CARBONATED WATER|2.96|1|CB SMARTWATER 1 LTR PET SINGLE|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00786162338006|BOTTLED WATER|G1 GROCERY|-80.810056|80.810075837400746|218|4
35.219587|6ee83d3858ebbca826e94be455c58e960ff7ef03|7.96|2015-01-30 16:58:00|80.810069425230125|3|78616233800|401|35.24504930456466|0|23|31|-80.85013|4|35.175855|NON CARBONATED WATER|2.96|1|CB SMARTWATER 1 LTR PET SINGLE|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00786162338006|BOTTLED WATER|G1 GROCERY|-80.810056|80.810075837400746|218|4
35.219587|842a9d07fb67d29e087724aa4bd517e97d647c6b|9.95|2015-02-21 15:47:00|80.810069425230125|3|78616233800|401|35.24504930456466|0|23|31|-80.85013|4|35.175855|NON CARBONATED WATER|4.95|1|CB SMARTWATER 1 LTR PET SINGLE|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00786162338006|BOTTLED WATER|G1 GROCERY|-80.810056|80.810075837400746|218|5
35.219587|231627504125a733db9006371063dfc073ebff7c|7.99|2015-01-15 21:28:00|80.810069425230125|3|78436948375|401|35.24504930456466|0|23|6911|-80.85013|1582|35.175855|DOG TOYS|0.0|18|LAMB CHOP DOG TOY|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00784369483758|PET NEEDS|GM|-80.810056|80.810075837400746|218|1
35.219587|03d7f786c9e60d6c371cdeded5b468c5c91ea998|3.25|2014-11-15 13:24:00|80.810069425230125|3|7203656080|401|35.24504930456466|0|23|318|-80.85013|52|35.175855|SHREDDED/GRATED CHEESE|0.0|3|HT FANCY SHRED MILD CHED CHES|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00072036560810|CHEESE|DAIRY|-80.810056|80.810075837400746|218|1
35.219587|561334d7594d8454f81841a1d605986c0923018c|6.59|2015-03-01 16:51:00|80.810069425230125|3|7940035291|401|35.245049308383152|0|23|3814|-80.826724|1070|35.195689|INVISIBLE-FEMALE|1.6|17|DOVE CLR TONE SOLID A/P PNK RS|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00079400362520|DEODORANT|HBC|-80.810056|80.810066102972343|412|1
35.219587|cf69f6852944c81cf893d9f3dd5180a028a033cf|2.49|2014-10-12 19:10:00|80.810069425230125|3|1380017219|401|35.24504930456466|0|23|1278|-80.85013|48|35.175855|SINGLE SERVE NUTRITIONAL|0.0|5|LC FETTUCINI ALFREDO|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00013800166517|FROZEN MEALS|FROZEN|-80.810056|80.810075837400746|218|1
35.219587|acd8d13a1d1191e6f6e9aa2e474a9bac6b9372bf|2.79|2014-09-14 18:06:00|80.810069425230125|3|1600042060|401|35.24504930456466|0|23|13|-80.85013|2|35.175855|ROLLS/BISCUIT MIXES|1.29|1|BC BISQUICK|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00016000420601|BAKING MIXES|G1 GROCERY|-80.810056|80.810075837400746|218|1
35.219587|9ee78cf4b32dbcdb52c74461d1fe243a1d3f5459|2.59|2014-12-11 19:13:00|80.810069425230125|3|1480000034|401|35.24504930456466|0|23|128|-80.85013|20|35.175855|APPLE JUICE-SHELF|0.0|1|MOTTS 100% PURE APPLE JUICE|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00014800000344|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.810056|80.810075837400746|218|1
35.219587|5019587febe0fa817c2047bdf8418a5baf826ddc|6.99|2014-11-06 18:52:00|80.810069425230125|3|81651201395|401|35.24504930456466|0|23|141|-80.85013|21|35.175855|TRAIL MIXES AND BLENDS|1.0|1|I/O CS MILK CHOC PEPP PRETZEL|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00816512013953|NUTS|G1 GROCERY|-80.810056|80.810075837400746|218|1
35.219587|d39fbda225a03fe0798382229ecbcd51501e65db|2.89|2015-02-16 19:05:00|80.810069425230125|3|7203655029|401|35.24504930456466|0|23|331|-80.85013|52|35.175855|NATURAL SLICED|1.22|3|HT PROVOLONE SLICES|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00072036550170|CHEESE|DAIRY|-80.810056|80.810075837400746|218|1
35.219587|e51cbc2d8dc9f48761faf4f49181809d7d93d515|2.99|2015-02-02 19:02:00|80.810069425230125|3|7172000611|401|35.24504930456466|0|23|52|-80.85013|7|35.175855|PKG NON CHOC|0.0|1|TOOTSIE ROLL MIDGEES|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00071720006115|CANDY|G1 GROCERY|-80.810056|80.810075837400746|218|1
35.219587|342ca37261116d71685a9353d7b710e298dd7d63|6.49|2014-12-01 19:51:00|80.810069425230125|3|1200080994|401|35.24504930456466|0|23|54|-80.85013|8|35.175855|DIET|1.5|23|DT MTN DEW FRIDGEMATE|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00012000809972|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.810075837400746|218|1
35.219587|687e92baaea096ad8c555d45a383db390ecc6d0d|13.58|2015-01-24 17:26:00|80.810069425230125|3|1200080994|401|35.24504930456466|0|23|54|-80.85013|8|35.175855|DIET|3.4|23|DT MTN DEW FRIDGEMATE|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00012000809972|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.810075837400746|218|2
35.219587|ee03301e868aebfecbbecb580192474a864eace7|6.79|2015-02-10 15:35:00|80.810069425230125|3|1200080994|401|35.24504930456466|0|23|54|-80.85013|8|35.175855|DIET|1.8|23|DT MTN DEW FRIDGEMATE|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00012000809972|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.810075837400746|218|1
35.219587|a95254ea83a94f634920533634e4058b32dc8283|6.99|2015-03-09 17:23:00|80.810069425230125|3|1200080994|401|35.24504930456466|0|23|54|-80.85013|8|35.175855|DIET|2.0|23|DT MTN DEW FRIDGEMATE|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00012000809972|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.810075837400746|218|1
35.219587|560eb8c7be425a2c5b8bde13145197b8bd3b3cf1|6.49|2014-09-10 20:40:00|80.810069425230125|3|1200080994|401|35.24504930456466|0|23|54|-80.85013|8|35.175855|DIET|3.74|23|DT MTN DEW FRIDGEMATE|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00012000809972|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.810075837400746|218|1
35.219587|75edb6db9e0380bb144a35932efe09159647488f|9.58|2014-12-14 18:40:00|80.810069425230125|3|1200010041|401|35.24504930456466|0|23|54|-80.85013|8|35.175855|DIET|2.4|23|DIET MTN DEW 16 OZ 6 PK|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00012000107061|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.810075837400746|218|2
35.219587|6419cc7e1f11782066ad319f8702a8e42e5d7abc|6.49|2014-09-20 21:51:00|80.810069425230125|3|1200080994|401|35.24504930456466|0|23|54|-80.85013|8|35.175855|DIET|1.5|23|DT MTN DEW FRIDGEMATE|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00012000809972|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.810075837400746|218|1
35.219587|818680fc25df2fb0b026555df8f42fb5d98adddd|6.49|2014-11-13 21:03:00|80.810069425230125|3|1200080994|401|35.24504930456466|0|23|54|-80.85013|8|35.175855|DIET|1.5|23|DT MTN DEW FRIDGEMATE|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00012000809972|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.810075837400746|218|1
35.219587|a2ffa84377caa37925acec566ddf4a3870025537|6.49|2014-11-01 20:34:00|80.810069425230125|3|1200080994|401|35.24504930456466|0|23|54|-80.85013|8|35.175855|DIET|1.5|23|DT MTN DEW FRIDGEMATE|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00012000809972|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.810075837400746|218|1
35.219587|0a0f9366b6741f8fc917de0a631144ca098e176b|9.58|2014-10-08 19:40:00|80.810069425230125|3|1200010041|401|35.24504930456466|0|23|54|-80.85013|8|35.175855|DIET|2.39|23|DIET MTN DEW 16 OZ 6 PK|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00012000107061|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.810075837400746|218|2
35.219587|085ad21df66a78c08bb4b387ac66675104cd49da|13.98|2015-02-26 19:19:00|80.810069425230125|3|1200080994|401|35.24504930456466|0|23|54|-80.85013|8|35.175855|DIET|3.5|23|DT MTN DEW FRIDGEMATE|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00012000809972|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.810075837400746|218|2
35.219587|e76419e356a0d4c5f07b0537563cb5a32850f173|6.49|2014-10-21 18:37:00|80.810069425230125|3|1200080994|401|35.24504930456466|0|23|54|-80.85013|8|35.175855|DIET|1.5|23|DT MTN DEW FRIDGEMATE|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00012000809972|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.810075837400746|218|1
35.219587|f4bec637af6cd62c1b3aa4bccba85d93b0a2f4a4|4.99|2015-02-08 12:56:00|80.810069425230125|3|4242101480|401|35.24504930456466|0|23|482|-80.85013|100|35.175855|PRECOOKED BACON|0.6|19|BOARS HEAD FULLY COOKED BACON|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00042421014808|BACON|CASE READY MEATS|-80.810056|80.810075837400746|218|1
35.219587|f5f6835078fa5ff5accb9c3a8374fe8aa0f3bc31|0.91|2014-11-18 16:16:00|80.810069425230125|3||401|35.24504930456466|0|23|502|-80.85013|64|35.175855|FRESH BANANAS|0.0|4|BANANAS, YELLOW|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00204011000008|FRESH PRODUCE|PRODUCE|-80.810056|80.810075837400746|218|1
35.219587|43fc0b9240e1d70822d2ebaf039b12467efc8dd5|0.27|2015-01-20 18:00:00|80.810069425230125|3||401|35.24504930456466|0|23|502|-80.85013|64|35.175855|FRESH BANANAS|0.0|4|BANANAS, YELLOW|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00204011000008|FRESH PRODUCE|PRODUCE|-80.810056|80.810075837400746|218|1
35.219587|a568977c786f7de7622c9b636eef6c45cf41b931|5.58|2014-12-17 19:40:00|80.810069425230125|3|5964200343|401|35.24504930456466|0|23|52|-80.85013|7|35.175855|PKG NON CHOC|0.0|1|DUBBLE BUBBLE ORIGINAL 1LB BAG|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00059642003436|CANDY|G1 GROCERY|-80.810056|80.810075837400746|218|2
35.219587|8b3cdd4e5211c71e771a6d74ba8a987747ab0e95|5.98|2014-12-06 18:49:00|80.810069425230125|3|1070010541|401|35.24504930456466|0|23|727|-80.85013|7|35.175855|SEASONAL CANDY-SINGLE FAC|0.98|1|I/O(C14)JOLLY RNCH CNDY CANE|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00010700105417|CANDY|G1 GROCERY|-80.810056|80.810075837400746|218|2
35.219587|595f103b39090b362307214421147e14961a005b|9.69|2015-01-09 19:58:00|80.810069425230125|3|1780057309|401|35.24504930456466|0|23|156|-80.85013|24|35.175855|NFS-DOG FOOD-DRY|0.0|1|PURINA ONE CHICKEN & RICE|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00017800475556|PET FOOD/SUPPLIES|G1 GROCERY|-80.810056|80.810075837400746|218|1
35.219587|08eee1b00167c3f48596b85f030eb6e55498e576|19.38|2014-12-13 19:55:00|80.810069425230125|3|1780057309|401|35.24504930456466|0|23|156|-80.85013|24|35.175855|NFS-DOG FOOD-DRY|0.0|1|PURINA ONE CHICKEN & RICE|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00017800475556|PET FOOD/SUPPLIES|G1 GROCERY|-80.810056|80.810075837400746|218|2
35.219587|7115c7dc2a22dbb0a53104c140ec785abec2db35|9.69|2014-11-11 22:14:00|80.810069425230125|3|1780057309|401|35.24504930456466|0|23|156|-80.85013|24|35.175855|NFS-DOG FOOD-DRY|0.0|1|PURINA ONE CHICKEN & RICE|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00017800475556|PET FOOD/SUPPLIES|G1 GROCERY|-80.810056|80.810075837400746|218|1
35.219587|09351c617eb91b046e7e6d1fd82b4b50e6cb6aea|9.99|2015-02-21 21:20:00|80.810069425230125|3|1820053047|401|35.245049308383152|0|23|455|-80.826724|82|35.195689|DOMESTIC PREMIUM 12PK&>|0.0|16|BUD LIGHT 12PK 12OZ CAN|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00018200530470|DOMESTIC BEER|BEER|-80.810056|80.810066102972343|412|1
35.219587|6f39cf2279be3dbc57aa46777c377f7508cfda73|9.69|2014-09-21 15:46:00|80.810069425230125|3|1780057309|401|35.24504930456466|0|23|156|-80.85013|24|35.175855|NFS-DOG FOOD-DRY|0.0|1|PURINA ONE CHICKEN & RICE|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00017800475556|PET FOOD/SUPPLIES|G1 GROCERY|-80.810056|80.810075837400746|218|1
35.219587|fc2d5bd08807fac541667c2d96564e9c8c9e233b|9.69|2015-02-25 15:13:00|80.810069425230125|3|1780057309|401|35.24504930456466|0|23|156|-80.85013|24|35.175855|NFS-DOG FOOD-DRY|0.0|1|PURINA ONE CHICKEN & RICE|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00017800475556|PET FOOD/SUPPLIES|G1 GROCERY|-80.810056|80.810075837400746|218|1
35.219587|033e5c3b61e98c4e2019f40ff8c731d5dff41d87|1.79|2014-10-10 23:19:00|80.810069425230125|3|2430004101|401|35.24504930456466|0|23|1044|-80.85013|173|35.175855|SW BAKD GOOD SNACK CAKES|0.0|7|LD HONEY BUNS|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00024300041020|SWEET BAKED GOODS|COMMERCIAL BAKERY|-80.810056|80.810075837400746|218|1
35.219587|4ddb7d95d32c6cff609c0af808dcdd0e3e5391dd|4.99|2014-09-20 21:50:00|80.810069425230125|3|72527434190|401|35.24504930456466|0|23|6785|-80.85013|1568|35.175855|MAGAZINES WEEKLY|0.0|18|US WEEKLY|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00725274341900|MAGAZINES|GM|-80.810056|80.810075837400746|218|1
35.219587|d700586a202de419506cc3afbdc19cab83c7f65e|4.99|2014-11-22 13:44:00|80.810069425230125|3|2840008313|401|35.24504930456466|0|23|204|-80.85013|31|35.175855|TORTILLA CHIPS|1.0|1|TOSTITOS RSTC FAMILY SIZE|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00028400083133|SNACKS|G1 GROCERY|-80.810056|80.810075837400746|218|1
35.219587|c095a81e23c623e6de909df3651be30916656df7|1.49|2014-12-17 12:20:00|80.810069425230125|3|2200001567|401|35.24504930456466|0|23|727|-80.85013|7|35.175855|SEASONAL CANDY-SINGLE FAC|0.0|1|I/O(C14)STRBURST FAVRED CNDYCN|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00022000015679|CANDY|G1 GROCERY|-80.810056|80.810075837400746|218|1
35.219587|5e6fa79946ce5af5f7d2cbc78e96f4e64e7e73fb|10.99|2014-11-12 19:10:00|80.810069425230125|3|3600038585|401|35.24504930456466|0|23|427|-80.85013|72|35.175855|NFS-TOILET TISSUE|0.0|1|COTTONELLE CLEAN CARE 9RL|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00036000385670|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.810056|80.810075837400746|218|1
35.219587|990e8228fdf36b91230ae5b39943c7de623cd30f|7.99|2015-01-05 18:22:00|80.810069425230125|3|5200020805|401|35.24504930456466|0|23|171|-80.85013|20|35.175855|ISOTONIC DRINKS|2.01|1|GATORADE G2 ORANGE 8PK|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00052000208726|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.810056|80.810075837400746|218|1
35.219587|aa5dc78c8d59cc2646f6d0cd575ce6b2802a1a39|15.98|2014-10-25 16:11:00|80.810069425230125|3|5200020805|401|35.24504930456466|0|23|171|-80.85013|20|35.175855|ISOTONIC DRINKS|4.02|1|GATORADE GLACIER FREEZ 8PK|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00052000200218|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.810056|80.810075837400746|218|2
35.219587|7d3202aba92f353c3cdeb26cc8c45274ab43372f|7.99|2015-02-20 18:28:00|80.810069425230125|3|5200020805|401|35.24504930456466|0|23|171|-80.85013|20|35.175855|ISOTONIC DRINKS|2.99|1|GATORADE GLACIER FREEZ 8PK|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00052000200218|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.810056|80.810075837400746|218|1
35.219587|5b920e125caf7face99e42df2c3b18d170e13f37|7.99|2015-02-18 14:48:00|80.810069425230125|3|5200020805|401|35.24504930456466|0|23|171|-80.85013|20|35.175855|ISOTONIC DRINKS|2.99|1|GATORADE GLACIER FREEZ 8PK|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00052000200218|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.810056|80.810075837400746|218|1
35.219587|a06c98ee4feacab5be68fca9f0bc7be410837b1d|7.99|2015-02-06 19:29:00|80.810069425230125|3|5200020805|401|35.24504930456466|0|23|171|-80.85013|20|35.175855|ISOTONIC DRINKS|2.01|1|GATORADE GLACIER FREEZ 8PK|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00052000200218|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.810056|80.810075837400746|218|1
35.219587|564de8f28d0e5500058960b624d49d1bb5607b29|4.99|2014-11-13 21:08:00|80.810069425230125|3|7203695714|401|35.24504930456466|0|23|1647|-80.85013|379|35.175855|PACKAGED MUFFINS|1.5|14|JUMBO PUMPKIN MUFFIN 4 CT.|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00072036959553|MUFFINS|BAKERY|-80.810056|80.810075837400746|218|1
35.219587|7db7b8752c3cc6a0c2336d8e91fbad81f4fcde84|1.19|2015-01-25 19:37:00|80.810069425230125|3|5100001031|401|35.24504930456466|0|23|212|-80.85013|33|35.175855|CONDENSED SOUP|0.0|1|CAMP COND CREAM OF MUSHROOM|54c57a5691b4897585400c0bd735288af5559f5e|1.759384112405368|35.240679762029046|00051000012616|SOUP|G1 GROCERY|-80.810056|80.810075837400746|218|1
35.585842|84c9f484732e3e2c19785d91fbcc8c89d4127374|11.92|2014-10-04 14:49:00|1.4102725052409182|4|20358600000|99|0.6210901099944839|0|1|978|-80.875654|202|35.585842|SMOKED MEATS|0.0|2|SMOKED PORK BUTTS|58508e37fa6d9d07c50484f476cddf589c957580|4.8863766728906|0.61833652052202714|00203586000000|SMOKED HAMS|MEAT|-80.875654|1.411546447003722|99|1
35.585842|b2ccb2a6f5a17a728454da17d7ea954e24e33b96|0.51|2014-12-16 12:15:00|1.4102725052409182|4||99|0.6210901099944839|0|1|502|-80.875654|64|35.585842|FRESH BANANAS|0.0|4|BANANAS, YELLOW|58508e37fa6d9d07c50484f476cddf589c957580|4.8863766728906|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.875654|1.411546447003722|99|1
35.585842|e0a734fb9760521d69fc84d3fff8c60e99a4245d|12.57|2015-02-03 15:25:00|1.4102725052409182|4|76026300010|99|0.6210901099944839|0|1|213|-80.875654|33|35.585842|SOUP MIXES|0.5|1|BEAR CREEK SOUP MIX CHED BROCC|58508e37fa6d9d07c50484f476cddf589c957580|4.8863766728906|0.61833652052202714|00760263000260|SOUP|G1 GROCERY|-80.875654|1.411546447003722|99|3
35.585842|031fc2688b806d333f88bfc8c68e524ed407818e|4.29|2014-11-26 15:17:00|80.891462859624312|4|71514140234|99|35.656559039462145|0|45|364|-80.895009|55|35.603432|ORGANIC AND CF EGGS|0.0|3|EGGLAND'S BEST CAGE FREE JUMBO|58508e37fa6d9d07c50484f476cddf589c957580|4.8863766728906|35.636605227883024|00715141402346|EGGS FRESH|DAIRY|-80.875654|80.875662178412369|274|1
35.585842|faf5ec93964f896a54ef5d90aa3e5213fb055043|17.99|2015-01-16 18:03:00|80.891462859624312|4|7203689916|99|35.656559039462145|0|45|588|-80.895009|136|35.603432|OTHER MERCH FRUIT BASKET|0.0|4|THE SAMPLER FRUIT BASKET|58508e37fa6d9d07c50484f476cddf589c957580|4.8863766728906|35.636605227883024|00072036899163|OTHER MERCHANDISE|PRODUCE|-80.875654|80.875662178412369|274|1
35.585842|ede3d89453542503813aabf98dbc3ff5a1347212|20.5|2015-02-19 10:58:00|80.891462859624312|4|20272300000|99|35.656558970421059|0|45|653|-80.861571|142|35.444615|FRESH VEAL PRIMALS|3.46|2|VEAL LOIN CHOP|58508e37fa6d9d07c50484f476cddf589c957580|4.8863766728906|35.636605227883024|00202723000002|VEAL|MEAT|-80.875654|80.875775837832649|340|2
35.23102|6ec31ccdd56b2fdc6839b57ef3aee6d6e8d3fb45|3.15|2014-09-16 21:30:00|80.843945456961976|2|7265500105|205|35.240053645736076|0|59|1278|-80.810056|48|35.219587|SINGLE SERVE NUTRITIONAL|1.15|5|HC CAFE STEAMERS CHKN MARSALA|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00072655001084|FROZEN MEALS|FROZEN|-80.8438|80.843800376399685|401|1
35.23102|740e08511b83334c120baa39533c14a21364e91d|5.45|2015-02-16 16:01:00|80.843945456961976|2|20328700000|205|35.240053645736076|0|59|641|-80.810056|137|35.219587|PREMIUM PORK|0.0|2|PORK LOIN RIB END CHOPS BNLS|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00203287000002|PORK|MEAT|-80.8438|80.843800376399685|401|1
35.23102|1986e0f08b471db5ec875ad646084345d138767f|6.09|2015-02-22 14:13:00|80.843945456961976|2|20328700000|205|35.240053645736076|0|59|641|-80.810056|137|35.219587|PREMIUM PORK|3.26|2|PORK LOIN RIB END CHOPS BNLS|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00203287000002|PORK|MEAT|-80.8438|80.843800376399685|401|1
35.23102|902dccd52a82b7cb1964f82664956f92680002f0|2.39|2014-12-28 13:45:00|80.843945456961976|2|7203663216|205|35.240053645388251|0|59|330|-80.844274|55|35.204336|EGGS|0.0|3|HT GRADE A    LARGE BROWN EGGS|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00072036632166|EGGS FRESH|DAIRY|-80.8438|80.843803092190811|61|1
35.23102|92ed4e9529de94eb0d94f70837bc1558c09d37eb|1.59|2014-11-16 17:15:00|1.4094857484078087|2|4280011400|205|0.6148972978359727|0|26|255|-80.8438|892|35.23102|VALUE PIZZA|0.59|5|TOTINO'S CHEESE PIZZA|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|0.61471665291522548|00042800113009|FROZEN PIZZA|FROZEN|-80.8438|1.4109904898237917|205|1
35.23102|810bea5d024b290eea4a4a05f74534bb05d4e139|1.29|2015-02-18 11:18:00|1.4094857484078087|2|7203657030|205|0.6148972978359727|0|26|322|-80.8438|53|35.23102|SOUR CREAM|0.49|3|HT LIGHT SOUR CREAM|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|0.61471665291522548|00072036600349|CULTURES|DAIRY|-80.8438|1.4109904898237917|205|1
35.23102|5c45b61a2c43c6965165fd516c1df82a0b14096d|1.97|2014-11-26 18:25:00|1.4094857484078087|2|7203656065|205|0.6148972978359727|0|26|315|-80.8438|52|35.23102|CHEESE-PROCESSED-SLICED|0.0|3|HT SINGLE WRAP CHEESE|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|0.61471665291522548|00072036560650|CHEESE|DAIRY|-80.8438|1.4109904898237917|205|1
35.23102|6da64374eb95d0c09af3b51edcc8e3d2676bea8d|2.97|2014-10-10 22:30:00|80.843945456961976|2|7203658035|205|35.240053645736076|0|59|358|-80.810056|100|35.219587|REGULAR BACON|0.0|19|HT REGULAR SLICED BACON|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00072036580351|BACON|CASE READY MEATS|-80.8438|80.843800376399685|401|1
35.23102|4a9b28c66e87596525219b54cf758e9bb230466e|1.69|2014-10-19 14:05:00|80.843945456961976|2|4600083251|205|35.240053645736076|0|59|1212|-80.810056|272|35.219587|HISP BEANS/PEPPERS|0.0|1|OEP CHILIES GREEN CHOPPED|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00046000832517|HISPANIC PREP. FOODS|G1 GROCERY|-80.8438|80.843800376399685|401|1
35.23102|3ddec9eb25e313b64ee04a97213eef98be5e0743|3.49|2014-11-02 10:11:00|1.4094857484078087|2|4812127620|205|0.6148972978359727|0|26|1037|-80.8438|164|35.23102|ENGLISH MUFFINS|1.74|7|THOMAS PUMPKIN EM PP|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|0.61471665291522548|00048121184193|BREAKFAST|COMMERCIAL BAKERY|-80.8438|1.4109904898237917|205|1
35.23102|a52593ed449140f116d6c0010e8e7f01159d2a0d|2.4|2014-09-25 19:06:00|80.843945456961976|2|3663202717|205|35.240053645736076|0|59|685|-80.810056|61|35.219587|GREEK|0.0|3|DANNON OIKOS KEY LIME TRAD|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00036632032218|YOGURT|DAIRY|-80.8438|80.843800376399685|401|2
35.23102|8135db9b29ae8bce537b6b6433fe857db7a5157e|5.59|2015-01-05 17:58:00|80.843945456961976|2|3700047451|205|35.240053645736076|0|59|4092|-80.810056|1080|35.219587|TOOTHPASTE-WHITENING|1.6|17|CREST 3D WH GLMRS VIBR MINT TP|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00037000891918|ORAL HYGIENE|HBC|-80.8438|80.843800376399685|401|1
35.23102|6f028115d1b16fb6d081a83b5c389a707da9cca9|10.36|2014-09-29 20:02:00|80.843945456961976|2|8000051306|205|35.240053645736076|0|59|189|-80.810056|29|35.219587|TUNA-POUCH|5.36|1|STARKIST TUNA PCH LS CHNK LGHT|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00080000505279|SEAFOOD-CANNED|G1 GROCERY|-80.8438|80.843800376399685|401|4
35.23102|ab8e9bbfbbd8095feb398d8711c2d4d079c279ff|5.04|2015-02-09 16:14:00|80.843945456961976|2|20337700000|205|35.240053645736076|0|59|641|-80.810056|137|35.219587|PREMIUM PORK|0.0|2|PORK LOIN CHOPS BNLS THIN|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00203377000004|PORK|MEAT|-80.8438|80.843800376399685|401|1
35.23102|1f5b1e47d8de35e0ad0742b15bf557bf547cb46d|4.65|2014-12-01 19:39:00|80.843945456961976|2|8000051306|205|35.240053645736076|0|59|189|-80.810056|29|35.219587|TUNA-POUCH|0.8999999999999999|1|STARKIST TUNA PCH LS CHNK LGHT|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00080000505279|SEAFOOD-CANNED|G1 GROCERY|-80.8438|80.843800376399685|401|3
35.23102|b323bc60ff4acbfdf0fbde10dda06352e6e9c45a|3.97|2014-11-01 21:40:00|1.4094857484078087|2|7203659020|205|0.6148972978359727|0|26|312|-80.8438|51|35.23102|BUTTER|0.0|3|HARRIS TEETER UNSALTED BUTTER|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|0.61471665291522548|00072036590213|BUTTER & MARGARINE|DAIRY|-80.8438|1.4109904898237917|205|1
35.23102|55b92ddec1e91a5249aaffd49ea406dc44135825|3.35|2014-10-07 16:33:00|80.843945456961976|2|7203656080|205|35.240053645736076|0|59|318|-80.810056|52|35.219587|SHREDDED/GRATED CHEESE|0.0|3|HT FANCY SHRED MILD CHED CHES|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00072036560810|CHEESE|DAIRY|-80.8438|80.843800376399685|401|1
35.23102|12433fa4087728bdb089d5406d94af1381310054|3.55|2015-02-02 20:09:00|80.843945456961976|2||205|35.240053645736076|0|59|505|-80.810056|64|35.219587|FRESH SOFT FRUIT|0.89|4|NECTARINES,TREE RIPE, XL|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00204378000000|FRESH PRODUCE|PRODUCE|-80.8438|80.843800376399685|401|1
35.23102|3729bfcea7137cad87ecf73fa0b38649ad61149d|12.95|2014-12-19 18:43:00|80.843945456961976|2|20138900000|205|35.240053645736076|0|59|296|-80.810056|49|35.219587|RANCHER BEEF|3.6|2|BEEF TENDERLOIN FILET MIGNON|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00201389000005|BEEF|MEAT|-80.8438|80.843800376399685|401|1
35.23102|38b56b8dbf2da99c2573dfc20a3d74f46f99aed1|2.59|2015-02-06 19:27:00|80.843945456961976|2||205|35.240053645736076|0|59|505|-80.810056|64|35.219587|FRESH SOFT FRUIT|0.97|4|NECTARINES,TREE RIPE, XL|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00204378000000|FRESH PRODUCE|PRODUCE|-80.8438|80.843800376399685|401|1
35.23102|3d4f127db0c152aaba12dade5a743c04bdd13dba|4.65|2014-09-12 06:26:00|80.843945456961976|2|97151|205|35.240053645736076|0|59|1589|-80.810056|369|35.219587|NFS BEVERAGE ESPRESSO|0.0|22|PUMPKIN SPICE LATTE GRANDE|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00000000971510|NFS STARBUCKS|COFFEE SHOP|-80.8438|80.843800376399685|401|1
35.23102|698830448656257b809c8088feec727518aa6901|1.79|2014-11-25 20:01:00|80.843945456961976|2|1200000157|205|35.240053645736076|0|59|31|-80.810056|4|35.219587|NON CARBONATED WATER|0.79|1|AQUAFINA WATER  1 LITER|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00012000001574|BOTTLED WATER|G1 GROCERY|-80.8438|80.843800376399685|401|1
35.23102|4e668d339e8f7effd39aad5684ef4857de31567a|7.79|2015-01-17 13:41:00|80.843945456961976|2|30045027125|205|35.240053645736076|0|59|4236|-80.810056|1200|35.219587|DEX ADULT/CHILDREN|1.8|17|TYL SEVERE COLD/FLU CAPLETS|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00300450270269|COUGH/COLD/SINUS|HBC|-80.8438|80.843800376399685|401|1
35.23102|6dda07a28bc34df3fcab226f47ed8d5ac11befa0|2.19|2014-09-13 16:20:00|80.843945456961976|2|7203670268|205|35.240053645388251|0|59|176|-80.844274|72|35.204336|NFS-DISPOSE CUPS|0.0|1|YH PLASTIC CUPS 18OZ|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00072036702685|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.8438|80.843803092190811|61|1
35.23102|c5d66d317df5bf32511b8d48e2cca0a2a6644e08|7.99|2015-02-07 16:22:00|80.843945456961976|2|8500000715|205|35.240053635406703|0|59|9983|-80.764523|889|35.341927|NFS-SPARKLING|0.0|13|TOTT'S BRUT|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00085000007150|SPARKLING|WINE|-80.8438|80.843816729561524|220|1
35.23102|c0f73971fb52b1e1fa67d823b0e906e155b97fcb|3.25|2015-01-29 20:18:00|80.843945456961976|2|4157005617|205|35.240053645736076|0|59|1265|-80.810056|57|35.219587|ALMOND MILK|0.0|3|ALMOND BREEZE UNSWEETENED VAN|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00041570056189|MILK|DAIRY|-80.8438|80.843800376399685|401|1
35.23102|3d6de398c0c4914e9c9313055d87c0d3c607a3ba|1.55|2015-01-19 17:27:00|80.843945456961976|2|78616201000|205|35.240053624559991|0|59|31|-80.847383|4|35.024464|NON CARBONATED WATER|0.55|1|VIT WATER ESSENTIAL 20 OZ|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00786162040008|BOTTLED WATER|G1 GROCERY|-80.8438|80.843823950459651|317|1
35.23102|ab65b34e09d96842c3248e2327784f0d700e974d|3.19|2014-10-19 13:24:00|1.4094857484078087|2|1800081778|205|0.6148972978359727|0|26|326|-80.8438|54|35.23102|COOKIES/BROWNIES-REFRIGERATED|0.69|3|PILLSURY RTB SUGAR|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|0.61471665291522548|00018000817726|DOUGH PRODUCTS|DAIRY|-80.8438|1.4109904898237917|205|1
35.23102|deb50f2b12083a379aeadb68216d50128d31733b|7.19|2015-01-14 20:11:00|80.843945456961976|2|20253500000|205|35.240053645736076|0|59|299|-80.810056|49|35.219587|ANGUS BEEF|0.0|2|ANGUS BEEF SIRLOIN STIR FRY|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00202533000001|BEEF|MEAT|-80.8438|80.843800376399685|401|1
35.23102|6b45d475f71f15c522b5d2fc2c504134b69e7a81|3.15|2014-11-18 16:05:00|80.843945456961976|2|7265500105|205|35.240053645736076|0|59|1278|-80.810056|48|35.219587|SINGLE SERVE NUTRITIONAL|0.0|5|HC CAFE STEAMER SWTSPC ORN CHK|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00072655001091|FROZEN MEALS|FROZEN|-80.8438|80.843800376399685|401|1
35.23102|1801bb32edd4a4f2364ef07c1c24e989b0900016|21.99|2015-02-13 16:35:00|80.843945456961976|2|20310200000|205|35.240053645736076|0|59|1153|-80.810056|87|35.219587|NFS-FRESH CUT ARRANGE|0.0|9|*ROSE ARRANGEMENTS|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00203102000002|FLORAL|FLORAL|-80.8438|80.843800376399685|401|1
35.23102|c716923b02bc282091c7bdb4cd964bcd7e280ad5|13.49|2014-10-13 21:13:00|80.843945456961976|2|89445500031|205|35.240053645736076|0|59|1435|-80.810056|19|35.219587|SHELF STABLE SPREADS|0.0|1|JUSTINS VANILLA ALMOND BUTTER|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00894455000377|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.8438|80.843800376399685|401|1
35.23102|8523b2f81c16ef0698e5fb40d46c5f5d75dfba82|1.99|2014-10-30 17:45:00|1.4094857484078087|2|7203648011|205|0.6148972978359727|0|26|274|-80.8438|44|35.23102|ICE|0.0|5|HT BAGGED ICE 10LB (456)|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|0.61471665291522548|00000000004560|ICE|FROZEN|-80.8438|1.4109904898237917|205|1
35.23102|0d1d78513e84d4ebe24e28416fdb60ad80a3d3dd|5.49|2015-02-14 19:43:00|80.843945456961976|2|7895150058|205|35.240053645736076|0|59|533|-80.810056|64|35.219587|FRESH PEPPERS|0.0|4|STOPLIGHT PEPPER 3PK|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00078951500580|FRESH PRODUCE|PRODUCE|-80.8438|80.843800376399685|401|1
35.23102|0eb4b8a6c07c1e3c105143e45d135d48454f582d|9.99|2014-11-01 18:39:00|80.843945456961976|2|8500002157|205|35.240053635406703|0|59|9979|-80.764523|888|35.341927|NFS-U/PREM-MALBEC|0.0|13|BAREFOOT MALBEC 1.5L|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00085000021576|ULTRA PREMIUM ($15-$19.99)|WINE|-80.8438|80.843816729561524|220|1
35.23102|40a24653a5e1d7d47b7a3b67d171a4ac8ea7715e|1.05|2014-10-28 16:15:00|80.843945456961976|2||205|35.240053645736076|0|59|502|-80.810056|64|35.219587|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00204011000008|FRESH PRODUCE|PRODUCE|-80.8438|80.843800376399685|401|1
35.23102|a293a15f7b9283e8ac984bf10287a3129d01341d|0.2|2015-03-06 06:37:00|80.843945456961976|2||205|35.240053645736076|0|59|502|-80.810056|64|35.219587|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00204011000008|FRESH PRODUCE|PRODUCE|-80.8438|80.843800376399685|401|1
35.23102|6923cc5d4519df3d533364221636c958aa0cad28|3.39|2014-12-11 20:40:00|80.843945456961976|2|3680013316|205|35.240053645736076|0|59|4418|-80.810056|1210|35.219587|ANTINAUSEA REMEDY-LIQUID|0.0|17|TC REG STR PEPTIC RELIEF-CHRRY|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00036800133167|STOMACH REMEDIES|HBC|-80.8438|80.843800376399685|401|1
35.23102|62c7f088667f4a8f83487e42d4968f20621f88c7|1.4|2015-02-11 17:51:00|80.843945456961976|2||205|35.240053624559991|0|59|501|-80.847383|64|35.024464|FRESH PEARS|0.16|4|ANJOU PEARS|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00204416000009|FRESH PRODUCE|PRODUCE|-80.8438|80.843823950459651|317|1
35.23102|13aab1885d9a67e12f9a8e73eeffa3771dbc449d|7.99|2014-09-13 16:19:00|80.843945456961976|2|32390001424|205|35.240053645388251|0|59|4236|-80.844274|1200|35.204336|DEX ADULT/CHILDREN|1.5|17|NYQUIL LIQUICAP|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00323900014398|COUGH/COLD/SINUS|HBC|-80.8438|80.843803092190811|61|1
35.23102|a4be63ff50cd6b4e0a409a99f258ce34c079dfaf|3.99|2015-01-14 06:31:00|80.843945456961976|2|7203695459|205|35.240053645736076|0|59|2003|-80.810056|495|35.219587|FFM GREEN SALADS|1.0|6|NEW CAESAR  W/CRTNS|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00072036954596|GREEN SALADS|DELI|-80.8438|80.843800376399685|401|1
35.23102|8163543d459dbbcdaa3b6b25657f4b0c598bf8c0|1.99|2015-01-08 16:44:00|80.843945456961976|2|1780054108|205|35.240053645736076|0|59|168|-80.810056|24|35.219587|NFS-CAT TREATS|0.0|1|WHISKER LICKIN MOUSERS TREATS|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00017800541084|PET FOOD/SUPPLIES|G1 GROCERY|-80.8438|80.843800376399685|401|1
35.23102|e617c58f4350c47bc317432b0a812ba7b0c6b0bd|1.44|2015-02-09 12:17:00|80.843945456961976|2||205|35.240053645388251|0|59|505|-80.844274|64|35.204336|FRESH SOFT FRUIT|0.0|4|RED PLUMS|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00204042000008|FRESH PRODUCE|PRODUCE|-80.8438|80.843803092190811|61|1
35.23102|fed60c8c36ada97b9d125964b15ce0f77d21ba8a|14.99|2015-01-24 22:09:00|80.843945456961976|2|1820053168|205|35.240053645736076|0|59|455|-80.810056|82|35.219587|DOMESTIC PREMIUM 12PK&>|0.0|16|BUD LIGHT 24PK 12OZ CANS|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00018200531682|DOMESTIC BEER|BEER|-80.8438|80.843800376399685|401|1
35.23102|13254d16b0a14d3fa7d365127342b116e8135294|3.99|2015-02-02 17:16:00|80.843945456961976|2|72243011016|205|35.240053624559991|0|59|577|-80.847383|136|35.024464|OTHER MERCH FR MSC JUICE|0.0|4|ORG. GT KOMBUCHA CRANBERRY|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00722430300160|OTHER MERCHANDISE|PRODUCE|-80.8438|80.843823950459651|317|1
35.23102|344db440bad28b5be3c42bbb14b77a22e6551cd1|6.99|2015-02-04 20:06:00|80.843945456961976|2|4242122579|205|35.240053645736076|0|59|358|-80.810056|100|35.219587|REGULAR BACON|1.0|19|BOARS HEAD SMOKED BACON 16 OZ|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00042421225792|BACON|CASE READY MEATS|-80.8438|80.843800376399685|401|1
35.23102|5b1136e7bd048307f00dfa4fe90b06af03faa590|2.35|2015-01-22 06:36:00|80.843945456961976|2||205|35.240053645736076|0|59|562|-80.810056|64|35.219587|FRESH CUT FRUIT|0.0|4|CANTALOUPE CHUNKS (IN-STORE)|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00204318000008|FRESH PRODUCE|PRODUCE|-80.8438|80.843800376399685|401|1
35.23102|9f73a3bc6fee314bc15b55b00ea595f076f83c1d|8.99|2014-12-24 18:14:00|80.843945456961976|2|85337000208|205|35.240053635406703|0|59|458|-80.764523|82|35.341927|CRAFT BEER|0.0|16|LONERIDER SWEET JOSIE 24/12|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00853370002088|DOMESTIC BEER|BEER|-80.8438|80.843816729561524|220|1
35.23102|13738639e39392f8991afdc480b338f8a63c5211|4.15|2014-10-03 06:22:00|80.843945456961976|2|97158|205|35.240053645736076|0|59|1589|-80.810056|369|35.219587|NFS BEVERAGE ESPRESSO|0.0|22|VANILLA LATTE GRANDE|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00000000971580|NFS STARBUCKS|COFFEE SHOP|-80.8438|80.843800376399685|401|1
35.23102|7b822eb71abe8303ed4b347f86cd41a0964132c6|4.15|2014-10-10 06:27:00|80.843945456961976|2|97158|205|35.240053645736076|0|59|1589|-80.810056|369|35.219587|NFS BEVERAGE ESPRESSO|0.0|22|VANILLA LATTE GRANDE|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00000000971580|NFS STARBUCKS|COFFEE SHOP|-80.8438|80.843800376399685|401|1
35.23102|9eeb6eb8bb03c16300700c578b15a476caa2ce45|9.99|2014-11-30 12:11:00|80.843945456961976|2|7203678030|205|35.240053645736076|0|59|458|-80.810056|82|35.219587|CRAFT BEER|0.0|16|HT CREATE YOUR OWN SAMPLER|5960cd72b65f296f250fabd676c633d584ec7957|0.6242031052505824|35.232478750868765|00072036780300|DOMESTIC BEER|BEER|-80.8438|80.843800376399685|401|1
35.17335|41c9e7eb1f54c422f3db293656b56b77049e42de|4.59|2014-10-16 16:43:00|80.709059419360486|3|2700061286|174|35.186342437510824|0|31|195|-80.709466|30|35.124987|SALAD & COOKING OIL|1.09|1|WESSON VEGETABLE OIL|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00027000612866|SHORTENING/OIL|G1 GROCERY|-80.70901|80.709018040149374|157|1
35.17335|ed45da41b0c0656aff2151c048476d5d74ec402b|1.89|2014-11-20 14:18:00|1.4094857484078087|3|2000000065|174|0.6138907664563474|0|26|1272|-80.70901|50|35.17335|BAG VEG STEAM|0.89|5|GG BOIL IN BAG ROSEMARY|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|0.61471665291522548|00020000481821|VEGETABLES-FROZEN|FROZEN|-80.70901|1.4086379605250285|174|1
35.17335|298ec7cc610010035149d7a532156c4dcfc2dc7b|3.78|2014-12-18 15:23:00|1.4094857484078087|3|2000000065|174|0.6138907664563474|0|26|1272|-80.70901|50|35.17335|BAG VEG STEAM|1.78|5|GG BOIL IN BAG ROSEMARY|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|0.61471665291522548|00020000481821|VEGETABLES-FROZEN|FROZEN|-80.70901|1.4086379605250285|174|2
35.17335|80df9fe608ba65e6e079279357416ece8a832e75|3.29|2014-12-30 12:31:00|1.4094857484078087|3|2840004768|174|0.6138907664563474|0|26|202|-80.70901|31|35.17335|PRETZELS|0.79|1|ROLD GOLD 3 CHEESE PRETZEL THN|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|0.61471665291522548|00028400232043|SNACKS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|4e2b22c227b212cd400849b1ee0ce18aaf932178|4.29|2015-02-05 17:47:00|80.709059419360486|3|2840015636|174|35.186342438884516|0|31|204|-80.661096|31|35.172688|TORTILLA CHIPS|1.79|1|DORTIOS NACHO CHEESE|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00028400156363|SNACKS|G1 GROCERY|-80.70901|80.709013348554933|474|1
35.17335|d7db1ddc50749184e06af7a3cf205bd2cf82c008|3.49|2014-09-15 15:59:00|1.4094857484078087|3|1410007438|174|0.6138907664563474|0|26|1253|-80.70901|12|35.17335|ALL OTHER COOKIES|1.75|1|PF SWEET SIMPLE SHORTBREAD|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|0.61471665291522548|00014100074441|COOKIES|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|a9a90a1929562515144b18e1dae2f18063fc461e|3.49|2014-09-13 15:58:00|1.4094857484078087|3|1410007438|174|0.6138907664563474|0|26|1253|-80.70901|12|35.17335|ALL OTHER COOKIES|1.75|1|PF SWEET SIMPLE SHORTBREAD|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|0.61471665291522548|00014100074441|COOKIES|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|c4fd09e8ade5467a4df5e5b47ebab2346114f73b|3.25|2015-01-15 16:01:00|1.4094857484078087|3|7203656080|174|0.6138907664563474|0|26|318|-80.70901|52|35.17335|SHREDDED/GRATED CHEESE|1.58|3|HT SHREDDED COLBY JACK|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|0.61471665291522548|00072036600745|CHEESE|DAIRY|-80.70901|1.4086379605250285|174|1
35.17335|cb5fa4d5bbfbd830236923ec4caf96a5b8b924f5|3.35|2014-10-23 15:12:00|80.709059419360486|3|7203656080|174|35.186342437510824|0|31|318|-80.709466|52|35.124987|SHREDDED/GRATED CHEESE|1.68|3|HT SHREDDED COLBY JACK|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00072036600745|CHEESE|DAIRY|-80.70901|80.709018040149374|157|1
35.17335|872f63f8efa81ef28e845975e13e05425e1c59ae|2.79|2015-02-19 13:18:00|1.4094857484078087|3|7203670356|174|0.6138907664563474|0|26|442|-80.70901|76|35.17335|NFS-COOKING-STORAGE BAGS|0.82|1|YH FREEZER BAGS QUART 20CT|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|0.61471665291522548|00072036703576|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|627a535af2a7ca60b6ebd86255227517dc7730ad|2.0|2014-10-05 11:59:00|1.4094857484078087|3|7203663118|174|0.6138907664563474|0|26|1262|-80.70901|57|35.17335|HALF N HALF WHIPPING CREAM|0.0|3|HT HALF & HALF|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|0.61471665291522548|00072036632043|MILK|DAIRY|-80.70901|1.4086379605250285|174|1
35.17335|8034859f67b9e7ca19478d394a4f560a65a3ecde|2.99|2014-09-18 17:01:00|80.709059419360486|3|7203670673|174|35.186342438884516|0|31|205|-80.661096|31|35.172688|REMAINING SNACKS|0.49|1|HTT SOCRISP PITA CHIPS RANCH|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00072036706744|SNACKS|G1 GROCERY|-80.70901|80.709013348554933|474|1
35.17335|ed947e868edd3df62757db3a7835bfb9eaaaf636|2.89|2015-03-07 15:07:00|80.709059419360486|3|7203655029|174|35.186342437510824|0|31|331|-80.709466|52|35.124987|NATURAL SLICED|0.92|3|HT PROVOLONE SLICES|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00072036550170|CHEESE|DAIRY|-80.70901|80.709018040149374|157|1
35.17335|84bd31c6280ad1594510d79a44bbbc3ff6114da9|2.0|2014-11-08 19:44:00|1.4094857484078087|3|7203663118|174|0.6138907664563474|0|26|1262|-80.70901|57|35.17335|HALF N HALF WHIPPING CREAM|0.0|3|HT HALF & HALF|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|0.61471665291522548|00072036632043|MILK|DAIRY|-80.70901|1.4086379605250285|174|1
35.17335|f87c8d568b31329f8c985e341b0f8229543bb9da|3.99|2015-01-22 18:07:00|80.709059419360486|3|7203604217|174|35.186342438884516|0|31|275|-80.661096|45|35.172688|SUPER PREMIUM ICE CREAM|0.0|5|HTT DBLE COCNT ALMD ICE CREAM|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00072036709189|ICE CREAM|FROZEN|-80.70901|80.709013348554933|474|1
35.17335|11066515e4c26e5827a534c73db4a334015bf70a|3.25|2014-11-13 13:40:00|80.709059419360486|3|7203656080|174|35.186342437510824|0|31|318|-80.709466|52|35.124987|SHREDDED/GRATED CHEESE|3.25|3|HT SHREDDED MOZZ/PROVLONE|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00072036705174|CHEESE|DAIRY|-80.70901|80.709018040149374|157|1
35.17335|e0a2ee2f4ce3bf8543dae97e8521c5e3fe86c03a|5.49|2015-02-28 18:19:00|1.4094857484078087|3|7597140209|174|0.6138907664563474|0|26|1845|-80.70901|425|35.17335|FFM PRESLICED CHEESE|0.0|6|F.F. SMOKED PROVOLONE CHEESE|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|0.61471665291522548|00072036010360|PRESLICED CHEESE|DELI|-80.70901|1.4086379605250285|174|1
35.17335|649ddddc57e3ac02bb25c95a4ec833f5090185a4|1.99|2015-02-05 17:41:00|80.709059419360486|3|7203603105|174|35.186342438884516|0|31|757|-80.661096|3|35.172688|BAKING NUTS|0.32|1|HT WALNUT PIECES|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00072036031051|BAKING SUPPLIES|G1 GROCERY|-80.70901|80.709013348554933|474|1
35.17335|a6666ff36c8d566e1ddbcf6f1505d05656be7b18|3.35|2014-10-23 15:14:00|80.709059419360486|3|7203656080|174|35.186342437510824|0|31|318|-80.709466|52|35.124987|SHREDDED/GRATED CHEESE|1.67|3|HT GOURMENT SHARP BLEND|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00072036600783|CHEESE|DAIRY|-80.70901|80.709018040149374|157|1
35.17335|5575bf819a693cf0562c61a06ee239452ff5426e|5.78|2014-12-26 18:33:00|80.709059419360486|3|7203655029|174|35.18634243773306|0|31|331|-80.739|52|35.141204|NATURAL SLICED|1.22|3|HT SLICED MUENSTER CHEESE|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00072036600387|CHEESE|DAIRY|-80.70901|80.709017483322825|171|2
35.17335|3742767cf21bae70843545c1f6b7cddbdf75c79e|2.65|2015-01-10 10:11:00|80.709059419360486|3|4119691401|174|35.18634243773306|0|31|1201|-80.739|33|35.141204|RTS CANNED|0.0|1|PROG RICH HRT CHCKEN WILD RICE|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00041196453850|SOUP|G1 GROCERY|-80.70901|80.709017483322825|171|1
35.17335|15cb9782e198e3d7e59713840effa3b506889ebe|1.89|2014-11-22 17:23:00|80.709059419360486|3|2000000065|174|35.18634243773306|0|31|1275|-80.739|50|35.141204|BOX VEG|0.89|5|GG BROCCOLI SPEAR NO SAUCE|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00020000174839|VEGETABLES-FROZEN|FROZEN|-80.70901|80.709017483322825|171|1
35.17335|7051cb1b72c9fafa716829eaeb7740aa8846f016|1.95|2014-10-18 15:45:00|80.709059419360486|3|2000000065|174|35.186342430473871|0|31|1275|-80.737839|50|35.297134|BOX VEG|0.28|5|GG SPINACH NO SAUCE|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00020000176819|VEGETABLES-FROZEN|FROZEN|-80.70901|80.709028394415171|258|1
35.17335|f4f7331fb301d22b8c63966d315f1d066611bfcb|3.49|2015-01-17 16:28:00|1.4094857484078087|3|2840023981|174|0.6138907664563474|0|26|203|-80.70901|31|35.17335|CHEESE SNACKS|1.75|1|CHEETOS MIX UPS XXTRA CHEESY|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|0.61471665291522548|00028400240123|SNACKS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|d3c7cfbf2cdf58a5caaf250747d3883727fa6893|4.29|2015-01-30 16:39:00|80.709059419360486|3|84357100478|174|35.186342438708223|0|31|197|-80.654118|31|35.123768|POPPED POPCORN|1.3|1|POP IND KETTLE CORN|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00843571004707|SNACKS|G1 GROCERY|-80.70901|80.709014250856526|473|1
35.17335|9641e3ee9e0cad16906d98582e9de8f18c5a88ff|8.58|2014-12-05 11:09:00|1.4094857484078087|3|84357100478|174|0.6138907664563474|0|26|197|-80.70901|31|35.17335|POPPED POPCORN|3.58|1|POP IND KETTLE CORN|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|0.61471665291522548|00843571004707|SNACKS|G1 GROCERY|-80.70901|1.4086379605250285|174|2
35.17335|19cd4e55d8175496a62ee84e182dbf7d83452c27|3.65|2015-03-04 13:14:00|80.709059419360486|3|3010067264|174|35.186342418414036|0|31|91|-80.760919|13|35.024332|SPRAYED BUTTER CRACKERS|1.15|1|KEEBLER TOWN HOUSE ORIGINAL|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00030100100553|CRACKERS|G1 GROCERY|-80.70901|80.709038415414284|343|1
35.17335|92fd4b7e0ce34ca1ac3f75f4f519aa78e8cad745|3.65|2014-11-29 16:01:00|1.4094857484078087|3|3010067264|174|0.6138907664563474|0|26|91|-80.70901|13|35.17335|SPRAYED BUTTER CRACKERS|1.15|1|TOWN HOUSE PRETZEL THINS PARMS|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|0.61471665291522548|00030100102335|CRACKERS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|e1c631656f2fe695b5af577af21f0b878cc8a4ef|2.69|2014-10-09 14:47:00|80.709059419360486|3|70935100013|174|35.186342437510824|0|31|556|-80.709466|64|35.124987|PACKAGED VEGETABLES|0.69|4|APIO BROCCOLI & CAULIFLOWER|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00709351000263|FRESH PRODUCE|PRODUCE|-80.70901|80.709018040149374|157|1
35.17335|50b7222944a76761136aba6eb696cd369e925403|2.69|2014-12-24 15:39:00|80.709059419360486|3|70935100013|174|35.18634243773306|0|31|556|-80.739|64|35.141204|PACKAGED VEGETABLES|0.19|4|APIO BROCCOLI & CAULIFLOWER|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00709351000263|FRESH PRODUCE|PRODUCE|-80.70901|80.709017483322825|171|1
35.17335|07cba93dd2e7c5f1627d40498f661efc96ed501a|3.0|2014-10-02 17:15:00|80.709059419360486|3|20600200000|174|35.186342438884516|0|31|1802|-80.661096|400|35.172688|FFM HAM|1.5|6|HONEY CURED HAM|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00206002000004|FFM MEAT|DELI|-80.70901|80.709013348554933|474|1
35.17335|9ecce4b426d8a6dfb9d9bc0c8d5ba6bd6b4d0d6c|19.98|2014-12-20 18:20:00|1.4094857484078087|3|4200044517|174|0.6138907664563474|0|26|426|-80.70901|72|35.17335|NFS-PAPER TOWELS|6.0|1|BRAWNY 6 BIG ROLL PICK A SIZE|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|0.61471665291522548|00042000445177|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.70901|1.4086379605250285|174|2
35.17335|012dd65ff00d3aab83cc06cf92b07928e73cbc48|9.94|2014-09-20 13:52:00|80.709059419360486|3|4200044517|174|35.186342438884516|0|31|426|-80.661096|72|35.172688|NFS-PAPER TOWELS|0.0|1|BRAWNY 6 BIG ROLL PICK A SIZE|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00042000445177|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.70901|80.709013348554933|474|2
35.17335|1142889b47de1fed1f9339c8d22ab8c1d25259f7|17.98|2014-10-18 14:43:00|80.709059419360486|3|4300005001|174|35.186342429992663|0|31|37|-80.780702|10|35.318911|PODS/CUPS/SINGLES|4.0|1|GEVALIA DRK ROYAL ROAST K PODS|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00043000049921|COFFEE|G1 GROCERY|-80.70901|80.70902889634543|167|2
35.17335|128d255ba3114f14df26fbca50d69ad747217b1a|4.38|2015-03-08 12:35:00|80.709059419360486|3|4800000086|174|35.186342431957513|0|31|187|-80.7007|29|35.06858|SALMON-CANNED|1.38|1|COS PINK SALMON SB|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00048000000866|SEAFOOD-CANNED|G1 GROCERY|-80.70901|80.709026752513196|273|2
35.17335|f60f312db488f47452397ed8ce87c7cf6ca13f70|3.65|2014-11-06 13:16:00|1.4094857484078087|3|4610000094|174|0.6138907664563474|0|26|318|-80.70901|52|35.17335|SHREDDED/GRATED CHEESE|1.15|3|SARGENTO CB 6 CHEESE ITALIAN|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|0.61471665291522548|00046100000915|CHEESE|DAIRY|-80.70901|1.4086379605250285|174|1
35.17335|62b46e753cc1da5ee5a8159f6c8cecb1188f00c8|0.83|2014-10-16 16:48:00|80.709059419360486|3||174|35.186342437510824|0|31|565|-80.709466|64|35.124987|REDUCED PRODUCE|0.0|4|PRODUCE REWRAP BY LB|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00204844000008|FRESH PRODUCE|PRODUCE|-80.70901|80.709018040149374|157|1
35.17335|7847857efc4a335bed2337f3b9daf7f9bbfc87cd|2.98|2015-01-24 22:19:00|80.709059419360486|3||174|35.186342430473871|0|31|565|-80.737839|64|35.297134|REDUCED PRODUCE|0.0|4|PRODUCE REWRAP BY CT|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00204845000007|FRESH PRODUCE|PRODUCE|-80.70901|80.709028394415171|258|2
35.17335|6f436e9010278d5db8f6b4c46c2196c40fb1dc9a|1.0|2015-01-24 20:19:00|80.709059419360486|3||174|35.186342424526778|0|31|565|-80.764523|64|35.341927|REDUCED PRODUCE|0.0|4|PRODUCE REWRAP BY CT|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00204845000007|FRESH PRODUCE|PRODUCE|-80.70901|80.709033867836567|220|1
35.17335|721b39409f2698b5b49cdce0334ae2aba0002b31|4.98|2015-03-08 11:59:00|80.709059419360486|3|4150880012|174|35.18634243215002|0|31|30|-80.64817|4|35.04711|CARBONATED WATER|0.98|1|SAN PELLEGRINO 750ML|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00041508800129|BOTTLED WATER|G1 GROCERY|-80.70901|80.709026527519597|129|2
35.17335|69e3d3e7654725018da78168ca8a4546017ca406|5.19|2015-01-27 15:35:00|80.709059419360486|3|7274500224|174|35.186342438884516|0|31|1224|-80.661096|107|35.172688|CHICKEN STRIPS|2.59|19|PERDUE SHORTCUTS HONEY ROASTD|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00072745002243|HEAT & EAT|CASE READY MEATS|-80.70901|80.709013348554933|474|1
35.17335|12c333b01b7ecab68121ecf6bfa1095b228fbb77|4.19|2015-03-08 11:18:00|80.709059419360486|3|73291322811|174|35.186342431612339|0|31|398|-80.562829|69|35.006282|NFS-BATHROOM CLEANERS|0.0|1|7TH GEN DISINFECT BATHRM CLNR|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00732913228119|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.70901|80.709027148551911|60|1
35.17335|5ffcf52875f770e56b7878af0b26c344577ea4f1|28.97|2014-10-18 14:09:00|80.709059419360486|3|78535701280|174|35.186342424526778|0|31|37|-80.764523|10|35.341927|PODS/CUPS/SINGLES|8.0|1|PEET'S 10CT HOUSE BLEND|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00785357012592|COFFEE|G1 GROCERY|-80.70901|80.709033867836567|220|3
35.17335|132a2138913040d47e2eac9ccbbd78f3980b2449|0.5|2014-10-02 17:16:00|80.709059419360486|3|7203698487|174|35.186342438884516|0|31|201|-80.661096|31|35.172688|POTATO CHIPS|0.0|1|HT ORIGINAL POTATO CHIPS|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00072036984876|SNACKS|G1 GROCERY|-80.70901|80.709013348554933|474|1
35.17335|41f017709f84e356999c4e56e204258c3a9477a9|3.23|2015-01-21 13:41:00|80.709059419360486|3|7726006141|174|35.186342424526778|0|31|727|-80.764523|7|35.341927|SEASONAL CANDY-SINGLE FAC|0.0|1|I/O(C15)RS DC RED VELVET SANTA|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00077260061416|CANDY|G1 GROCERY|-80.70901|80.709033867836567|220|3
35.17335|7af4e0181feb9e5540cb5f84c28fe743581ae186|3.39|2014-10-16 16:50:00|80.709059419360486|3|4450034122|174|35.186342437510824|0|31|357|-80.709466|104|35.124987|SMOKED SAUSAGE ROPES|1.45|19|HILLSHIRE POLSKA KIELBASA|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00044500341225|DINNER SAUSAGE|CASE READY MEATS|-80.70901|80.709018040149374|157|1
35.17335|fcf758534a57a2dabd6de55cf9dfb30aa96f4c09|2.29|2015-02-21 13:54:00|80.709059419360486|3|7203663996|174|35.18634243773306|0|31|342|-80.739|57|35.141204|FRESH MILK|0.52|3|HARRIS TEETER WHOLE MILK|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00072036639967|MILK|DAIRY|-80.70901|80.709017483322825|171|1
35.17335|1dc5938838ede72085356fb32ecdc01e2361ac8b|15.8|2014-12-13 11:17:00|1.4094857484078087|3|7203663995|174|0.6138907664563474|0|26|342|-80.70901|57|35.17335|FRESH MILK|1.96|3|HARRIS TEETER 2% MILK|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|0.61471665291522548|00072036639981|MILK|DAIRY|-80.70901|1.4086379605250285|174|4
35.17335|89b8d87c1f6b704ce2544f8a0dbc00370c5afc5c|6.98|2015-02-07 14:52:00|1.4094857484078087|3|7203663995|174|0.6138907664563474|0|26|342|-80.70901|57|35.17335|FRESH MILK|0.72|3|HARRIS TEETER 2% MILK|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|0.61471665291522548|00072036639981|MILK|DAIRY|-80.70901|1.4086379605250285|174|2
35.17335|aafe01b096777b9c693853e3142e66335cee51eb|7.98|2014-09-27 12:20:00|1.4094857484078087|3|7203663995|174|0.6138907664563474|0|26|342|-80.70901|57|35.17335|FRESH MILK|1.02|3|HARRIS TEETER 2% MILK|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|0.61471665291522548|00072036639981|MILK|DAIRY|-80.70901|1.4086379605250285|174|2
35.17335|5a44497ff2f69be87c9377fd0db5d97af292cb7b|7.98|2014-10-11 16:14:00|1.4094857484078087|3|7203663995|174|0.6138907664563474|0|26|342|-80.70901|57|35.17335|FRESH MILK|1.02|3|HARRIS TEETER 2% MILK|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|0.61471665291522548|00072036639981|MILK|DAIRY|-80.70901|1.4086379605250285|174|2
35.17335|30ed6b00997474e8723dfe473f26af20f6f1a3f7|3.75|2015-01-06 16:14:00|80.709059419360486|3|4610000094|174|35.186342439156661|0|31|333|-80.62331|52|35.140781|PARMESAN CHEESE|1.25|3|SARGENTO ARTISAN PARMESAN|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|35.187384292804154|00046100000595|CHEESE|DAIRY|-80.70901|80.709010791965582|39|1
35.17335|e3b7c7bfeae60ab4b31ef09ff761900fe029596c|7.1|2014-11-29 15:49:00|1.4094857484078087|3|7433610102|174|0.6138907664563474|0|26|342|-80.70901|57|35.17335|FRESH MILK|2.16|3|HIGHLAND CREST 2% REDUCE FAT|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|0.61471665291522548|00074336101021|MILK|DAIRY|-80.70901|1.4086379605250285|174|2
35.17335|20e707a1523cec4833004db795536f295e8f620c|2.99|2015-02-23 15:28:00|1.4094857484078087|3|7433610102|174|0.6138907664563474|0|26|342|-80.70901|57|35.17335|FRESH MILK|0.0|3|HIGHLAND CREST 2% REDUCE FAT|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|0.61471665291522548|00074336101021|MILK|DAIRY|-80.70901|1.4086379605250285|174|1
35.17335|c419d3031bd315c019f9a889ab6093f5cd1c7489|6.98|2015-01-17 16:29:00|1.4094857484078087|3|7203663995|174|0.6138907664563474|0|26|342|-80.70901|57|35.17335|FRESH MILK|0.92|3|HARRIS TEETER 2% MILK|5a84427792e2a46a6d6c79cd82e3a93ad3389cf5|0.897746171222875|0.61471665291522548|00072036639981|MILK|DAIRY|-80.70901|1.4086379605250285|174|2
35.175855|35b217d0c251fa0ae91e2cb21e9e10d9de1e593e|8.49|2015-02-28 14:58:00|80.850140887259911|2|3100065020|218|35.184131225048482|0|50|1280|-80.848528|48|35.053394|MULTI SERVE MEALS|0.0|5|BER CKN ALF VEGGIE PENNE|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00031000650094|FROZEN MEALS|FROZEN|-80.85013|80.850142830593981|11|1
35.175855|51668969ab45f5746368eebca2a452323c5a2500|3.49|2015-01-18 13:23:00|80.850140887259911|2|4588822215|218|35.184131225048482|0|50|6730|-80.848528|1564|35.053394|RETRACTABLE BALL POINT PEN|0.0|18|Z-GRIP RETRACT BALLPOINT PEN|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00045888222151|SCHOOL & OFFICE SUPPLY|GM|-80.85013|80.850142830593981|11|1
35.175855|57c7cc4c073f319339cef32aa3fafb25ed2aff53|4.58|2015-01-31 16:29:00|80.850140887259911|2|20165700000|218|35.184131225048482|0|50|297|-80.848528|49|35.053394|GROUND BEEF|1.02|2|HT GROUND BEEF CHUCK 80% LEAN|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00201657000003|BEEF|MEAT|-80.85013|80.850142830593981|11|1
35.175855|95b49d21d7d388fe739f2b630f7c17caa6a1ecd7|8.29|2015-01-08 15:23:00|80.850140887259911|2|20165700000|218|35.184131225048482|0|50|297|-80.848528|49|35.053394|GROUND BEEF|0.9099999999999999|2|HT GROUND BEEF CHUCK 80% LEAN|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00201657000003|BEEF|MEAT|-80.85013|80.850142830593981|11|2
35.175855|087af954efab07b0f3921ca3ca77a7020a8db804|11.81|2014-12-28 15:48:00|80.850140887259911|2|20165700000|218|35.184131225048482|0|50|297|-80.848528|49|35.053394|GROUND BEEF|1.38|2|HT GROUND BEEF CHUCK 80% LEAN|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00201657000003|BEEF|MEAT|-80.85013|80.850142830593981|11|2
35.175855|9eba03b7313cd47577e0ef32efdcfa5ea14e2bf5|4.53|2014-12-20 15:32:00|80.850140887259911|2|20165700000|218|35.184131227095108|0|50|297|-80.816172|49|35.059823|GROUND BEEF|0.5|2|HT GROUND BEEF CHUCK 80% LEAN|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00201657000003|BEEF|MEAT|-80.85013|80.850140673078798|66|1
35.175855|78d842ba1cc265d10f436c2b52ec3ed482d6e2b0|4.35|2015-02-21 15:15:00|80.850140887259911|2|20323600000|218|35.184131225048482|0|50|641|-80.848528|137|35.053394|PREMIUM PORK|0.0|2|PORK LOIN END CHOPS BONE-IN|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00203236000008|PORK|MEAT|-80.85013|80.850142830593981|11|1
35.175855|04def45f0d8ff86afadc786de4d70d2b5a39bd55|4.49|2014-11-15 15:00:00|80.850140887259911|2|7203695649|218|35.184131225048482|0|50|1699|-80.848528|387|35.053394|EVERYDAY (COOKIES)|0.0|14|HT CHOCO, CHOCO FROSTED COOKIE|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00072036956514|COOKIES|BAKERY|-80.85013|80.850142830593981|11|1
35.175855|be42e53419144deaa7a9667f3d10159f1387b2d7|7.99|2014-09-28 15:10:00|80.850140887259911|2|38151901250|218|35.184131225048482|0|50|3628|-80.848528|1055|35.053394|WOMEN-ROOT TOUCH UP|2.0|17|NICE/EZ ROOT 4R DRK AUBURN|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00381519012525|HAIR COLORING/PERM|HBC|-80.85013|80.850142830593981|11|1
35.175855|d27b738002d3a039eadbd878bd4ba3a2a643efd4|7.3|2014-11-29 15:34:00|80.850140887259911|2|4610000094|218|35.184131227095108|0|50|318|-80.816172|52|35.059823|SHREDDED/GRATED CHEESE|0.0|3|SARGENTO CB 6 CHEESE ITALIAN|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00046100000915|CHEESE|DAIRY|-80.85013|80.850140673078798|66|2
35.175855|5c6c37f00a35acfd2e8d421f1b3e31b1acb3bc60|0.85|2014-10-05 14:23:00|80.850140887259911|2|7203663222|218|35.184131225048482|0|50|330|-80.848528|55|35.053394|EGGS|0.0|3|HT GRADE A    LARGE EGGS 6 CT.|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00072036632227|EGGS FRESH|DAIRY|-80.85013|80.850142830593981|11|1
35.175855|3fabd323919d75fe0bf75b0ac3c1d231531f80fa|12.19|2014-10-18 15:52:00|80.850140887259911|2|1380023260|218|35.184131227095108|0|50|1280|-80.816172|48|35.059823|MULTI SERVE MEALS|0.0|5|STOUFF CKN ALFREDO LRG FAMILY|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00013800232700|FROZEN MEALS|FROZEN|-80.85013|80.850140673078798|66|1
35.175855|965c93f59571fafbe278e2e99c54d72879b5e342|14.07|2014-09-20 15:12:00|80.850140887259911|2|4900002468|218|35.184131227095108|0|50|54|-80.816172|8|35.059823|DIET|3.57|23|DIET COKE .5 LITER/6 PK.|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.85013|80.850140673078798|66|3
35.175855|3c726470cc6f3a18edb6ecd5014e438c3c57df3b|9.38|2014-10-12 14:59:00|80.850140887259911|2|4900002468|218|35.184131225048482|0|50|54|-80.848528|8|35.053394|DIET|2.38|23|DIET COKE .5 LITER/6 PK.|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.85013|80.850142830593981|11|2
35.175855|b87f9216ff1e66da7a34c8630f11e03942e4eae0|9.98|2015-02-08 15:49:00|80.850140887259911|2|4900002468|218|35.184131225048482|0|50|54|-80.848528|8|35.053394|DIET|0.0|23|DIET COKE .5 LITER/6 PK.|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.85013|80.850142830593981|11|2
35.175855|a678b290753cc3f3ab3f2f6073ca86bd2bc71691|9.38|2014-11-22 15:31:00|80.850140887259911|2|4900002468|218|35.184131225048482|0|50|54|-80.848528|8|35.053394|DIET|0.0|23|DIET COKE .5 LITER/6 PK.|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.85013|80.850142830593981|11|2
35.175855|3bf087bd48b02084a26f1b540bdc5c798b7c215e|9.98|2015-03-09 17:46:00|80.850140887259911|2|4900002468|218|35.184131225048482|0|50|54|-80.848528|8|35.053394|DIET|4.98|23|DIET COKE .5 LITER/6 PK.|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.85013|80.850142830593981|11|2
35.175855|c3a8929f7478d1b0536af707fb7c3b7f132fd063|14.97|2015-01-25 16:21:00|80.850140887259911|2|4900002468|218|35.184131225048482|0|50|54|-80.848528|8|35.053394|DIET|2.31|23|DIET COKE .5 LITER/6 PK.|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.85013|80.850142830593981|11|3
35.175855|b66ff85865e1d2a2535d4f6e8f060c6165ed4b2a|14.07|2014-10-26 14:40:00|80.850140887259911|2|4900002468|218|35.184131225048482|0|50|54|-80.848528|8|35.053394|DIET|2.35|23|DIET COKE .5 LITER/6 PK.|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.85013|80.850142830593981|11|3
35.175855|90532e48a9623597f87bea278718b24a37cecdcc|9.98|2015-02-14 15:25:00|80.850140887259911|2|4900002468|218|35.184131225048482|0|50|54|-80.848528|8|35.053394|DIET|2.0|23|DIET COKE .5 LITER/6 PK.|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.85013|80.850142830593981|11|2
35.175855|4c22148f0cf762d7d6234d86abe5f64272fc73d4|14.07|2014-12-14 15:56:00|80.850140887259911|2|4900002468|218|35.184131225048482|0|50|54|-80.848528|8|35.053394|DIET|0.0|23|DIET COKE .5 LITER/6 PK.|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.85013|80.850142830593981|11|3
35.175855|74550c02384d0838d05077de7a7f80371c84436b|14.07|2014-11-05 15:03:00|80.850140887259911|2|4900002468|218|35.184131227095108|0|50|54|-80.816172|8|35.059823|DIET|2.34|23|DIET COKE .5 LITER/6 PK.|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.85013|80.850140673078798|66|3
35.175855|730a7a2c2aedef4e24ca109b57bad072595e1ea2|14.07|2014-12-07 15:20:00|80.850140887259911|2|4900002468|218|35.184131225048482|0|50|54|-80.848528|8|35.053394|DIET|2.35|23|DIET COKE .5 LITER/6 PK.|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.85013|80.850142830593981|11|3
35.175855|714456d25b25027ebee248baf05829855cf27e7a|9.38|2014-09-11 17:26:00|80.850140887259911|2|4900002468|218|35.184131225048482|0|50|54|-80.848528|8|35.053394|DIET|2.34|23|DIET COKE .5 LITER/6 PK.|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.85013|80.850142830593981|11|2
35.175855|b0c98ec5809226baabe82381690bb581a7a63e54|8.99|2014-12-04 17:08:00|80.850140887259911|2|7289010011|218|35.184131225048482|0|50|459|-80.848528|83|35.053394|IMPORT BEER|0.0|16|AMSTEL LIGHT 6PK 12OZ BTL|5bd01cd61c23873f76504700fc2106b37bdace07|0.5718676235812749|35.186025810841215|00072890100115|IMPORT BEER|BEER|-80.85013|80.850142830593981|11|1
35.037115|fef10999f524e64da4076b77ac76edfee9634f10|1.55|2014-10-25 15:08:00|1.4091206135396188|2|78616201000|27|0.611513017149893|0|47|31|-80.8062|4|35.037115|NON CARBONATED WATER|0.55|1|VIT WATER ZERO RISE|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00786162002983|BOTTLED WATER|G1 GROCERY|-80.8062|1.4103342460250419|27|1
35.037115|92ca833089d94d35099a3257f0ac7252bfdf520b|1.59|2014-09-20 13:15:00|1.4091206135396188|2|78616201000|27|0.611513017149893|0|47|31|-80.8062|4|35.037115|NON CARBONATED WATER|0.59|1|VIT WATER ZERO RISE|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00786162002983|BOTTLED WATER|G1 GROCERY|-80.8062|1.4103342460250419|27|1
35.037115|b534c2d4cf4b3c9a8aa2b7c9843da04652267a20|0.75|2014-12-14 12:04:00|80.811922674510953|2||27|35.038660345157815|0|12|1617|-80.848528|373|35.053394|ROLLS BULK|0.0|14|BULK ROLLS|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00072036955555|ROLLS|BAKERY|-80.8062|80.806200040759364|11|1
35.037115|e24775010e468a5c2bb7061944a43257fb7d9e89|1.97|2015-02-28 15:23:00|1.4091206135396188|2|7203697723|27|0.611513017149893|0|47|223|-80.8062|35|35.037115|SUGAR SUBSTITUTES|0.2|1|HT SWEETENER - SUCRALOSE|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00072036977236|SUGAR/SUBSTITUTES|G1 GROCERY|-80.8062|1.4103342460250419|27|1
35.037115|948a1a6c47ff0c40290216f0790afb0e64ba5488|3.98|2015-02-14 17:18:00|1.4091206135396188|2|7294075600|27|0.611513017149893|0|47|257|-80.8062|39|35.037115|TOMATOES|0.98|1|TUTTOROSSO TOMATO WHL PLUM|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00072940754008|VEGETABLES-CAN/JAR|G1 GROCERY|-80.8062|1.4103342460250419|27|2
35.037115|79fcc3b5942df035d7c18d2db9acece1a321e0ab|1.77|2015-01-31 16:41:00|1.4091206135396188|2|7203657031|27|0.611513017149893|0|47|322|-80.8062|53|35.037115|SOUR CREAM|0.18|3|HT LIGHT SOUR CREAM|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00072036590343|CULTURES|DAIRY|-80.8062|1.4103342460250419|27|1
35.037115|229daf732add01264b6e326a3bde29ce79454c77|5.69|2015-01-25 15:13:00|1.4091206135396188|2|7203663043|27|0.611513017149893|0|47|974|-80.8062|201|35.037115|FRESH TURKEY|2.85|2|HT 85% LEAN GROUND TURKEY|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00072036630438|POULTRY|MEAT|-80.8062|1.4103342460250419|27|1
35.037115|db7556e198606f9e08af5e610e4a2117dbe27b3c|0.79|2015-01-17 14:26:00|1.4091206135396188|2|7203688001|27|0.611513017149893|0|47|527|-80.8062|64|35.037115|FRESH CARROTS|0.0|4|HT WHOLE CARROTS 1LB BAG|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00072036880017|FRESH PRODUCE|PRODUCE|-80.8062|1.4103342460250419|27|1
35.037115|f6bd11c0b1eafd930ca517fa248e458187a80b44|0.79|2015-01-09 17:39:00|1.4091206135396188|2|7203688001|27|0.611513017149893|0|47|527|-80.8062|64|35.037115|FRESH CARROTS|0.0|4|HT WHOLE CARROTS 1LB BAG|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00072036880017|FRESH PRODUCE|PRODUCE|-80.8062|1.4103342460250419|27|1
35.037115|0020c8148f64094d2a74c583255732107feb8176|4.58|2014-10-12 12:25:00|1.4091206135396188|2|4118804070|27|0.611513017149893|0|47|257|-80.8062|39|35.037115|TOMATOES|1.14|1|FURMANO TOMATO PETITE 28|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00041188046749|VEGETABLES-CAN/JAR|G1 GROCERY|-80.8062|1.4103342460250419|27|2
35.037115|c583ba0db6d5f7aeebfa9c833e62b4b39d203bd8|3.29|2015-01-30 19:20:00|1.4091206135396188|2|5210007127|27|0.611513017149893|0|47|220|-80.8062|34|35.037115|PEPPER|0.0|1|MC CRUSHED RED PEPPER FAM SIZE|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00052100071275|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.8062|1.4103342460250419|27|1
35.037115|caf04662a102c54fdf27e0180c80a87504d9827e|7.35|2014-11-16 11:51:00|1.4091206135396188|2|4470002268|27|0.611513017149893|0|47|481|-80.8062|100|35.037115|CENTER CUT BACON|3.68|19|OSCAR MAYER CTR SLICED BACON|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00044700022689|BACON|CASE READY MEATS|-80.8062|1.4103342460250419|27|1
35.037115|1d0e8eba5c991664b5492efa38b9233419ed6530|21.99|2014-10-17 15:41:00|80.811922674510953|2|9870908850|27|35.038660345146859|0|12|9985|-80.699909|890|35.002628|NFS-LUX-CAB SAUVIGNON|0.0|13|CATENA CABERNET SAUVIGNON RSV|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00098709088504|LUXURY (OVER $20)|WINE|-80.8062|80.806200228358577|477|1
35.037115|7291e17a0b37b48703d8795b49f7bfbdcfdee140|1.69|2015-01-09 11:54:00|80.811922674510953|2|4900000044|27|35.03866032912331|0|12|54|-80.662946|8|35.412407|DIET|0.0|23|CB COKE ZERO 20 OZ|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00049000040869|CARBONATED BEVERAGES|BEVERAGE|-80.8062|80.806208597970979|68|1
35.037115|a0562fc8713ced244c06d339cd6eb3fc784b6d1c|1.69|2015-01-22 13:15:00|80.811922674510953|2|4900000044|27|35.038660345157815|0|12|54|-80.848528|8|35.053394|DIET|0.0|23|CB COKE ZERO 20 OZ|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00049000040869|CARBONATED BEVERAGES|BEVERAGE|-80.8062|80.806200040759364|11|1
35.037115|6854bb8264d95ace83078a8bffff294fb0c0dc83|4.99|2014-12-30 16:26:00|1.4091206135396188|2|3700047984|27|0.611513017149893|0|47|726|-80.8062|73|35.037115|NFS-BODY WASHES|2.5|1|GILL DRY SKIN HYDRATOR&BDYWSH|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00037000479840|PERSONAL SOAP/BATH ADDITIVES|G1 GROCERY|-80.8062|1.4103342460250419|27|1
35.037115|7990e2abe9d4eacb3a2f6ac5bc3ebe470077e077|4.99|2014-10-18 15:27:00|1.4091206135396188|2|4242101480|27|0.611513017149893|0|47|482|-80.8062|100|35.037115|PRECOOKED BACON|0.6|19|BOARS HEAD FULLY COOKED BACON|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00042421014808|BACON|CASE READY MEATS|-80.8062|1.4103342460250419|27|1
35.037115|2382bf661c791d6760d780781da74c92cab9aadc|3.74|2015-01-05 13:06:00|80.811922674510953|2|20598400000|27|35.038660343461636|0|12|1822|-80.80146|410|35.17739|BH CHICKEN|0.68|6|BOARS HEAD EVERROAST CKN BRST|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00205984000002|BH MEAT|DELI|-80.8062|80.806202796705563|208|1
35.037115|db2940312d753709f436456a763b8adf45081a41|0.79|2014-11-30 11:38:00|1.4091206135396188|2||27|0.611513017149893|0|47|532|-80.8062|64|35.037115|FRESH CUCUMBERS|0.0|4|COO CUCUMBERS S/S|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00204062000002|FRESH PRODUCE|PRODUCE|-80.8062|1.4103342460250419|27|1
35.037115|ea19ca88092a8ae7a7cafd8954386ea0465c0f73|0.79|2015-02-21 15:13:00|1.4091206135396188|2||27|0.611513017149893|0|47|532|-80.8062|64|35.037115|FRESH CUCUMBERS|0.0|4|COO CUCUMBERS S/S|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00204062000002|FRESH PRODUCE|PRODUCE|-80.8062|1.4103342460250419|27|1
35.037115|397e7f54a1af69baddb8f22978ce71186c668c54|0.79|2015-03-08 12:07:00|1.4091206135396188|2||27|0.611513017149893|0|47|532|-80.8062|64|35.037115|FRESH CUCUMBERS|0.0|4|COO CUCUMBERS S/S|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00204062000002|FRESH PRODUCE|PRODUCE|-80.8062|1.4103342460250419|27|1
35.037115|1675314d34805d10e594e77f7be797cebf58527e|0.79|2014-11-09 13:18:00|1.4091206135396188|2||27|0.611513017149893|0|47|532|-80.8062|64|35.037115|FRESH CUCUMBERS|0.2|4|COO CUCUMBERS S/S|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00204062000002|FRESH PRODUCE|PRODUCE|-80.8062|1.4103342460250419|27|1
35.037115|a43ec23fb720990ff64067bbb62c2c5e98686de7|28.38|2014-12-13 19:27:00|1.4091206135396188|2|20220200000|27|0.611513017149893|0|47|299|-80.8062|49|35.037115|ANGUS BEEF|7.1|2|ANGUS BEEF FILET MIGNON|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00202204000002|BEEF|MEAT|-80.8062|1.4103342460250419|27|2
35.037115|92b1eaf2289d2e901d7e8c078e67280cf3c64ae2|1.67|2014-11-12 17:51:00|1.4091206135396188|2|3663201899|27|0.611513017149893|0|47|343|-80.8062|59|35.037115|PUDDINGS|0.77|3|CREAMERY CHERRY CHEESECAKE|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00036632018939|SNACKS/SPREADS/DIPS-DAIRY|DAIRY|-80.8062|1.4103342460250419|27|1
35.037115|9cb0eaa5efcf6888797287da185886bd785f7d9e|3.42|2015-01-26 09:55:00|80.811922674510953|2|20413100000|27|35.038660345140997|0|12|500|-80.992182|64|35.103409|FRESH APPLES|0.17|4|FUJI APPLES|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00891658001316|FRESH PRODUCE|PRODUCE|-80.8062|80.806200281440724|88|2
35.037115|1c07e231345bd104f14267a2f5076d9f1e5e45d9|6.99|2015-01-11 11:18:00|1.4091206135396188|2|7203663045|27|0.611513017149893|0|47|974|-80.8062|201|35.037115|FRESH TURKEY|0.0|2|HT 99% LEAN GRND TURKEY BREAST|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00072036630452|POULTRY|MEAT|-80.8062|1.4103342460250419|27|1
35.037115|50ce5208f5fc0921b2df24b078eb9e5b2bb76b69|3.58|2014-10-26 10:22:00|1.4091206135396188|2|4850001775|27|0.611513017149893|0|47|335|-80.8062|56|35.037115|ORANGE JUICE-REGRIGERATED|1.58|3|TROPICANA PP ORIGINAL 12 OZ|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00048500017753|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.8062|1.4103342460250419|27|2
35.037115|794c2e5445856dd4abb3e0a2fae078e5d8d404b3|1.29|2015-02-06 17:21:00|1.4091206135396188|2||27|0.611513017149893|0|47|508|-80.8062|64|35.037115|FRESH GRAPEFRUIT|0.29|4|RED GRAPEFRUIT LRG|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00204027000009|FRESH PRODUCE|PRODUCE|-80.8062|1.4103342460250419|27|1
35.037115|f150f2cd182b9ece6f9c285c76308fb817f9973b|0.44|2015-01-07 17:51:00|1.4091206135396188|2||27|0.611513017149893|0|47|502|-80.8062|64|35.037115|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00204011000008|FRESH PRODUCE|PRODUCE|-80.8062|1.4103342460250419|27|1
35.037115|13a33f26d60f8f1f1f74db9ddca3a91cd1d113b5|0.55|2014-12-07 11:51:00|80.811922674510953|2||27|35.038660345157815|0|12|502|-80.848528|64|35.053394|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00204011000008|FRESH PRODUCE|PRODUCE|-80.8062|80.806200040759364|11|1
35.037115|148d8728a7310f2ecdadac6f6554de5e2e777549|2.97|2015-01-06 19:10:00|80.811922674510953|2|20597100000|27|35.03866034184891|0|12|1821|-80.661096|410|35.172688|BH TURKEY|0.54|6|BOARS HEAD LOW SODIUM TURKEY|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00205971000008|BH MEAT|DELI|-80.8062|80.806203905984418|474|1
35.037115|8c545d1e7b0b11b650921aa492fd1b4510cad233|3.65|2014-10-01 10:09:00|80.811922674510953|2|95546|27|35.038660343743494|0|12|1582|-80.709466|369|35.124987|NFS BEVERAGE TEA|0.0|22|CHAI TEA LATTE GRANDE|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00000000955460|NFS STARBUCKS|COFFEE SHOP|-80.8062|80.806202553845253|157|1
35.037115|26880d139045b304353dd12875dfac53232c6494|1.5|2015-02-08 14:47:00|1.4091206135396188|2|20892500000|27|0.611513017149893|0|47|645|-80.8062|201|35.037115|FRESH POULTRY SAUSAGE|0.0|2|CHICKEN ITALIAN HOT SAUSAGE|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00208915000003|POULTRY|MEAT|-80.8062|1.4103342460250419|27|1
35.037115|8056ac2a8878b68dc82174fbb03b090d4203eb55|12.95|2014-12-14 12:07:00|80.811922674510953|2|76211191510|27|35.038660345157815|0|12|1583|-80.848528|370|35.053394|VIA|3.89|22|KCUP CHRISTMAS 12 CT|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00762111915108|STARBUCKS|COFFEE SHOP|-80.8062|80.806200040759364|11|1
35.037115|fe4d1b5ecbb65ce2a2cc39bd7090dac30e92180c|0.8|2014-12-12 08:06:00|80.811922674510953|2|97049|27|35.038660345157815|0|12|1589|-80.848528|369|35.053394|NFS BEVERAGE ESPRESSO|0.16|22|ADD ESPRESSO SHOTS|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00000000970490|NFS STARBUCKS|COFFEE SHOP|-80.8062|80.806200040759364|11|1
35.037115|58b277495228ea454b1f162d234440cd59ffb48d|4.2|2014-11-10 08:32:00|80.811922674510953|2|96825|27|35.038660342422133|0|12|1581|-80.810056|369|35.219587|NFS BEVERAGE BREWED|0.0|22|BREWED COFFEE GRANDE|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00000000968250|NFS STARBUCKS|COFFEE SHOP|-80.8062|80.806203551618239|401|2
35.037115|2849e8c54abe56a70997f551d84dd1a66ba29ab8|2.1|2015-01-09 08:46:00|80.811922674510953|2|96825|27|35.038660344073158|0|12|1581|-80.837892|369|34.937113|NFS BEVERAGE BREWED|0.0|22|BREWED COFFEE GRANDE|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00000000968250|NFS STARBUCKS|COFFEE SHOP|-80.8062|80.806202236570869|372|1
35.037115|8c69d0a906c07e725faac8a1cf14871d43dac9e6|1.79|2014-09-15 08:53:00|80.811922674510953|2|2500000024|27|35.038660344192806|0|12|335|-80.825175|56|35.152722|ORANGE JUICE-REGRIGERATED|0.79|3|SIMPLY ORANGE JUICE CALCIUM|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00025000000355|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.8062|80.806202109660063|160|1
35.037115|fb75784772c4d1d0b4a57cf40c6645280ee304e5|1.79|2014-09-17 08:47:00|80.811922674510953|2|2500000024|27|35.038660344192806|0|12|335|-80.825175|56|35.152722|ORANGE JUICE-REGRIGERATED|0.0|3|SIMPLY ORANGE JUICE CALCIUM|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00025000000355|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.8062|80.806202109660063|160|1
35.037115|a3a970865a3756a64b51fabdcad096337d448d6e|20.97|2014-10-09 18:02:00|80.811922674510953|2|3798298222|27|35.038660345157815|0|12|2017|-80.848528|505|35.053394|STRETCHED CURD CHEESE|14.04|6|PALAZZINA MOZZARELLA BALLS|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00037982982222|SPECIALTY CHEESE|DELI|-80.8062|80.806200040759364|11|3
35.037115|06eefa9dcf5a543751ebc26c6228b6f73f77961f|1.59|2015-02-10 13:36:00|80.811922674510953|2|1200000129|27|35.038660345157815|0|12|54|-80.848528|8|35.053394|DIET|0.25|23|DIET SUNKIST ORANGE 20 OZ|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00078000122404|CARBONATED BEVERAGES|BEVERAGE|-80.8062|80.806200040759364|11|1
35.037115|8b5ba781fd1d73d1f810e8e3231cdd4340c51c69|1.55|2014-12-22 08:43:00|80.811922674510953|2|78616201000|27|35.038660332886963|0|12|31|-80.861571|4|35.444615|NON CARBONATED WATER|0.55|1|VIT WATER ZERO POWER- C|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00786162003737|BOTTLED WATER|G1 GROCERY|-80.8062|80.806207521550036|340|1
35.037115|5b546c68cbd3872d38d6f21fe434fb28e36f0dc6|1.55|2014-11-14 12:06:00|80.811922674510953|2|78616201000|27|35.038660344704311|0|12|31|-80.97058|4|35.03469|NON CARBONATED WATER|0.55|1|VIT WATER ZERO POWER- C|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00786162003737|BOTTLED WATER|G1 GROCERY|-80.8062|80.806201446532981|82|1
35.037115|0552502bfbf3a055e22bceca9bef6c5ff4f544ef|3.19|2014-10-04 08:34:00|1.4091206135396188|2|61126971646|27|0.611513017149893|0|47|97|-80.8062|8|35.037115|ENERGY DRINKS|0.0|23|CB RED BULL SF 12 OZ CAN|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|0.61242566243833529|00611269716467|CARBONATED BEVERAGES|BEVERAGE|-80.8062|1.4103342460250419|27|1
35.037115|41f21014bafbb52d4fee0e3ed3121a9931ee767b|1.0|2014-10-16 12:30:00|80.811922674510953|2|61300873089|27|35.038660331623902|0|12|99|-80.893784|32|35.478031|LIQUID TEA|0.0|1|PP ARIZONA ARNOLD PALMER|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00613008730895|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.8062|80.806207899162558|179|1
35.037115|91d8a196d28b49728334deedff6f93ce5cfdbae5|2.35|2015-02-20 07:58:00|80.811922674510953|2|96826|27|35.038660338129866|0|12|1581|-80.737839|369|35.297134|NFS BEVERAGE BREWED|0.0|22|BREWED COFFEE VENTI|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00000000968260|NFS STARBUCKS|COFFEE SHOP|-80.8062|80.806205692321541|258|1
35.037115|c39848eddd6c41da8e8ab4ebbeb0a99d77043c5d|1.55|2014-12-11 13:54:00|80.811922674510953|2|78616201000|27|35.038660344192806|0|12|31|-80.825175|4|35.152722|NON CARBONATED WATER|0.55|1|VIT WATER ZERO REVIVE|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00786162003744|BOTTLED WATER|G1 GROCERY|-80.8062|80.806202109660063|160|1
35.037115|eb2f3cfdb8b135d030393ac8a8e692db8d6f81ae|1.59|2014-10-06 13:15:00|80.811922674510953|2|78616201000|27|35.038660335030933|0|12|31|-80.86175|4|35.40953|NON CARBONATED WATER|0.59|1|VIT WATER ZERO REVIVE|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00786162003744|BOTTLED WATER|G1 GROCERY|-80.8062|80.806206832970517|209|1
35.037115|8233f482dbf288f3be3557075ca81b71ab312bf8|6.99|2014-09-13 12:39:00|80.811922674510953|2|7172807100|27|35.038660345129848|0|12|848|-80.816172|104|35.059823|NAT/ORG DINNER SAUSAGE|0.0|19|BILINSKI ORG SPINACH SAUSAGE|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00071728071009|DINNER SAUSAGE|CASE READY MEATS|-80.8062|80.806200361375488|66|1
35.037115|f6b1ed45f447e061973cb566ebbc5de76c4e9c51|1.57|2015-01-20 17:19:00|80.811922674510953|2||27|35.038660342520188|0|12|500|-80.8438|64|35.23102|FRESH APPLES|0.16|4|GALA APPLES|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00204135000007|FRESH PRODUCE|PRODUCE|-80.8062|80.806203487388444|205|1
35.037115|c6100a5da4f198069146e6cac1713f3d3da00498|1.55|2014-11-13 15:44:00|80.811922674510953|2|78616201000|27|35.038660335195132|0|12|31|-80.782849|4|35.372142|NON CARBONATED WATER|0.55|1|VIT WATER ZERO XXX|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00786162002969|BOTTLED WATER|G1 GROCERY|-80.8062|80.806206777350098|122|1
35.037115|c98b81eee1562e9b6ef903dd178ab160e1787d18|1.69|2015-02-09 13:38:00|80.811922674510953|2|4900000044|27|35.038660342520188|0|12|54|-80.8438|8|35.23102|DIET|0.0|23|CB DIET DR PEPPER 20OZ NR|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00078000083408|CARBONATED BEVERAGES|BEVERAGE|-80.8062|80.806203487388444|205|1
35.037115|b288f4fc2394c8963a2e32207e6ec65b6d2dee86|3.65|2014-12-03 07:02:00|80.811922674510953|2|96844|27|35.038660343743494|0|12|1589|-80.709466|369|35.124987|NFS BEVERAGE ESPRESSO|0.0|22|CAFFE LATTE GRANDE|5c1bb2ba133cb9fcd458b9a9abcf929a13257725|0.10677961855545227|35.037868710371079|00000000968440|NFS STARBUCKS|COFFEE SHOP|-80.8062|80.806202553845253|157|1
35.585842|9c4c7a6074982b6e6a0cef5243ce3f9952499a60|2.99|2015-03-06 17:12:00|1.4102725052409182|2|7044650000|99|0.6210901099944839|0|1|498|-80.875654|111|35.585842|PICKLES & SAUERKRAUT|0.9|19|BOARS HEAD SAUERKRAUT 32 OZ|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|0.61833652052202714|00070446500006|MISC. PACKAGED MEATS|CASE READY MEATS|-80.875654|1.411546447003722|99|1
35.585842|ee27b1af7670384ce7d05314d3d933ae8ac1e0ac|7.58|2014-12-28 17:43:00|80.849735164501183|2|7127930104|99|35.606598881305828|0|11|555|-80.992182|64|35.103409|PACKAGED SALADS|0.0|4|F.E. CAESAR SUPREME COMPLETE|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|35.604954314503821|00071279301044|FRESH PRODUCE|PRODUCE|-80.875654|80.875795288845453|88|2
35.585842|fecc1c8cf94c1efbccf6c6db5658de839a63f388|7.58|2014-09-29 19:13:00|80.849735164501183|2|7127930104|99|35.606598881305828|0|11|555|-80.992182|64|35.103409|PACKAGED SALADS|0.0|4|F.E. CAESAR SUPREME COMPLETE|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|35.604954314503821|00071279301044|FRESH PRODUCE|PRODUCE|-80.875654|80.875795288845453|88|2
35.585842|4a9a63ffc650195b6d76f5d1d9d211b417c7acbc|1.67|2014-11-29 21:01:00|80.849735164501183|2|7172053046|99|35.606599069352981|0|11|53|-80.8438|7|35.23102|THEATER BOX|0.0|1|JUNIOR MINTS THEATRE BOX|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|35.604954314503821|00071720530467|CANDY|G1 GROCERY|-80.875654|80.87574430929304|205|1
35.585842|38e963adc49d391106234eb349efee2e4e15c547|4.29|2015-02-25 16:05:00|1.4102725052409182|2|4178000011|99|0.6210901099944839|0|1|201|-80.875654|31|35.585842|POTATO CHIPS|1.3|1|UTZ CRAB CHIPS|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|0.61833652052202714|00041780001580|SNACKS|G1 GROCERY|-80.875654|1.411546447003722|99|1
35.585842|837b3cc2e2d9927acbb1126f9ef6f2f07bb44a24|3.69|2014-12-01 15:59:00|1.4102725052409182|2|4400001570|99|0.6210901099944839|0|1|1256|-80.875654|13|35.585842|WHOLESOME CRACKERS|0.69|1|RITZ TOASTED CHIPS CHEDDAR|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|0.61833652052202714|00044000015701|CRACKERS|G1 GROCERY|-80.875654|1.411546447003722|99|1
35.585842|6fab9ab02aa2d870eb0ff8312f22a44e20429336|8.99|2014-11-21 17:39:00|1.4102725052409182|2|7203688106|99|0.6210901099944839|0|1|583|-80.875654|136|35.585842|NUTS|0.0|4|HT WHOLE NATURAL ALMOND TRAY|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|0.61833652052202714|00072036881069|OTHER MERCHANDISE|PRODUCE|-80.875654|1.411546447003722|99|1
35.585842|fb8dac6c5b66cea5cf9cd3bc2eef761f9fe554a2|6.99|2015-03-05 14:56:00|80.849735164501183|2|4900002890|99|35.606599103399475|0|11|54|-80.945176|8|35.323246|DIET|3.5|23|CHERRY COKE ZERO 12OZ FPK CAN|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|35.604954314503821|00049000047516|CARBONATED BEVERAGES|BEVERAGE|-80.875654|80.875731576455948|166|1
35.585842|4c172ba7692b4d242d07681e19fe44d3a2ee978b|1.79|2014-12-23 15:51:00|1.4102725052409182|2|5210003850|99|0.6210901099944839|0|1|80|-80.875654|34|35.585842|SEASONING PACKETS|0.0|1|MC BEEF STROGANOFF|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|0.61833652052202714|00052100038506|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.875654|1.411546447003722|99|1
35.585842|a4cfa690504cc3dde824b2c2db4f6aa278f33a98|4.31|2014-12-18 15:47:00|1.4102725052409182|2||99|0.6210901099944839|0|1|529|-80.875654|64|35.585842|FRESH ASPARAGUS|0.48|4|GREEN  ASPARAGUS|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|0.61833652052202714|00204080000008|FRESH PRODUCE|PRODUCE|-80.875654|1.411546447003722|99|1
35.585842|72258a31655ae5a8998eebfb4823cc283846c4f1|3.95|2015-01-04 17:07:00|80.849735164501183|2|1410007467|99|35.606598881305828|0|11|1026|-80.992182|162|35.103409|WHEAT|0.0|7|PEP FH HNY WHEAT WP BRD  PP|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|35.604954314503821|00014100098959|SLICED BREAD|COMMERCIAL BAKERY|-80.875654|80.875795288845453|88|1
35.585842|3e509bc63f9265be39ccd21efa85a983d04c5852|2.32|2014-12-28 17:44:00|80.849735164501183|2||99|35.606598881305828|0|11|500|-80.992182|64|35.103409|FRESH APPLES|0.0|4|RED DEL APPLE, WA  48|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|35.604954314503821|00233284000002|FRESH PRODUCE|PRODUCE|-80.875654|80.875795288845453|88|1
35.585842|231012d56504c41db705844acfd22f9d1221a6ba|2.0|2014-12-05 15:42:00|1.4102725052409182|2|812|99|0.6210901099944839|0|1|1639|-80.875654|377|35.585842|BULK (DONUTS)|0.0|14|NEW BULK DONUT CODE|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|0.61833652052202714|00000000008120|DONUTS|BAKERY|-80.875654|1.411546447003722|99|2
35.585842|9f5bd34459e7166df9cdf50ec6e770d102f37839|3.99|2014-11-04 15:08:00|1.4102725052409182|2|7203697785|99|0.6210901099944839|0|1|2022|-80.875654|505|35.585842|BLUE VEINED CHEESE|0.0|6|HT BLUE CHEESE CRMBLD|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|0.61833652052202714|00072036977854|SPECIALTY CHEESE|DELI|-80.875654|1.411546447003722|99|1
35.585842|b287524662e2136f28295dcd60da77c15e6c63e5|2.99|2014-12-30 12:28:00|1.4102725052409182|2|3338365583|99|0.6210901099944839|0|1|522|-80.875654|64|35.585842|FRESH TOMATOES|0.2|4|SWEET GRAPE TOMATO (PINT)|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|0.61833652052202714|00814369011214|FRESH PRODUCE|PRODUCE|-80.875654|1.411546447003722|99|1
35.585842|ec4e58f2c8f7192a42fcb4fb01dd19d509d8d10f|2.99|2015-02-03 13:20:00|1.4102725052409182|2|3338365583|99|0.6210901099944839|0|1|522|-80.875654|64|35.585842|FRESH TOMATOES|0.49|4|SWEET GRAPE TOMATO (PINT)|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|0.61833652052202714|00814369011214|FRESH PRODUCE|PRODUCE|-80.875654|1.411546447003722|99|1
35.585842|69de6e7ea8bbc1366d43d0bd2bfb79b379942ecc|2.29|2014-10-23 14:40:00|1.4102725052409182|2|88937912601|99|0.6210901099944839|0|1|80|-80.875654|34|35.585842|SEASONING PACKETS|0.0|1|RED FORK SC LEM HERB ASPARAGUS|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|0.61833652052202714|00889379126012|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.875654|1.411546447003722|99|1
35.585842|ddd97e9019fae2c8c2a5d9bd6cea3916742207a1|2.19|2015-01-04 15:10:00|1.4102725052409182|2|7478063991|99|0.6210901099944839|0|1|30|-80.875654|4|35.585842|CARBONATED WATER|0.0|1|PERRIER 1LT PET CITRON|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|0.61833652052202714|00074780643184|BOTTLED WATER|G1 GROCERY|-80.875654|1.411546447003722|99|1
35.585842|5573679b0bd1e0b5e9d8bf5880c5d7a0de2cfc64|2.19|2014-10-27 15:35:00|1.4102725052409182|2|7478063991|99|0.6210901099944839|0|1|30|-80.875654|4|35.585842|CARBONATED WATER|0.4|1|PERRIER 1LT PET CITRON|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|0.61833652052202714|00074780643184|BOTTLED WATER|G1 GROCERY|-80.875654|1.411546447003722|99|1
35.585842|f0f912841170cad36b200580435aed3e1e4f3da1|4.98|2015-01-23 09:34:00|1.4102725052409182|2|7478063991|99|0.6210901099944839|0|1|30|-80.875654|4|35.585842|CARBONATED WATER|0.98|1|PERRIER 1LT PET CITRON|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|0.61833652052202714|00074780643184|BOTTLED WATER|G1 GROCERY|-80.875654|1.411546447003722|99|2
35.585842|31855e20b37d0c3a05931e729e581850a839750e|2.19|2014-10-11 18:55:00|1.4102725052409182|2|7478063991|99|0.6210901099944839|0|1|30|-80.875654|4|35.585842|CARBONATED WATER|0.4|1|PERRIER 1 LT PET REG|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|0.61833652052202714|00074780639910|BOTTLED WATER|G1 GROCERY|-80.875654|1.411546447003722|99|1
35.585842|3b2d6062dab1ec3c22f8d91e7576f3a3546a57f5|7.96|2014-10-01 17:07:00|1.4102725052409182|2|7478063991|99|0.6210901099944839|0|1|30|-80.875654|4|35.585842|CARBONATED WATER|0.8|1|PERRIER 1 LT PET REG|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|0.61833652052202714|00074780639910|BOTTLED WATER|G1 GROCERY|-80.875654|1.411546447003722|99|4
35.585842|9dfb1d5402ac5f93a1547fcd624067c5e8bb3be4|5.97|2014-09-12 19:54:00|1.4102725052409182|2|7478063991|99|0.6210901099944839|0|1|30|-80.875654|4|35.585842|CARBONATED WATER|1.47|1|PERRIER 1 LT PET REG|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|0.61833652052202714|00074780639910|BOTTLED WATER|G1 GROCERY|-80.875654|1.411546447003722|99|3
35.585842|03a8385e68a10fbde5df0bd7352b9eea522ba2b9|4.38|2014-11-19 17:34:00|1.4102725052409182|2|7478063991|99|0.6210901099944839|0|1|30|-80.875654|4|35.585842|CARBONATED WATER|0.8|1|PERRIER 1 LT PET REG|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|0.61833652052202714|00074780639910|BOTTLED WATER|G1 GROCERY|-80.875654|1.411546447003722|99|2
35.585842|f67b9f2a6a106b04ddcb9f2dc58431ba35c3c9ca|3.38|2014-10-02 14:00:00|1.4102725052409182|2||99|0.6210901099944839|0|1|503|-80.875654|64|35.585842|FRESH GRAPES|0.23|4|GREEN GRAPES, SEEDLESS 12/16|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|0.61833652052202714|00204022000004|FRESH PRODUCE|PRODUCE|-80.875654|1.411546447003722|99|1
35.585842|18d5cc4f54f94dbb227365db2f478ffede03da02|2.27|2014-10-23 11:48:00|1.4102725052409182|2|2200015586|99|0.6210901099944839|0|1|45|-80.875654|7|35.585842|PEG GUM|0.0|1|ORBIT PEPPERMINT|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|0.61833652052202714|00022000155863|CANDY|G1 GROCERY|-80.875654|1.411546447003722|99|1
35.585842|072f1f0535b1c6c1ecc9eeb10e1927771f158f5c|0.46|2014-10-09 19:55:00|1.4102725052409182|2||99|0.6210901099944839|0|1|502|-80.875654|64|35.585842|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.875654|1.411546447003722|99|1
35.585842|c0b93e3d04c366316a84f88d205ad2d2c7c8cfaa|8.0|2014-11-28 21:28:00|80.849735164501183|2||99|35.606599069352981|0|11|509|-80.8438|64|35.23102|FRESH CITRUS-REMAINING|0.0|4|COO LIMES, LRG|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|35.604954314503821|00204048000002|FRESH PRODUCE|PRODUCE|-80.875654|80.87574430929304|205|16
35.585842|166459d6fe30e8507ffb1b6c32ea2cbfae21e124|6.0|2014-12-29 19:20:00|80.849735164501183|2||99|35.606599069352981|0|11|509|-80.8438|64|35.23102|FRESH CITRUS-REMAINING|0.0|4|COO LIMES, LRG|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|35.604954314503821|00204048000002|FRESH PRODUCE|PRODUCE|-80.875654|80.87574430929304|205|12
35.585842|5346968b6e782a3ebd9ff415136a17870fdb8e43|18.99|2015-02-06 13:23:00|80.849735164501183|2|7119000600|99|35.606598881305828|0|11|156|-80.992182|24|35.103409|NFS-DOG FOOD-DRY|2.0|1|RACH RAY NUTRSH BEEF&RCE 14 LB|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|35.604954314503821|00071190006028|PET FOOD/SUPPLIES|G1 GROCERY|-80.875654|80.875795288845453|88|1
35.585842|ec0e1b2eda45449fbc1cb4c31e73b2919154afd1|16.99|2015-03-08 21:55:00|80.849735164501183|2|7203695339|99|35.606598881305828|0|11|1654|-80.992182|381|35.103409|DESSERT CAKES|0.0|14|"8"" TRIPLE LYR ASST VARIETY CK"|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|35.604954314503821|00072036953391|CAKES|BAKERY|-80.875654|80.875795288845453|88|1
35.585842|d87f4838b82f036fc6940a2ba62bebeb2d631259|4.98|2014-11-01 21:32:00|80.849735164501183|2|60504939530|99|35.606599069352981|0|11|509|-80.8438|64|35.23102|FRESH CITRUS-REMAINING|0.0|4|LEMONS, SMALL 1LB BAG|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|35.604954314503821|00605049395300|FRESH PRODUCE|PRODUCE|-80.875654|80.87574430929304|205|2
35.585842|ce2654ba9c8aa45aca5d5cc255f6a377b1528184|15.58|2014-10-22 06:47:00|1.4102725052409182|2|1291912212|99|0.6210901099944839|0|1|36|-80.875654|10|35.585842|PREMIUM GROUND|2.8|1|SEATTLE'S 4 BEST HENRY'S BLEND|5c55104496090402a36b467ab28346c8d1e3b074|1.4342723412938778|0.61833652052202714|00012919122612|COFFEE|G1 GROCERY|-80.875654|1.411546447003722|99|2
35.059823|255912371b8db0bf3579262a58a776fdca285a7f|1.9|2014-09-16 20:05:00|1.4091206135396188|2||66|0.6119093465164359|0|47|502|-80.816172|64|35.059823|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5d9fb253b347a91c85cbb997da7014c4e3bd9b98|0.6518340734283655|0.61242566243833529|00204011000008|FRESH PRODUCE|PRODUCE|-80.816172|1.4105082902580508|66|1
35.059823|9ea4ef739c01265a3648448af91f7dd8f06fec60|0.93|2014-10-03 11:08:00|80.816179662140996|2||66|35.069256528795776|0|41|565|-80.848528|64|35.053394|REDUCED PRODUCE|0.0|4|PRODUCE REWRAP BY LB|5d9fb253b347a91c85cbb997da7014c4e3bd9b98|0.6518340734283655|35.070508771677183|00204844000008|FRESH PRODUCE|PRODUCE|-80.816172|80.816174455744203|11|1
35.059823|de07ca2eeae9ef7a062855a0b9686af7a5925ce2|1.0|2014-09-21 19:31:00|80.816179662140996|2|3700038592|66|35.069256528795776|0|41|4169|-80.848528|1085|35.053394|TRAIL SIZE TOOTHPASTE|0.0|17|CREST PLUS SCOPE PASTE TRAVEL|5d9fb253b347a91c85cbb997da7014c4e3bd9b98|0.6518340734283655|35.070508771677183|00037000385929|TRIAL SIZE|HBC|-80.816172|80.816174455744203|11|1
35.059823|393c02bbbdd73377a2c443a92a7a9b6f6bb9e56c|1.79|2014-10-06 12:48:00|80.816179662140996|2|7203663158|66|35.069256528795776|0|41|495|-80.848528|108|35.053394|NON REFRIGERATED|0.9|19|HT CORN TORTILLA 30CT|5d9fb253b347a91c85cbb997da7014c4e3bd9b98|0.6518340734283655|35.070508771677183|00072036631589|TORTILLAS|CASE READY MEATS|-80.816172|80.816174455744203|11|1
35.059823|30f6ebd3d0cbd548efcc58f2feb84fde616a60c5|3.99|2014-10-15 12:16:00|80.816179662140996|2|7203663089|66|35.069256528795776|0|41|345|-80.848528|57|35.053394|ORGANIC MILK|0.0|3|HTO ORGANIC CRTN MILK FAT FREE|5d9fb253b347a91c85cbb997da7014c4e3bd9b98|0.6518340734283655|35.070508771677183|00072036630896|MILK|DAIRY|-80.816172|80.816174455744203|11|1
35.059823|5399f520f5acc63fc5af2ba2d38f93f6551a858c|3.99|2014-09-12 20:06:00|1.4091206135396188|2|8500002183|66|0.6119093465164359|0|47|9936|-80.816172|885|35.059823|NFS POP MERLOT|0.0|13|LIBERTY CREEK MERLOT TETRA|5d9fb253b347a91c85cbb997da7014c4e3bd9b98|0.6518340734283655|0.61242566243833529|00085000021835|POPULAR (4-$7.99)|WINE|-80.816172|1.4105082902580508|66|1
35.059823|ad3369fa8bc3d7add33f781aa2f14d314f86ab51|8.99|2014-10-19 15:53:00|1.4091206135396188|2|7199009532|66|0.6119093465164359|0|47|458|-80.816172|82|35.059823|CRAFT BEER|0.0|16|BLUE MOON SEASONAL 6PK|5d9fb253b347a91c85cbb997da7014c4e3bd9b98|0.6518340734283655|0.61242566243833529|00071990095321|DOMESTIC BEER|BEER|-80.816172|1.4105082902580508|66|1
35.059823|007ed1c2ea4e5f07cc7b2b2d12accc08bb442cb1|4.99|2014-09-27 17:30:00|1.4091206135396188|2||66|0.6119093465164359|0|47|558|-80.816172|64|35.059823|SPECIALTY-VEGETABLES|0.0|4|#STALK BRUSSEL SPROUTS|5d9fb253b347a91c85cbb997da7014c4e3bd9b98|0.6518340734283655|0.61242566243833529|00233083000005|FRESH PRODUCE|PRODUCE|-80.816172|1.4105082902580508|66|1
35.059823|ada292656583414ebd10ed336d61cc9cb146e1de|11.99|2014-09-28 18:06:00|80.816179662140996|2|8130800132|66|35.069256528795776|0|41|9983|-80.848528|889|35.053394|NFS-SPARKLING|0.0|13|CUPCAKE PROSECCO|5d9fb253b347a91c85cbb997da7014c4e3bd9b98|0.6518340734283655|35.070508771677183|00081308001326|SPARKLING|WINE|-80.816172|80.816174455744203|11|1
35.059823|195a1e5fb2bfa29594a19f221c5fa1a0e5338de3|1.69|2014-09-13 16:33:00|1.4091206135396188|2|4900000044|66|0.6119093465164359|0|47|54|-80.816172|8|35.059823|DIET|0.0|23|CB COKE ZERO 20 OZ|5d9fb253b347a91c85cbb997da7014c4e3bd9b98|0.6518340734283655|0.61242566243833529|00049000040869|CARBONATED BEVERAGES|BEVERAGE|-80.816172|1.4105082902580508|66|1
35.059823|d4a626a761727e52d5ae7918dc5fbf26a46a4e14|1.69|2014-10-10 10:30:00|1.4091206135396188|2|4900000044|66|0.6119093465164359|0|47|54|-80.816172|8|35.059823|DIET|0.0|23|CB COKE ZERO 20 OZ|5d9fb253b347a91c85cbb997da7014c4e3bd9b98|0.6518340734283655|0.61242566243833529|00049000040869|CARBONATED BEVERAGES|BEVERAGE|-80.816172|1.4105082902580508|66|1
35.059823|a22a8e6ad686857fc11d44105f81ad043e5e6783|4.89|2014-10-02 14:04:00|1.4091206135396188|2|7203660021|66|0.6119093465164359|0|47|355|-80.816172|104|35.059823|FRESH GRILLING SAUSAGE|0.0|19|HT GROUND SAUSAGE MILD|5d9fb253b347a91c85cbb997da7014c4e3bd9b98|0.6518340734283655|0.61242566243833529|00072036600264|DINNER SAUSAGE|CASE READY MEATS|-80.816172|1.4105082902580508|66|1
35.059823|532d79270ffaab8d853dc6e193128ba6cd1d2ad9|1.98|2014-10-01 19:33:00|1.4091206135396188|2|3400000031|66|0.6119093465164359|0|47|47|-80.816172|7|35.059823|REGISTER BARS|0.49|1|(FE)REESE'S NUTRAGEOUS BAR|5d9fb253b347a91c85cbb997da7014c4e3bd9b98|0.6518340734283655|0.61242566243833529|00034000000050|CANDY|G1 GROCERY|-80.816172|1.4105082902580508|66|2
35.059823|09607b4d146d407c6e32639881b873524fabb47c|1.99|2014-09-19 14:02:00|80.816179662140996|2|2840003912|66|35.069256528795776|0|41|206|-80.848528|31|35.053394|FRONT END SNACKS|0.0|1|FRITO LAY CASHEWS|5d9fb253b347a91c85cbb997da7014c4e3bd9b98|0.6518340734283655|35.070508771677183|00028400039123|SNACKS|G1 GROCERY|-80.816172|80.816174455744203|11|1
35.059823|785349c356dd3278a01e55a44ed2902d41c89a00|2.99|2014-09-16 20:05:00|1.4091206135396188|2|7203636062|66|0.6119093465164359|0|47|31|-80.816172|4|35.059823|NON CARBONATED WATER|0.0|1|HT NATURAL SPRING WATER|5d9fb253b347a91c85cbb997da7014c4e3bd9b98|0.6518340734283655|0.61242566243833529|00072036360663|BOTTLED WATER|G1 GROCERY|-80.816172|1.4105082902580508|66|1
35.059823|d7b2b229f44638183add09690209ace19dfecf19|5.97|2014-09-12 20:05:00|1.4091206135396188|2|7203676359|66|0.6119093465164359|0|47|345|-80.816172|57|35.059823|ORGANIC MILK|0.0|3|HTO ORGANIC WHOLE MILK GAL|5d9fb253b347a91c85cbb997da7014c4e3bd9b98|0.6518340734283655|0.61242566243833529|00072036763594|MILK|DAIRY|-80.816172|1.4105082902580508|66|1
35.116751|cb6b2aca748e0cd4bd98b1994623d9129b398779|1.69|2015-02-21 12:41:00|80.825044058860698|4|4900000044|294|35.132488594128802|0|29|54|-80.844274|8|35.204336|DIET|0.0|23|CB DIET COKE CONTOUR 20 OZ NR|5e74f6152deccca1dc4f3e9592cecd37cc5bc3b8|1.0874301175903438|35.157881615307893|00049000000450|CARBONATED BEVERAGES|BEVERAGE|-80.824767|80.824782834502798|61|1
35.141204|ee9b7b3d5998cbda4d4442d60e7fe7414dfa3362|5.98|2014-12-09 16:54:00|80.739023103730261|4|1600081341|171|35.163057780515956|0|16|8|-80.66939|2|35.28326|BROWNIE MIXES|0.99|1|BC WALNUT BROWNIE MIX|5e9c901adb2468cb8dbee345ee0c25101fd986b0|1.5100458916245902|35.169056414731678|00016000813410|BAKING MIXES|G1 GROCERY|-80.739|80.739047979970366|46|2
34.937113|b17528837cfb82924eb5e0818ead22d08f746925|15.49|2015-02-06 15:55:00|1.41290891556208|2|30187136703|372|0.6097676529913135|0|33|3255|-80.837892|1020|34.937113|FACIAL LOTION|0.0|17|L'CERAVE FACIAL MOISTURIZER AM|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00301871366036|FACIAL CLEANSER & MOISTURIZER|HBC|-80.837892|1.4108873757715839|372|1
34.937113|45c72b67e171770e2457a39d9117ac871bb78a65|17.31|2014-12-06 09:53:00|1.41290891556208|2|20188000000|372|0.6097676529913135|0|33|299|-80.837892|49|34.937113|ANGUS BEEF|0.0|2|ANGUS BEEF BNLS CHUCK ROAST|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00201880000009|BEEF|MEAT|-80.837892|1.4108873757715839|372|1
34.937113|c991d25643ca73824b37295fe7d9c8d183c3fcce|18.45|2015-01-10 09:57:00|1.41290891556208|2|20188000000|372|0.6097676529913135|0|33|299|-80.837892|49|34.937113|ANGUS BEEF|6.16|2|ANGUS BEEF BNLS CHUCK ROAST|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00201880000009|BEEF|MEAT|-80.837892|1.4108873757715839|372|1
34.937113|336fc48a534ef6b948e4b3909cfe45d99eb6f909|16.47|2015-03-07 09:49:00|1.41290891556208|2|20188000000|372|0.6097676529913135|0|33|299|-80.837892|49|34.937113|ANGUS BEEF|0.0|2|ANGUS BEEF BNLS CHUCK ROAST|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00201880000009|BEEF|MEAT|-80.837892|1.4108873757715839|372|1
34.937113|4ac9985bc75e1c728a5896b4eaaad6a913b286e7|18.69|2014-12-20 10:03:00|1.41290891556208|2|20188000000|372|0.6097676529913135|0|33|299|-80.837892|49|34.937113|ANGUS BEEF|0.0|2|ANGUS BEEF BNLS CHUCK ROAST|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00201880000009|BEEF|MEAT|-80.837892|1.4108873757715839|372|1
34.937113|839966d2a99da70087118886d3fd4084d69d1e66|2.19|2015-02-26 17:49:00|1.41290891556208|2|7203656071|372|0.6097676529913135|0|33|316|-80.837892|52|34.937113|CREAM CHEESE|0.69|3|HT STAWBERRY CREAM CHEESE|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00072036559982|CHEESE|DAIRY|-80.837892|1.4108873757715839|372|1
34.937113|daff2fb6fe93ce758108d5d98e7a3ed365bfa3d0|3.79|2015-03-09 18:35:00|1.41290891556208|2|3700034885|372|0.6097676529913135|0|33|425|-80.837892|72|34.937113|NFS-PAPER NAPKINS|1.29|1|BOUNTY QUILTED NAPKINS 200CT|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00037000348856|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.837892|1.4108873757715839|372|1
34.937113|3abac4d48a33ae713af9e259e85d67a643e1aa43|1.79|2014-10-08 14:37:00|1.41290891556208|2|4100000362|372|0.6097676529913135|0|33|213|-80.837892|33|34.937113|SOUP MIXES|0.0|1|LIPTON ONION SOUP & DIP MIX|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00041000003622|SOUP|G1 GROCERY|-80.837892|1.4108873757715839|372|1
34.937113|3a56774fcc6dd842dc5ff6495569407f3d985092|1.79|2014-11-22 09:58:00|1.41290891556208|2|4100000362|372|0.6097676529913135|0|33|213|-80.837892|33|34.937113|SOUP MIXES|0.29|1|LIPTON ONION SOUP & DIP MIX|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00041000003622|SOUP|G1 GROCERY|-80.837892|1.4108873757715839|372|1
34.937113|44d78eec1d926581a250a5aa460011664a7376dc|3.79|2014-12-04 09:20:00|1.41290891556208|2|3700034885|372|0.6097676529913135|0|33|425|-80.837892|72|34.937113|NFS-PAPER NAPKINS|1.29|1|BOUNTY QUILTED NAPKINS 200CT|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00037000348856|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.837892|1.4108873757715839|372|1
34.937113|5d62ff05f3c9f7bdb9870acc13cd62bfe5c65c5d|4.97|2014-12-14 09:02:00|1.41290891556208|2|4127102450|372|0.6097676529913135|0|33|341|-80.837892|57|34.937113|CREAMERS|0.0|3|ITNAT'L DELIGHT SF FRENCH VAN|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00041271005073|MILK|DAIRY|-80.837892|1.4108873757715839|372|1
34.937113|8c778a731e92ffdd0c85f6a5f79e7be1d2085391|4.15|2014-11-01 09:35:00|1.41290891556208|2|4400000488|372|0.6097676529913135|0|33|89|-80.837892|12|34.937113|GRAHAM CRACKERS|0.65|1|HONEYMAID GRAHAMS|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00044000004637|COOKIES|G1 GROCERY|-80.837892|1.4108873757715839|372|1
34.937113|fb070cfd712eda2dc131b9b30173cca4f36c68f7|4.15|2014-12-07 11:11:00|1.41290891556208|2|4400000488|372|0.6097676529913135|0|33|89|-80.837892|12|34.937113|GRAHAM CRACKERS|0.65|1|HONEYMAID FRESH STACKS|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00044000026820|COOKIES|G1 GROCERY|-80.837892|1.4108873757715839|372|1
34.937113|61f8bb9e015af0fc533ca3a7eafaf43d40f57d25|4.99|2014-10-05 17:19:00|1.41290891556208|2|4242116078|372|0.6097676529913135|0|33|1855|-80.837892|430|34.937113|BH SALAMI/CHUBBS|1.0|6|BOARS HEAD PEPPERONI NC STICK|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00042421160789|SPECIALTY MEAT|DELI|-80.837892|1.4108873757715839|372|1
34.937113|6496a5b8e7b21fa511fd6e45bb515d7aae67293b|1.75|2014-09-26 14:11:00|1.41290891556208|2|96824|372|0.6097676529913135|0|33|1581|-80.837892|369|34.937113|NFS BEVERAGE BREWED|0.0|22|BREWED  COFFEE TALL.|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00000000968240|NFS STARBUCKS|COFFEE SHOP|-80.837892|1.4108873757715839|372|1
34.937113|9ff2f4884d7630685b2360cc3006d6a8ddf1029b|5.5|2014-12-01 16:26:00|1.41290891556208|2|930018709|372|0.6097676529913135|0|33|162|-80.837892|25|34.937113|PICKLES|0.0|1|MT OLV SPEAR KOSHER DILL FP|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00009300000802|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.837892|1.4108873757715839|372|2
34.937113|713fb28c6fb1f71eef93c8bcb34064fa07509736|5.29|2015-02-01 13:48:00|1.41290891556208|2|5150024177|372|0.6097676529913135|0|33|125|-80.837892|19|34.937113|PEANUT BUTTER|0.0|1|JIF CREAMY PEANUT BUTTER|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00051500241776|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.837892|1.4108873757715839|372|1
34.937113|7bb9ba1e0c354e9a15b75ccc411bbb3f48d0ac37|5.29|2015-01-25 15:43:00|1.41290891556208|2|5150024177|372|0.6097676529913135|0|33|125|-80.837892|19|34.937113|PEANUT BUTTER|0.0|1|JIF CREAMY PEANUT BUTTER|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00051500241776|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.837892|1.4108873757715839|372|1
34.937113|7e50af78bbe4754f5d6a22f2c6df8f7feca0017c|5.29|2014-11-09 15:02:00|1.41290891556208|2|5150024177|372|0.6097676529913135|0|33|125|-80.837892|19|34.937113|PEANUT BUTTER|1.3|1|JIF CREAMY PEANUT BUTTER|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00051500241776|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.837892|1.4108873757715839|372|1
34.937113|8f2302a019cb206491c630298f56bd88eaa1e44c|0.6|2014-09-17 13:58:00|1.41290891556208|2|5000000124|372|0.6097676529913135|0|33|154|-80.837892|24|34.937113|NFS-CAT FOOD WET|0.0|1|FANCY FEAST DELIGHTS TRKY&CHS|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00050000585489|PET FOOD/SUPPLIES|G1 GROCERY|-80.837892|1.4108873757715839|372|1
34.937113|72bbfb0611291f3cc0ba199ce0cbad6c3a8b0040|0.55|2015-01-18 14:10:00|1.41290891556208|2|5000000124|372|0.6097676529913135|0|33|154|-80.837892|24|34.937113|NFS-CAT FOOD WET|0.05|1|FANCY FEAST DELIGHTS CHK&CHS|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00050000585434|PET FOOD/SUPPLIES|G1 GROCERY|-80.837892|1.4108873757715839|372|1
34.937113|942c7a087132304cd9dfc8d7e359e7f709712a02|1.39|2014-10-10 15:28:00|1.41290891556208|2|5210076069|372|0.6097676529913135|0|33|80|-80.837892|34|34.937113|SEASONING PACKETS|0.0|1|MC GRILL MATES MESQUITE MARNDE|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00052100025780|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.837892|1.4108873757715839|372|1
34.937113|d860c6850cc14f43ad761c59eeadbb388f9d148b|2.79|2014-11-24 14:00:00|1.41290891556208|2|5150024136|372|0.6097676529913135|0|33|125|-80.837892|19|34.937113|PEANUT BUTTER|0.0|1|JIF TO GO 8 PK|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00051500241363|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.837892|1.4108873757715839|372|1
34.937113|3761a4ad90b8635a8d48cc3e737e71c46fb5cb8b|0.55|2015-03-02 18:04:00|1.41290891556208|2|5000000124|372|0.6097676529913135|0|33|154|-80.837892|24|34.937113|NFS-CAT FOOD WET|0.0|1|FANCY FEAST GOURMET CHICKEN|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00050000429943|PET FOOD/SUPPLIES|G1 GROCERY|-80.837892|1.4108873757715839|372|1
34.937113|c7f3b0fc4769237976cd6d42ec4df5339f42f6a9|1.1|2015-02-11 15:23:00|1.41290891556208|2|5000000124|372|0.6097676529913135|0|33|154|-80.837892|24|34.937113|NFS-CAT FOOD WET|0.0|1|FANCY FEAST BEEF/CHICKEN|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00050000429745|PET FOOD/SUPPLIES|G1 GROCERY|-80.837892|1.4108873757715839|372|2
34.937113|c28a792ea3230016e14a14949db4daf85d336f92|0.55|2015-01-20 14:34:00|80.762257539052428|2|5000000124|372|34.954807759443746|0|54|154|-80.847383|24|35.024464|NFS-CAT FOOD WET|0.05|1|FANCY FEAST BEEF/CHICKEN|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|34.983028186791387|00050000429745|PET FOOD/SUPPLIES|G1 GROCERY|-80.837892|80.837910724874504|317|1
34.937113|5f8d5741b6edb0adc4eec2920e1d35c704fc9af8|0.55|2014-11-05 14:45:00|80.762257539052428|2|5000000124|372|34.954807758683685|0|54|154|-80.850065|24|35.030252|NFS-CAT FOOD WET|0.0|1|FANCY FEAST SEAFOOD FEAST|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|34.983028186791387|00050000429349|PET FOOD/SUPPLIES|G1 GROCERY|-80.837892|80.837911764959472|470|1
34.937113|0bfd3642edd3735b4c34929bb5522b8ca922a7f2|0.55|2014-10-31 17:08:00|80.762257539052428|2|5000000124|372|34.954807758683685|0|54|154|-80.850065|24|35.030252|NFS-CAT FOOD WET|0.0|1|FANCY FEAST SAVORY SALMON|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|34.983028186791387|00050000429448|PET FOOD/SUPPLIES|G1 GROCERY|-80.837892|80.837911764959472|470|1
34.937113|e7478641b1a13951b45b5d13ec9ecb570a4fcf1b|0.99|2014-09-28 11:58:00|1.41290891556208|2|87694000301|372|0.6097676529913135|0|33|154|-80.837892|24|34.937113|NFS-CAT FOOD WET|0.09|1|VARIETY PET SALMON CASSEROLE|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00876940003063|PET FOOD/SUPPLIES|G1 GROCERY|-80.837892|1.4108873757715839|372|1
34.937113|cb96edb186289744d63631cb7b2c4b60a4bb2e28|3.58|2014-12-22 08:32:00|1.41290891556208|2|3600025824|372|0.6097676529913135|0|33|424|-80.837892|72|34.937113|NFS-FACIAL TISSUE|0.0|1|KLEENEX UL FACIAL TISSUE WHITE|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00036000258615|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.837892|1.4108873757715839|372|2
34.937113|27e8a6c558d8d2e814d64d7b6184ec8d392115c2|3.58|2015-01-30 15:27:00|1.41290891556208|2|3600025824|372|0.6097676529913135|0|33|424|-80.837892|72|34.937113|NFS-FACIAL TISSUE|0.0|1|KLEENEX UL FACIAL TISSUE WHITE|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00036000258615|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.837892|1.4108873757715839|372|2
34.937113|e520bc5dc2f13bc62d5d6b64eeb893392347cd38|5.37|2015-01-14 10:47:00|1.41290891556208|2|3600025824|372|0.6097676529913135|0|33|424|-80.837892|72|34.937113|NFS-FACIAL TISSUE|0.0|1|KLEENEX UL FACIAL TISSUE WHITE|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00036000258615|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.837892|1.4108873757715839|372|3
34.937113|54aec0b2627c46b4884aaa787f6982e3dcd4d255|3.58|2014-12-17 16:34:00|1.41290891556208|2|3600025824|372|0.6097676529913135|0|33|424|-80.837892|72|34.937113|NFS-FACIAL TISSUE|0.0|1|KLEENEX UL FACIAL TISSUE WHITE|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00036000258615|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.837892|1.4108873757715839|372|2
34.937113|2b97ebaaf786cab31375879adbdd4ba84a97fbe9|5.0|2014-11-19 15:43:00|1.41290891556208|2|3600025824|372|0.6097676529913135|0|33|424|-80.837892|72|34.937113|NFS-FACIAL TISSUE|0.42|1|KLEENEX UL FACIAL TISSUE WHITE|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00036000258615|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.837892|1.4108873757715839|372|3
34.937113|6c8fae27295701ca51b222e091cd108b2635c956|1.79|2015-02-23 18:35:00|1.41290891556208|2|3600025824|372|0.6097676529913135|0|33|424|-80.837892|72|34.937113|NFS-FACIAL TISSUE|0.0|1|KLEENEX UL FACIAL TISSUE WHITE|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00036000258615|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.837892|1.4108873757715839|372|1
34.937113|3f3badbf2a976daf6dfc7c30269ad6965c7c70f7|2.99|2014-10-27 14:48:00|1.41290891556208|2|4200035501|372|0.6097676529913135|0|33|425|-80.837892|72|34.937113|NFS-PAPER NAPKINS|0.0|1|VANITY FAIR FOLDED NAPKIN|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00042000355094|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.837892|1.4108873757715839|372|1
34.937113|1a0f5727e72ba3ab29901d096d289621104f334f|10.49|2015-03-06 10:44:00|1.41290891556208|2|7365111723|372|0.6097676529913135|0|33|160|-80.837892|25|34.937113|OLIVES|1.5|1|MARIO OLIVE QUEEN 21 OZ|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00073651117236|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.837892|1.4108873757715839|372|1
34.937113|c61c2cb2bcf8339ddab084c7710e259f7c0362aa|10.49|2014-12-17 13:27:00|1.41290891556208|2|7365111723|372|0.6097676529913135|0|33|160|-80.837892|25|34.937113|OLIVES|1.5|1|MARIO OLIVE QUEEN 21 OZ|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00073651117236|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.837892|1.4108873757715839|372|1
34.937113|4a6c96f5ce5e87a58e16af892c89a360e02cf448|1.15|2015-01-04 09:19:00|1.41290891556208|2|7203663222|372|0.6097676529913135|0|33|330|-80.837892|55|34.937113|EGGS|0.0|3|HT GRADE A    LARGE EGGS 6 CT.|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00072036632227|EGGS FRESH|DAIRY|-80.837892|1.4108873757715839|372|1
34.937113|deec35effbe55ccb381da7b05d83bbeb0c5a5226|2.19|2014-09-12 15:30:00|1.41290891556208|2|7203670343|372|0.6097676529913135|0|33|443|-80.837892|76|34.937113|NFS-GARBAGE BAGS|0.41|1|YH SML GARBAGE ODOR CNT|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00072036703507|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.837892|1.4108873757715839|372|1
34.937113|9aed5e204655ede4a65e6d33cbe5ea889dcdf2fc|0.85|2014-09-15 15:47:00|1.41290891556208|2|7203663222|372|0.6097676529913135|0|33|330|-80.837892|55|34.937113|EGGS|0.0|3|HT GRADE A    LARGE EGGS 6 CT.|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00072036632227|EGGS FRESH|DAIRY|-80.837892|1.4108873757715839|372|1
34.937113|e59370d855ff0123019e966c99004e2b1f0e3f99|9.99|2014-12-15 15:07:00|1.41290891556208|2|8520000062|372|0.6097676529913135|0|33|9933|-80.837892|884|34.937113|NFS FV OTHER WHITE|0.0|13|SUTTER HOME MOSCATO 1.5L|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00085200000623|FIGHTING VARIETL($0-$3.99)|WINE|-80.837892|1.4108873757715839|372|1
34.937113|0b3eeaf0e20aa7fdbeed28d3d37ba91246f3d996|14.99|2014-10-25 19:07:00|1.41290891556208|2|8500000653|372|0.6097676529913135|0|33|9925|-80.837892|883|34.937113|NFS-ECONOMY GLASS|0.0|13|LIVINGSTON RED ROSE 3L|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00085000006535|ECONOMY (GLASS 3L & UP)|WINE|-80.837892|1.4108873757715839|372|1
34.937113|88ae2c8f00d506dc3257c7610cfe1610ff403735|0.64|2014-09-21 15:42:00|1.41290891556208|2||372|0.6097676529913135|0|33|502|-80.837892|64|34.937113|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00204011000008|FRESH PRODUCE|PRODUCE|-80.837892|1.4108873757715839|372|1
34.937113|109e4a9654d24c7eeca5b57c537e2878722d0aa6|0.53|2015-01-08 16:14:00|1.41290891556208|2||372|0.6097676529913135|0|33|502|-80.837892|64|34.937113|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00204011000008|FRESH PRODUCE|PRODUCE|-80.837892|1.4108873757715839|372|1
34.937113|2f3b7b2b60103cec289b321cf345f34b673b98ad|0.61|2014-10-14 13:36:00|1.41290891556208|2||372|0.6097676529913135|0|33|502|-80.837892|64|34.937113|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00204011000008|FRESH PRODUCE|PRODUCE|-80.837892|1.4108873757715839|372|1
34.937113|d2f4d9b8f8931eb30e61ac4a09d41d6c14129cdc|0.58|2014-11-11 13:06:00|80.762257539052428|2||372|34.954807759443746|0|54|502|-80.847383|64|35.024464|FRESH BANANAS|0.0|4|BANANAS, YELLOW|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|34.983028186791387|00204011000008|FRESH PRODUCE|PRODUCE|-80.837892|80.837910724874504|317|1
34.937113|9bb998cb801c3d91f4ec0424cac5470d09a461f2|4.89|2014-11-01 18:01:00|1.41290891556208|2|7365111741|372|0.6097676529913135|0|33|160|-80.837892|25|34.937113|OLIVES|0.0|1|MARIO OLIVE QUEEN STFD PIM|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00073651117410|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.837892|1.4108873757715839|372|1
34.937113|db16f9bb3048e73b3e397487f2f7f09e2c0dd86d|22.93|2014-10-11 09:41:00|1.41290891556208|2|20898900000|372|0.6097676529913135|0|33|1421|-80.837892|201|34.937113|SMART CHICKEN VEGETABLE FED|0.0|2|SMART CHICKEN BONELESS BREAST|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00208989000008|POULTRY|MEAT|-80.837892|1.4108873757715839|372|2
34.937113|9c6cde6ba5fc6aada8aa79120b527ab1c7f25567|9.98|2015-02-25 15:35:00|1.41290891556208|2|20898900000|372|0.6097676529913135|0|33|1421|-80.837892|201|34.937113|SMART CHICKEN VEGETABLE FED|0.0|2|SMART CHICKEN BONELESS BREAST|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00208989000008|POULTRY|MEAT|-80.837892|1.4108873757715839|372|1
34.937113|16cf6349fdc32e09e94a4fc2e7a0d2fea473c27a|5.19|2014-11-15 09:40:00|1.41290891556208|2|20165500000|372|0.6097676529913135|0|33|297|-80.837892|49|34.937113|GROUND BEEF|0.0|2|HT PREMIUM GRND BEEF 80% LEAN|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00201655000005|BEEF|MEAT|-80.837892|1.4108873757715839|372|1
34.937113|de75a3bc7cb9b4c0973e87350039f20791b5b6cd|2.49|2014-09-24 15:35:00|1.41290891556208|2|7878350610|372|0.6097676529913135|0|33|527|-80.837892|64|34.937113|FRESH CARROTS|0.0|4|MATCHSTICK CARROTS, PKG|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00078783506101|FRESH PRODUCE|PRODUCE|-80.837892|1.4108873757715839|372|1
34.937113|eefa649f29a88022d2d196ea12d6a38a85dca3e5|8.89|2015-02-04 14:20:00|80.762257539052428|2|515|372|34.954807758683685|0|54|33|-80.850065|10|35.030252|COFFEE BULK|0.0|1|HT TRADER BULK COFFEE PLU|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|34.983028186791387|00000000005150|COFFEE|G1 GROCERY|-80.837892|80.837911764959472|470|1
34.937113|b2036e1a11c662faf9771f41c7274d34d44ae858|6.5|2015-01-07 14:12:00|80.762257539052428|2|4127102564|372|34.954807758683685|0|54|341|-80.850065|57|35.030252|CREAMERS|0.96|3|ITNAT'L SF FRENCH VANILLA|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|34.983028186791387|00041271025057|MILK|DAIRY|-80.837892|80.837911764959472|470|2
34.937113|de4053fd384328c5fb63f764bd4ed17feaf08e16|3.15|2014-09-26 14:08:00|1.41290891556208|2|4127102564|372|0.6097676529913135|0|33|341|-80.837892|57|34.937113|CREAMERS|0.0|3|ITNAT'L SF FRENCH VANILLA|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00041271025057|MILK|DAIRY|-80.837892|1.4108873757715839|372|1
34.937113|d0921c08307eea50ac236d21eea5e3bdff787eb7|3.25|2015-02-09 18:02:00|1.41290891556208|2|4127102564|372|0.6097676529913135|0|33|341|-80.837892|57|34.937113|CREAMERS|0.48|3|ITNAT'L SF FRENCH VANILLA|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00041271025057|MILK|DAIRY|-80.837892|1.4108873757715839|372|1
34.937113|f8585d7918d8b3e6a0f31b45afb985a009261f40|3.25|2015-03-05 15:38:00|1.41290891556208|2|4127102564|372|0.6097676529913135|0|33|341|-80.837892|57|34.937113|CREAMERS|1.26|3|ITNAT'L SF FRENCH VANILLA|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00041271025057|MILK|DAIRY|-80.837892|1.4108873757715839|372|1
34.937113|1953eb1accd08ffe1d8c2414c2000e8a21c3c62c|3.49|2014-10-01 14:09:00|1.41290891556208|2|4127102564|372|0.6097676529913135|0|33|341|-80.837892|57|34.937113|CREAMERS|0.49|3|ITNAT'L SF FRENCH VANILLA|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00041271025057|MILK|DAIRY|-80.837892|1.4108873757715839|372|1
34.937113|a6c09ecc50e0b1f347d319236ad4e1768029b634|3.0|2014-09-13 08:08:00|1.41290891556208|2|76211193803|372|0.6097676529913135|0|33|1598|-80.837892|369|34.937113|NFS MERCHANDISE|0.0|22|REUSABLE CUP 16OZ|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00762111938039|NFS STARBUCKS|COFFEE SHOP|-80.837892|1.4108873757715839|372|3
34.937113|1e0c5beb6e24f78256817151e877f040d526d6ad|4.45|2014-11-07 14:42:00|1.41290891556208|2|96974|372|0.6097676529913135|0|33|1597|-80.837892|369|34.937113|NFS BEVERAGE BLEND|0.0|22|CARAMEL FRAPPUCCINO GRANDE|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00000000969740|NFS STARBUCKS|COFFEE SHOP|-80.837892|1.4108873757715839|372|1
34.937113|8032b9715bb2ec2ce15034560ab84b255f26219c|4.45|2014-10-08 18:38:00|1.41290891556208|2|96974|372|0.6097676529913135|0|33|1597|-80.837892|369|34.937113|NFS BEVERAGE BLEND|0.0|22|CARAMEL FRAPPUCCINO GRANDE|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00000000969740|NFS STARBUCKS|COFFEE SHOP|-80.837892|1.4108873757715839|372|1
34.937113|aefc6246edd41e232acd80da3de057062da41cd3|4.45|2014-10-29 18:34:00|1.41290891556208|2|96974|372|0.6097676529913135|0|33|1597|-80.837892|369|34.937113|NFS BEVERAGE BLEND|1.45|22|CARAMEL FRAPPUCCINO GRANDE|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00000000969740|NFS STARBUCKS|COFFEE SHOP|-80.837892|1.4108873757715839|372|1
34.937113|a13e1cee6e558cc6dc277a8947567aa67a3a73ff|4.45|2015-01-21 18:31:00|1.41290891556208|2|96974|372|0.6097676529913135|0|33|1597|-80.837892|369|34.937113|NFS BEVERAGE BLEND|0.0|22|CARAMEL FRAPPUCCINO GRANDE|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00000000969740|NFS STARBUCKS|COFFEE SHOP|-80.837892|1.4108873757715839|372|1
34.937113|36115379a5678a1e8f759351f0f946a0a068e096|1.94|2014-12-10 13:07:00|1.41290891556208|2|7203698758|372|0.6097676529913135|0|33|31|-80.837892|4|34.937113|NON CARBONATED WATER|0.0|1|HT SPRING WATER|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00072036987587|BOTTLED WATER|G1 GROCERY|-80.837892|1.4108873757715839|372|2
34.937113|c3091f77181ec57675ac436dcbed1d7f9c16a9e3|3.58|2015-02-07 09:43:00|1.41290891556208|2||372|0.6097676529913135|0|33|540|-80.837892|64|34.937113|FRESH CELERY|0.0|4|COO CELERY (RPC) 24'S|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00204070000001|FRESH PRODUCE|PRODUCE|-80.837892|1.4108873757715839|372|2
34.937113|ce137cb4040433adb6fe69386f55b55afbdbd341|2.75|2014-10-11 08:10:00|1.41290891556208|2|96326|372|0.6097676529913135|0|33|1599|-80.837892|370|34.937113|PASTRY|0.0|22|BOWL OF OATMEAL|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00000000963260|STARBUCKS|COFFEE SHOP|-80.837892|1.4108873757715839|372|1
34.937113|3b0d9b919664f6168d3a1f13bb06df0e49970c20|2.75|2014-09-27 08:06:00|1.41290891556208|2|96326|372|0.6097676529913135|0|33|1599|-80.837892|370|34.937113|PASTRY|0.0|22|BOWL OF OATMEAL|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00000000963260|STARBUCKS|COFFEE SHOP|-80.837892|1.4108873757715839|372|1
34.937113|79d4a4e8b52e6fd25b0ef54c3fca37043e47d831|4.19|2015-01-03 15:21:00|1.41290891556208|2|1600027578|372|0.6097676529913135|0|33|61|-80.837892|9|34.937113|RTE CEREAL ADULT|0.0|1|FIBER ONE CEREAL|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00016000275058|CEREAL|G1 GROCERY|-80.837892|1.4108873757715839|372|1
34.937113|6fb216d4fd5348801a598f06f22a52ba3e1e285a|2.35|2014-11-22 07:41:00|1.41290891556208|2|96826|372|0.6097676529913135|0|33|1581|-80.837892|369|34.937113|NFS BEVERAGE BREWED|0.0|22|BREWED COFFEE VENTI|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00000000968260|NFS STARBUCKS|COFFEE SHOP|-80.837892|1.4108873757715839|372|1
34.937113|bdcfc5cd5071bf27fc7f7d0e1344416b41f97a07|2.35|2015-01-10 07:43:00|1.41290891556208|2|96826|372|0.6097676529913135|0|33|1581|-80.837892|369|34.937113|NFS BEVERAGE BREWED|0.0|22|BREWED COFFEE VENTI|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00000000968260|NFS STARBUCKS|COFFEE SHOP|-80.837892|1.4108873757715839|372|1
34.937113|21040c58ae98dbb191965c9095e82df6511001ca|2.35|2015-01-31 07:48:00|1.41290891556208|2|96826|372|0.6097676529913135|0|33|1581|-80.837892|369|34.937113|NFS BEVERAGE BREWED|0.0|22|BREWED COFFEE VENTI|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00000000968260|NFS STARBUCKS|COFFEE SHOP|-80.837892|1.4108873757715839|372|1
34.937113|348147550096862450d106076dafb512a3b0528a|2.35|2014-11-01 07:49:00|1.41290891556208|2|96826|372|0.6097676529913135|0|33|1581|-80.837892|369|34.937113|NFS BEVERAGE BREWED|0.0|22|BREWED COFFEE VENTI|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00000000968260|NFS STARBUCKS|COFFEE SHOP|-80.837892|1.4108873757715839|372|1
34.937113|527bce209c27300c2a58afeed9a59c062b704c85|2.35|2014-12-06 07:41:00|1.41290891556208|2|96826|372|0.6097676529913135|0|33|1581|-80.837892|369|34.937113|NFS BEVERAGE BREWED|0.0|22|BREWED COFFEE VENTI|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00000000968260|NFS STARBUCKS|COFFEE SHOP|-80.837892|1.4108873757715839|372|1
34.937113|01fbe0773577633923b4428dacc53d49a8582110|2.35|2014-12-20 07:49:00|1.41290891556208|2|96826|372|0.6097676529913135|0|33|1581|-80.837892|369|34.937113|NFS BEVERAGE BREWED|0.0|22|BREWED COFFEE VENTI|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00000000968260|NFS STARBUCKS|COFFEE SHOP|-80.837892|1.4108873757715839|372|1
34.937113|ddf88b769577f17593afdc4779a753813ea71481|2.35|2014-11-08 08:06:00|1.41290891556208|2|96826|372|0.6097676529913135|0|33|1581|-80.837892|369|34.937113|NFS BEVERAGE BREWED|0.0|22|BREWED COFFEE VENTI|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00000000968260|NFS STARBUCKS|COFFEE SHOP|-80.837892|1.4108873757715839|372|1
34.937113|dc9e000eb92b578e45c29aae04debd0f56a452bc|2.35|2015-03-07 08:07:00|1.41290891556208|2|96826|372|0.6097676529913135|0|33|1581|-80.837892|369|34.937113|NFS BEVERAGE BREWED|0.0|22|BREWED COFFEE VENTI|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00000000968260|NFS STARBUCKS|COFFEE SHOP|-80.837892|1.4108873757715839|372|1
34.937113|cc9e76441b80f06b92417da69cad6f4a0a6535bb|2.35|2014-11-15 07:40:00|1.41290891556208|2|96826|372|0.6097676529913135|0|33|1581|-80.837892|369|34.937113|NFS BEVERAGE BREWED|0.0|22|BREWED COFFEE VENTI|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00000000968260|NFS STARBUCKS|COFFEE SHOP|-80.837892|1.4108873757715839|372|1
34.937113|76a5db39974a3f7a3bd32d3959d2394de62411b4|12.59|2014-10-29 16:07:00|1.41290891556208|2|73221630004|372|0.6097676529913135|0|33|4195|-80.837892|1200|34.937113|COUGH & COLD REMEDY-ADULT|0.0|17|ZICAM COLD RM CHRY-30004|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00732216300048|COUGH/COLD/SINUS|HBC|-80.837892|1.4108873757715839|372|1
34.937113|54e573342c933b4515ad2d54fad71a86866f4376|4.45|2015-03-09 18:38:00|1.41290891556208|2|97078|372|0.6097676529913135|0|33|1597|-80.837892|369|34.937113|NFS BEVERAGE BLEND|0.0|22|CARAMEL LIGHT FRAPP GRANDE|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00000000970780|NFS STARBUCKS|COFFEE SHOP|-80.837892|1.4108873757715839|372|1
34.937113|7c3c27149c7c265ee891f07ded8cbcf855ac66a1|4.45|2014-12-10 13:10:00|1.41290891556208|2|97078|372|0.6097676529913135|0|33|1597|-80.837892|369|34.937113|NFS BEVERAGE BLEND|0.0|22|CARAMEL LIGHT FRAPP GRANDE|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00000000970780|NFS STARBUCKS|COFFEE SHOP|-80.837892|1.4108873757715839|372|1
34.937113|2312a59347fff7e8138999aa286868a06ff9f3c5|3.95|2015-02-07 07:46:00|1.41290891556208|2|96973|372|0.6097676529913135|0|33|1597|-80.837892|369|34.937113|NFS BEVERAGE BLEND|0.0|22|CARAMEL FRAPPUCCINO TALL|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|0.61055446569467375|00000000969730|NFS STARBUCKS|COFFEE SHOP|-80.837892|1.4108873757715839|372|1
34.937113|b3afebe7d765b1492f06dab384b28d58b43273a0|12.850000000000001|2014-12-19 17:41:00|80.762257539052428|2|20169200000|372|34.954807754123038|0|54|297|-80.848528|49|35.053394|GROUND BEEF|0.0|2|GROUND BEEF 96% LEAN|5ea9c0f2503ffdbce025ac723f8bff46271eae64|1.2226656062174164|34.983028186791387|00201692000006|BEEF|MEAT|-80.837892|80.837917117093994|11|2
35.478031|32702db382db4566873d36a273088d70e6160952|1.99|2014-12-28 20:23:00|80.8939826282094|1|7203688096|179|35.491662991994396|0|2|526|-80.8955|64|35.4437|FRESH MUSHROOMS|0.0|4|HT SLICED WHITE MUSHROOMS|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00072036880963|FRESH PRODUCE|PRODUCE|-80.893784|80.893790090795775|272|1
35.478031|a63e2e365e12cb934471bec4931749a77ce68891|1.99|2015-02-11 16:19:00|80.8939826282094|1|7203688096|179|35.491662992623695|0|2|526|-80.861571|64|35.444615|FRESH MUSHROOMS|0.49|4|HT SLICED WHITE MUSHROOMS|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00072036880963|FRESH PRODUCE|PRODUCE|-80.893784|80.893787349746532|340|1
35.478031|b54fa68536d0a11810c4e13874eb493f68f86cc7|1.99|2014-10-28 11:39:00|80.8939826282094|1|7203676415|179|35.491662990721132|0|2|1465|-80.86175|42|35.40953|ORGANIC FROZEN FRUIT|0.0|5|HTO ORGANIC WHOLE MXED BERRIES|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00072036763846|FROZEN FRUIT|FROZEN|-80.893784|80.893793458029279|209|1
35.478031|873526aa82acfcad5fb332bc2108d5ce52cb8d8d|1.99|2015-01-25 17:22:00|80.8939826282094|1|7203688096|179|35.491662991994396|0|2|526|-80.8955|64|35.4437|FRESH MUSHROOMS|0.0|4|HT SLICED WHITE MUSHROOMS|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00072036880963|FRESH PRODUCE|PRODUCE|-80.893784|80.893790090795775|272|1
35.478031|3bde0118d0faaf2220079dc7dbb0945551d7c35f|1.99|2014-11-25 15:53:00|80.8939826282094|1|7203688096|179|35.491662990721132|0|2|526|-80.86175|64|35.40953|FRESH MUSHROOMS|0.2|4|HT SLICED WHITE MUSHROOMS|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00072036880963|FRESH PRODUCE|PRODUCE|-80.893784|80.893793458029279|209|1
35.478031|1cac73251b3ea37e2017a4ddf7e783d0c93a60b1|1.99|2015-03-09 17:03:00|80.8939826282094|1|7203688096|179|35.491662992623695|0|2|526|-80.861571|64|35.444615|FRESH MUSHROOMS|0.0|4|HT SLICED WHITE MUSHROOMS|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00072036880963|FRESH PRODUCE|PRODUCE|-80.893784|80.893787349746532|340|1
35.478031|381094969740bc8cb066dc20a2bcbb4be4faf98d|1.99|2015-02-24 19:52:00|80.8939826282094|1|7203688096|179|35.491662992623695|0|2|526|-80.861571|64|35.444615|FRESH MUSHROOMS|0.0|4|HT SLICED WHITE MUSHROOMS|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00072036880963|FRESH PRODUCE|PRODUCE|-80.893784|80.893787349746532|340|1
35.478031|0c461a55ccf550dee619627eff94e53beeff7253|1.99|2014-09-28 17:33:00|80.8939826282094|1|7203688096|179|35.491662990721132|0|2|526|-80.86175|64|35.40953|FRESH MUSHROOMS|0.49|4|HT SLICED WHITE MUSHROOMS|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00072036880963|FRESH PRODUCE|PRODUCE|-80.893784|80.893793458029279|209|1
35.478031|0acc15abcf6f61077b9f22daf30076cb8a7e48a6|3.85|2014-10-05 20:16:00|80.8939826282094|1|7203663089|179|35.491662990721132|0|2|345|-80.86175|57|35.40953|ORGANIC MILK|0.0|3|HTO ORGANIC CRTN MILK 2%|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00072036630889|MILK|DAIRY|-80.893784|80.893793458029279|209|1
35.478031|efdcfd0b5bf5ad9a91fd6bc96f61b585ff7b2cb4|2.79|2014-09-14 16:06:00|80.8939826282094|1|7203663125|179|35.491662990721132|0|2|1262|-80.86175|57|35.40953|HALF N HALF WHIPPING CREAM|0.0|3|HT HEAVY WHIPPING CREAM|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00072036630988|MILK|DAIRY|-80.893784|80.893793458029279|209|1
35.478031|0701035815ec97f56c1834ab5d833d3f51d45b8b|4.88|2015-02-22 11:19:00|80.8939826282094|1||179|35.491662990721132|0|2|501|-80.86175|64|35.40953|FRESH PEARS|0.0|4|RED PEARS|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00204417000008|FRESH PRODUCE|PRODUCE|-80.893784|80.893793458029279|209|1
35.478031|9ab1f272ca48e0856877c4e5817ac3373158d3f9|2.89|2014-11-09 12:52:00|80.8939826282094|1|7240000720|179|35.491662990721132|0|2|126|-80.86175|19|35.40953|PRESERVES/MARMALADE|0.0|1|POLANER ALL FRUIT STRAWBERRY|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00072400007200|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.893784|80.893793458029279|209|1
35.478031|3c6a700e474e4416aa40b30f8feb645b286781be|7.59|2015-01-21 10:45:00|80.8939826282094|1|7274580478|179|35.491662992623695|0|2|353|-80.861571|110|35.444615|FROZEN CASE MEAT|0.0|19|PERDUE CHICKEN BREAST TENDERS|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00072745804311|FROZEN CASE MEAT|CASE READY MEATS|-80.893784|80.893787349746532|340|1
35.478031|d1f90ec951b344e0e5ec55c170221d51de921ee7|7.59|2014-11-22 14:52:00|80.8939826282094|1|7274580478|179|35.491662990721132|0|2|353|-80.86175|110|35.40953|FROZEN CASE MEAT|0.0|19|PERDUE CHICKEN BREAST PATTIE|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00072745804113|FROZEN CASE MEAT|CASE READY MEATS|-80.893784|80.893793458029279|209|1
35.478031|d131c79f09837376a3af966442abeac079b554b8|4.99|2014-11-17 15:25:00|80.8939826282094|1|71575610004|179|35.491662990721132|0|2|561|-80.86175|64|35.40953|FR PROD ORGANIC PRODUCE|0.0|4|ORG RED RASPBERRIES 6 OZ|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00715756100040|FRESH PRODUCE|PRODUCE|-80.893784|80.893793458029279|209|1
35.478031|882091ebd88fc79035098be3f25145d06a05001f|5.29|2015-01-12 14:05:00|80.8939826282094|1|74236560635|179|35.491662990721132|0|2|332|-80.86175|52|35.40953|STRING/SNACK|1.3|3|HORIZON STRING CHEESE|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00742365606359|CHEESE|DAIRY|-80.893784|80.893793458029279|209|1
35.478031|1fb92776e9802e7381a0b60ed06533dda48952cd|3.29|2015-02-10 10:10:00|80.8939826282094|1|2840018382|179|35.491662992623695|0|2|201|-80.861571|31|35.444615|POTATO CHIPS|0.79|1|BAKED RUFFLES REGULAR|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00028400184793|SNACKS|G1 GROCERY|-80.893784|80.893787349746532|340|1
35.478031|36e0f2c6c4724a22eb3e9fafddb34f6b5b539611|2.99|2015-01-17 17:46:00|80.8939826282094|1|1800000338|179|35.491662991994396|0|2|1268|-80.8955|54|35.4437|BAGELS AND MUFFINS|0.0|3|PILLSBURY READY PIZZA CRUST|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00018000003389|DOUGH PRODUCTS|DAIRY|-80.893784|80.893790090795775|272|1
35.478031|8f3bfcc913e6c8b2c4ae31325f52a3496362dd53|5.98|2014-09-24 18:22:00|80.8939826282094|1|1800000338|179|35.491662990721132|0|2|1268|-80.86175|54|35.40953|BAGELS AND MUFFINS|0.0|3|PILLSBURY READY PIZZA CRUST|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00018000003389|DOUGH PRODUCTS|DAIRY|-80.893784|80.893793458029279|209|2
35.478031|cc86fa8fb995da3f7ba42f77a9cdd294c0976fa2|1.89|2014-11-03 14:19:00|80.8939826282094|1|2000000065|179|35.491662990721132|0|2|1275|-80.86175|50|35.40953|BOX VEG|0.0|5|GG BROCCOLI SPEAR NO SAUCE|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00020000174839|VEGETABLES-FROZEN|FROZEN|-80.893784|80.893793458029279|209|1
35.478031|fbadcbdcdb168a666704c94d9a3a84db0b7d5b83|2.79|2015-02-01 17:32:00|80.8939826282094|1|4133500053|179|35.491662991994396|0|2|184|-80.8955|28|35.4437|SALAD DRESSINGS-LIQUID|0.0|1|KENS DRS CNKY BLUE CHEESE|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00041335001256|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.893784|80.893790090795775|272|1
35.478031|75e554988894ab085a3fb5bdce994d77ad8960ec|6.3|2015-02-08 17:31:00|80.8939826282094|1|7265500105|179|35.491662991994396|0|2|1278|-80.8955|48|35.4437|SINGLE SERVE NUTRITIONAL|1.3|5|HC CAFE STEAMERS BASIL CHICKEN|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00072655001145|FROZEN MEALS|FROZEN|-80.893784|80.893790090795775|272|2
35.478031|a8f791572df829d144d9422771a6a911f6b9f8e5|6.99|2014-12-10 14:47:00|80.8939826282094|1|7790050241|179|35.491662992623695|0|2|1271|-80.861571|41|35.444615|PROTEIN BREAKFAST|0.0|5|J D DL 4CT TSEC FLATBREAD|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00077900650246|BREAKFAST FOODS FROZEN|FROZEN|-80.893784|80.893787349746532|340|1
35.478031|e81ced783437a4d013763ac3173f8a6a1af3f9a2|4.99|2014-12-04 17:16:00|80.8939826282094|1|3338365592|179|35.491662990721132|0|2|561|-80.86175|64|35.40953|FR PROD ORGANIC PRODUCE|0.0|4|ORG GRAPE TOMATOES|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00716310521844|FRESH PRODUCE|PRODUCE|-80.893784|80.893793458029279|209|1
35.478031|1f990a59cff05865ca56d21b3fd73645aaa67ce0|3.99|2015-03-02 11:24:00|80.8939826282094|1|3338324028|179|35.491662991994396|0|2|504|-80.8955|64|35.4437|FRESH BERRIES|2.0|4|BLACKBERRIES 5.6 OZ|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00033383240268|FRESH PRODUCE|PRODUCE|-80.893784|80.893790090795775|272|1
35.478031|d4c928279b98a99902a1696f819791f03575572b|13.98|2014-12-31 16:00:00|80.8939826282094|1|3338324000|179|35.491662991994396|0|2|504|-80.8955|64|35.4437|FRESH BERRIES|3.49|4|BLACKBERRIES 12 OZ|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00033383240015|FRESH PRODUCE|PRODUCE|-80.893784|80.893790090795775|272|2
35.478031|760125f8030297c53dd5309f0ac02b1f68b37fad|1.29|2014-10-10 10:35:00|80.8939826282094|1|7203670959|179|35.491662990721132|0|2|257|-80.86175|39|35.40953|TOMATOES|0.0|1|HTO TOMATO GREEN CHILIES.|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00072036709592|VEGETABLES-CAN/JAR|G1 GROCERY|-80.893784|80.893793458029279|209|1
35.478031|6869c711fb7da806363cb44e46f6a89c91425f5f|12.19|2015-02-16 16:38:00|80.8939826282094|1|1380023260|179|35.491662990721132|0|2|1280|-80.86175|48|35.40953|MULTI SERVE MEALS|0.0|5|STOUFF BAKED ZITI LRG FAMILY|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00013800197368|FROZEN MEALS|FROZEN|-80.893784|80.893793458029279|209|1
35.478031|7b71493d4cf195c73f54dea71173040f58645538|12.99|2014-10-16 18:58:00|80.8939826282094|1|1813831702|179|35.491662990721132|0|2|9961|-80.86175|887|35.40953|NFS-S/PREM-MERLOT|0.0|13|DYNAMITE MERLOT|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00018138317020|SUPER PREMIUM ($11-$14.99)|WINE|-80.893784|80.893793458029279|209|1
35.478031|d1bb744e97d953c7199a0471070a247d90a84aa7|6.49|2014-11-23 11:04:00|80.8939826282094|1|1708247047|179|35.491662991994396|0|2|215|-80.8955|31|35.4437|JERKY SNACKS|1.0|1|J LINK'S PREM CUT PRM RIB CUT|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00017082470478|SNACKS|G1 GROCERY|-80.893784|80.893790090795775|272|1
35.478031|aca9c15a49fa7eaafcdcdb0a43bee30e2d040623|1.29|2014-09-27 12:26:00|80.8939826282094|1|78616200387|179|35.491662990721132|0|2|31|-80.86175|4|35.40953|NON CARBONATED WATER|0.29|1|FRUITWATER BLACK RASPBERRY|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00786162003874|BOTTLED WATER|G1 GROCERY|-80.893784|80.893793458029279|209|1
35.478031|65923488074fd93e9b9011f12a33a6e5119abf92|2.99|2015-02-16 15:01:00|80.8939826282094|1|89899901000|179|35.491662990721132|0|2|31|-80.86175|4|35.40953|NON CARBONATED WATER|0.99|1|VITA COCO PURE COCONUT|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00898999010007|BOTTLED WATER|G1 GROCERY|-80.893784|80.893793458029279|209|1
35.478031|c72c367f510748477649cba72cc96169c32ae577|3.15|2015-01-25 17:15:00|80.8939826282094|1|2580002320|179|35.491662991994396|0|2|1278|-80.8955|48|35.4437|SINGLE SERVE NUTRITIONAL|0.65|5|WW SMART ONES MINI CHSEBURGERS|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00025800026715|FROZEN MEALS|FROZEN|-80.893784|80.893790090795775|272|1
35.478031|ecc79a483c931406de3b63f786b3085bdaf7d721|6.58|2014-12-06 12:04:00|80.8939826282094|1|2840018382|179|35.491662990721132|0|2|201|-80.86175|31|35.40953|POTATO CHIPS|0.0|1|BAKED TOSTITOS SCOOPS|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00028400184762|SNACKS|G1 GROCERY|-80.893784|80.893793458029279|209|2
35.478031|4d600120aa33680a7222d0fd5fd2142b3ec0e4b6|2.49|2014-09-23 18:31:00|80.8939826282094|1|7203688048|179|35.491662990721132|0|2|526|-80.86175|64|35.40953|FRESH MUSHROOMS|0.49|4|HT SLICED BABY BELLAS|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00072036880482|FRESH PRODUCE|PRODUCE|-80.893784|80.893793458029279|209|1
35.478031|23863f52ec27b2ff54d89b2f697070d0db362156|2.99|2015-02-04 15:25:00|80.8939826282094|1|3338365583|179|35.491662991994396|0|2|522|-80.8955|64|35.4437|FRESH TOMATOES|1.5|4|SWEET GRAPE TOMATO (PINT)|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00072036880284|FRESH PRODUCE|PRODUCE|-80.893784|80.893790090795775|272|1
35.478031|73f4fa44243098a99b41baba3c9dc469b05c6e39|25.74|2014-12-13 12:42:00|80.8939826282094|1|7535307312|179|35.491662990721132|0|2|6253|-80.86175|1550|35.40953|TAPES/DUCT TAPE|0.0|18|CARTON TAPE 48MMX50M CLEAR|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00075353073124|HARDWARE|GM|-80.893784|80.893793458029279|209|6
35.478031|e3a1e429fd93a8d843b493092b95b6e43d5e747e|18.99|2014-12-24 11:41:00|80.8939826282094|1|89105600087|179|35.491662990721132|0|2|62|-80.86175|7|35.40953|SPECIALTY BAR/BOX CHOCOLATE|2.0|1|I/OFUNKY CHUNKY CHOC CARM PCRN|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00891056000874|CANDY|G1 GROCERY|-80.893784|80.893793458029279|209|1
35.478031|90be96a85d29c7dda8b23a09d5d636d235119723|2.89|2015-01-04 10:52:00|80.8939826282094|1|1200037401|179|35.491662990721132|0|2|854|-80.86175|32|35.40953|LIQUID ICED COFFEES|0.0|1|STARBUCKS REFRESH STRW LEMONAD|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00012000374012|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.893784|80.893793458029279|209|1
35.478031|5eb5a11b80c6d8ab8e7127a22fde44fd713c9675|4.29|2014-11-13 10:07:00|80.8939826282094|1|2840015636|179|35.491662992623695|0|2|204|-80.861571|31|35.444615|TORTILLA CHIPS|1.79|1|DORTIOS NACHO CHEESE|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00028400156363|SNACKS|G1 GROCERY|-80.893784|80.893787349746532|340|1
35.478031|4f38074fc9602377727a2bd9ba0c0003b72eb7ca|7.99|2015-02-01 15:11:00|80.8939826282094|1|2100061161|179|35.491662992623695|0|2|314|-80.861571|52|35.444615|CHEESE-PROCESSED-OTHER|1.0|3|KRAFT VELVEETA CHEESE|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00021000611614|CHEESE|DAIRY|-80.893784|80.893787349746532|340|1
35.478031|d34e58157289245df1fff8e4f7aa6894044840c2|5.99|2014-12-23 20:46:00|80.8939826282094|1|7041101343|179|35.491662991994396|0|2|215|-80.8955|31|35.4437|JERKY SNACKS|1.0|1|OBERTO NTRL BACON JERKY|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00070411603725|SNACKS|G1 GROCERY|-80.893784|80.893790090795775|272|1
35.478031|84f9a38a833b79a583c17b9fb356998b8b66f4ec|11.98|2014-11-16 12:53:00|80.8939826282094|1|7041101343|179|35.491662990721132|0|2|215|-80.86175|31|35.40953|JERKY SNACKS|3.0|1|OBERTO NTRL BEEF JRKY-TERIYAKI|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00070411013432|SNACKS|G1 GROCERY|-80.893784|80.893793458029279|209|2
35.478031|ddd0a1e5b16dbb3b55b1f40447862ce9e4d446af|2.99|2015-02-21 18:29:00|80.8939826282094|1|4000023132|179|35.491662990721132|0|2|727|-80.86175|7|35.40953|SEASONAL CANDY-SINGLE FAC|0.49|1|I/O(E15)STARBRST FAVRED JLY BN|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00040000231325|CANDY|G1 GROCERY|-80.893784|80.893793458029279|209|1
35.478031|787be40b027439809ee76edb5a031e66fff3f4f2|5.98|2015-02-02 15:14:00|80.8939826282094|1|3700000309|179|35.491662990721132|0|2|4070|-80.86175|1080|35.40953|TOOTHPASTE-BAKING SODA|0.98|17|CREST BAKING SODA& PER-32024|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00037000320241|ORAL HYGIENE|HBC|-80.893784|80.893793458029279|209|2
35.478031|f395db0d09fa7239462c02f66d5f012a4b49d7b9|6.58|2015-02-14 12:04:00|80.8939826282094|1|84667500117|179|35.491662991994396|0|2|1260|-80.8955|1|35.4437|TODDLER HAND HELD|1.64|1|PLUM TEENSY FRUITS BERRY|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00846675001177|BABY FOOD|G1 GROCERY|-80.893784|80.893790090795775|272|2
35.478031|d89bf855ea9c0a6066d2a7e7636c52d377010831|4.29|2015-01-09 09:38:00|80.8939826282094|1|7341000305|179|35.491662992623695|0|2|1026|-80.861571|162|35.444615|WHEAT|2.14|7|ARN CNTRY OATMEAL BREAD WP PP|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00073410003558|SLICED BREAD|COMMERCIAL BAKERY|-80.893784|80.893787349746532|340|1
35.478031|acf1b4a65ac31861c5a78295b1347f0e0c5d8193|3.99|2014-11-21 18:46:00|80.8939826282094|1|2392320200|179|35.491662990721132|0|2|1260|-80.86175|1|35.40953|TODDLER HAND HELD|0.0|1|E B SESAME STREET HNY STK CRNC|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00023923203013|BABY FOOD|G1 GROCERY|-80.893784|80.893793458029279|209|1
35.478031|9b6c5331159c97bce47533f665fe4ebd515a067b|2.35|2014-12-02 11:55:00|80.8939826282094|1|1500004873|179|35.491662990721132|0|2|1259|-80.86175|1|35.40953|TODDLER MEALS|0.0|1|GERB LIL ENT MACARONI CHEESE|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00015000048730|BABY FOOD|G1 GROCERY|-80.893784|80.893793458029279|209|1
35.478031|05c3080ca1b49b797b344bf7f089694b052366bc|1.69|2014-12-27 11:36:00|80.8939826282094|1|1708200003|179|35.491662991994396|0|2|206|-80.8955|31|35.4437|FRONT END SNACKS|0.2|1|J LINKS ORIGINAL BEEF STEAKS|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00017082000033|SNACKS|G1 GROCERY|-80.893784|80.893790090795775|272|1
35.478031|87a2e3430fe294137348404e812c93602c30d8d3|2.19|2015-01-01 11:26:00|80.8939826282094|1|38137008256|179|35.491662991994396|0|2|4834|-80.8955|1235|35.4437|COTTON/SWABS|0.0|17|JOHNSONS SAFETY SWABS-08256|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00381370082569|FIRST AID|HBC|-80.893784|80.893790090795775|272|1
35.478031|b845490797c90cc8c5f921201fb618f73c8a0d42|4.89|2015-01-01 17:48:00|80.8939826282094|1|74236526435|179|35.491662992623695|0|2|345|-80.861571|57|35.444615|ORGANIC MILK|0.0|3|HORIZON REDUCE FAT DHA|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00742365264351|MILK|DAIRY|-80.893784|80.893787349746532|340|1
35.478031|683205074a4f5755b93598e4653c69c6149fde67|4.49|2015-03-07 17:49:00|80.8939826282094|1|74236526405|179|35.491662991994396|0|2|345|-80.8955|57|35.4437|ORGANIC MILK|0.0|3|HORIZON ORGANIC WHOLE MILK|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00742365264450|MILK|DAIRY|-80.893784|80.893790090795775|272|1
35.478031|f251d672009f42d9227c7c93a56f7f1a7eb0dd04|2.39|2014-10-09 18:11:00|80.8939826282094|1|600980280204|179|35.491662990721132|0|2|30|-80.86175|4|35.40953|CARBONATED WATER|0.0|1|TRU COCO COCONUT WATR&MANGO JC|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|06009802802045|BOTTLED WATER|G1 GROCERY|-80.893784|80.893793458029279|209|1
35.478031|0c5baf97bff11b1ecd0e59dfa390c2a0f95ed198|11.99|2014-09-13 18:33:00|80.8939826282094|1|80489001212|179|35.491662990721132|0|2|194|-80.86175|30|35.40953|OLIVE OIL|3.0|1|SAN LEANDRO ORGANIC OIL|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00804890012125|SHORTENING/OIL|G1 GROCERY|-80.893784|80.893793458029279|209|1
35.478031|499d95f6fb87ced5f76d2169358edde5a27914b2|8.78|2014-12-21 15:50:00|80.8939826282094|1|5100020921|179|35.491662990721132|0|2|173|-80.86175|27|35.40953|CANNED POULTRY|1.78|1|SWANSON GRILLED CHUNK CHICKEN|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00051000209221|PREPARED FOODS-RTS|G1 GROCERY|-80.893784|80.893793458029279|209|2
35.478031|c5e21a7b1823a6e9467c2ec57b5d9d9fb7050348|5.79|2015-01-29 13:09:00|80.8939826282094|1|7007480240|179|35.491662991994396|0|2|3|-80.8955|1|35.4437|FORMULA RTF|0.8|1|PEDIALYTE GRAPE FLAVOR|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00070074802404|BABY FOOD|G1 GROCERY|-80.893784|80.893790090795775|272|1
35.478031|15764c2ba71e4d40a009beaebb87c9d8f9cab3ec|3.99|2015-01-17 13:12:00|80.8939826282094|1|85281048912|179|35.491662991994396|0|2|364|-80.8955|55|35.4437|ORGANIC AND CF EGGS|0.0|3|LOL CAGE FREE A LRG BRWN EGGS|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00852810489120|EGGS FRESH|DAIRY|-80.893784|80.893790090795775|272|1
35.478031|6d12d184b0c14d71fab1847a77adafabce9be913|15.99|2014-09-18 18:52:00|80.8939826282094|1|7023666063|179|35.491662990721132|0|2|751|-80.86175|87|35.40953|NFS-BOUQUETS|0.0|9|$15.99 BOUQUET|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00070236660637|FLORAL|FLORAL|-80.893784|80.893793458029279|209|1
35.478031|733fee425533c9f106a4ddb4a1093a029f9ee7e1|16.99|2014-11-08 14:50:00|80.8939826282094|1|1951839226|179|35.491662991994396|0|2|742|-80.8955|87|35.4437|"NFS-BLOOMING 4"""|0.0|9|"5"" ORCHID IN BIO POT"|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00019518392262|FLORAL|FLORAL|-80.893784|80.893790090795775|272|1
35.478031|a6f72edb618307591a5c36d17e8b7bb6e2abbf7d|5.29|2014-11-12 10:08:00|80.8939826282094|1|3680034644|179|35.491662992623695|0|2|4338|-80.861571|1205|35.444615|PAIN RELIEVER-CHILDREN|0.0|17|TC INFANT PAIN RLF DROPS GRAPE|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00036800346444|PAIN RELIEF|HBC|-80.893784|80.893787349746532|340|1
35.478031|894d1ffb5dfdf03cb836880b6bae82d5f185dc07|4.89|2014-11-08 17:11:00|80.8939826282094|1|74236526435|179|35.491662990721132|0|2|345|-80.86175|57|35.40953|ORGANIC MILK|0.0|3|HORIZON WHOLE  DHA|60333193007241337434451bcf0f7f7e0539edde|0.9419377890696846|35.490689277687849|00742365264474|MILK|DAIRY|-80.893784|80.893793458029279|209|1
35.061685|4e37b208dcb685ca9f0207224004c7e2cf8e88ca|9.29|2014-11-20 15:11:00|1.4132775322775095|2|76211188813|475|0.611941844547108|0|58|37|-80.994596|10|35.061685|PODS/CUPS/SINGLES|2.3|1|STARBUCKS HOUSE BLEND KCUP|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00762111888136|COFFEE|G1 GROCERY|-80.994596|1.4136223765226292|475|1
35.061685|d7b320b91946ae8161e9c10df91858dd41f0840e|2.79|2014-09-12 13:36:00|1.4132775322775095|2|7203688211|475|0.611941844547108|0|58|555|-80.994596|64|35.061685|PACKAGED SALADS|0.0|4|HT PREMIUM ROMAINE|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00072036882110|FRESH PRODUCE|PRODUCE|-80.994596|1.4136223765226292|475|1
35.061685|ff460adabd9edd58dfaea2734f8d8c536ea779df|7.38|2015-01-13 17:21:00|1.4132775322775095|2||475|0.611941844547108|0|58|503|-80.994596|64|35.061685|FRESH GRAPES|0.0|4|GREEN GRAPES, SEEDLESS 12/16|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00204022000004|FRESH PRODUCE|PRODUCE|-80.994596|1.4136223765226292|475|1
35.061685|dc86262d9bc3e283252cf2e1401b61e2129a5929|3.99|2015-01-05 16:13:00|1.4132775322775095|2|75166677005|475|0.611941844547108|0|58|522|-80.994596|64|35.061685|FRESH TOMATOES|0.0|4|NATURESWEET CHERUBS 10.5 OZ|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00751666770058|FRESH PRODUCE|PRODUCE|-80.994596|1.4136223765226292|475|1
35.061685|8ed5bc1f12a8cb2e6cceaee1ea278497e0c6e432|3.99|2014-10-13 17:15:00|1.4132775322775095|2|75166677005|475|0.611941844547108|0|58|522|-80.994596|64|35.061685|FRESH TOMATOES|0.0|4|NATURESWEET CHERUBS 10.5 OZ|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00751666770058|FRESH PRODUCE|PRODUCE|-80.994596|1.4136223765226292|475|1
35.061685|2d3801283bafb042c48fb695718011f16f6a25b6|3.99|2014-12-21 16:22:00|1.4132775322775095|2|75166677005|475|0.611941844547108|0|58|522|-80.994596|64|35.061685|FRESH TOMATOES|0.0|4|NATURESWEET CHERUBS 10.5 OZ|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00751666770058|FRESH PRODUCE|PRODUCE|-80.994596|1.4136223765226292|475|1
35.061685|8b344a31a1c4bff2009d2d006f04e61972a73bda|3.99|2015-03-03 17:27:00|1.4132775322775095|2|75166677005|475|0.611941844547108|0|58|522|-80.994596|64|35.061685|FRESH TOMATOES|0.0|4|NATURESWEET CHERUBS 10.5 OZ|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00751666770058|FRESH PRODUCE|PRODUCE|-80.994596|1.4136223765226292|475|1
35.061685|f3595b8475d15b9ac0ba6425d0da51bce871609f|3.99|2014-12-02 19:55:00|1.4132775322775095|2|75166677005|475|0.611941844547108|0|58|522|-80.994596|64|35.061685|FRESH TOMATOES|0.0|4|NATURESWEET CHERUBS 10.5 OZ|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00751666770058|FRESH PRODUCE|PRODUCE|-80.994596|1.4136223765226292|475|1
35.061685|781f963ff0ee3e0403960914f79a3f9484ef1299|2.69|2015-02-11 15:38:00|80.994598860450068|2|7680851558|475|35.08002036854041|0|53|149|-80.97058|23|35.03469|WHSE PASTA CORE|0.0|1|BARILLA PASTA LASAGNE|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|35.072594466811061|00895059000619|PASTA|G1 GROCERY|-80.994596|80.994599868442151|82|1
35.061685|5aa685427a95fdb49c1284c903ec2e2440696645|5.19|2015-02-08 19:28:00|1.4132775322775095|2|74236526435|475|0.611941844547108|0|58|345|-80.994596|57|35.061685|ORGANIC MILK|0.0|3|HORIZON ORGANIC FF DHA|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00742365003295|MILK|DAIRY|-80.994596|1.4136223765226292|475|1
35.061685|1fdf4cf8917e197e92b847479d19b3319bec19cc|4.89|2014-11-05 19:28:00|1.4132775322775095|2|74236526435|475|0.611941844547108|0|58|345|-80.994596|57|35.061685|ORGANIC MILK|0.0|3|HORIZON ORGANIC FF DHA|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00742365003295|MILK|DAIRY|-80.994596|1.4136223765226292|475|1
35.061685|e852f15a2a9547586f2f8a744d0a13b5bfd0cd54|4.89|2015-01-12 12:26:00|1.4132775322775095|2|74236526435|475|0.611941844547108|0|58|345|-80.994596|57|35.061685|ORGANIC MILK|0.0|3|HORIZON ORGANIC FF DHA|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00742365003295|MILK|DAIRY|-80.994596|1.4136223765226292|475|1
35.061685|0ab93d14c420f9e03350d27543d1043739504099|7.96|2014-11-13 15:42:00|80.994598860450068|2|7365121405|475|35.08002036854041|0|53|160|-80.97058|25|35.03469|OLIVES|0.99|1|MARIO OLIVE RIPE SLICED 2.25|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|35.072594466811061|00073651214058|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.994596|80.994599868442151|82|4
35.061685|57082f754d329cd5942133c4e592edea0e7609a9|7.27|2014-12-14 08:28:00|1.4132775322775095|2|20037600000|475|0.611941844547108|0|58|1801|-80.994596|400|35.061685|FFM TURKEY|0.0|6|TURKEY BREAST|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00200376000004|FFM MEAT|DELI|-80.994596|1.4136223765226292|475|1
35.061685|ba42ce5b9846ffc3b4db435b215efacba1c9a12f|0.99|2015-01-21 17:15:00|1.4132775322775095|2|5210009860|475|0.611941844547108|0|58|75|-80.994596|34|35.061685|GRAVY MIXES|0.0|1|MC CORMICK GF BROWN GRAVY|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00052100026923|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.994596|1.4136223765226292|475|1
35.061685|3fc1493b858f28d76cba495ad118b1fee4f4de77|4.99|2015-02-22 09:52:00|1.4132775322775095|2|7104000015|475|0.611941844547108|0|58|332|-80.994596|52|35.061685|STRING/SNACK|0.0|3|POLLY-O STRING CHEESE 2%|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00071040000602|CHEESE|DAIRY|-80.994596|1.4136223765226292|475|1
35.061685|14f7f96824892d53634f104421532cdcc287e3ce|4.99|2015-02-15 08:44:00|1.4132775322775095|2|7104000015|475|0.611941844547108|0|58|332|-80.994596|52|35.061685|STRING/SNACK|0.0|3|POLLY-O STRING CHEESE 2%|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00071040000602|CHEESE|DAIRY|-80.994596|1.4136223765226292|475|1
35.061685|cd44bd14f80608dd5374f70114400524772c58e5|2.99|2014-09-15 12:23:00|1.4132775322775095|2|1228951006|475|0.611941844547108|0|58|523|-80.994596|64|35.061685|FRESH POTATOES|0.0|4|SS STEAMABL RED POTATO 24OZ|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00012289510064|FRESH PRODUCE|PRODUCE|-80.994596|1.4136223765226292|475|1
35.061685|a8fccfe93ad94ed9ff3752364068a94e7de255c5|4.49|2014-11-10 16:45:00|1.4132775322775095|2|76770700167|475|0.611941844547108|0|58|312|-80.994596|51|35.061685|BUTTER|1.12|3|KERRYGOLD SPREADABLE BUTTER|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00767707001678|BUTTER & MARGARINE|DAIRY|-80.994596|1.4136223765226292|475|1
35.061685|277757b28b219c428939e82cf2d45e1719815fef|4.49|2014-12-06 19:46:00|1.4132775322775095|2|74236526405|475|0.611941844547108|0|58|345|-80.994596|57|35.061685|ORGANIC MILK|0.0|3|HORIZON ORGANIC FF MILK|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00742365264054|MILK|DAIRY|-80.994596|1.4136223765226292|475|1
35.061685|ed83638f7a037563909eb698a3e1c8613e16d3e8|4.49|2015-02-01 18:41:00|80.994598860450068|2|74236526405|475|35.08002036854041|0|53|345|-80.97058|57|35.03469|ORGANIC MILK|0.0|3|HORIZON ORGANIC FF MILK|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|35.072594466811061|00742365264054|MILK|DAIRY|-80.994596|80.994599868442151|82|1
35.061685|9d8b0d17e018d8912c52f97daee57bd5e1902a72|7.78|2015-02-25 14:59:00|80.994598860450068|2|4610000084|475|35.080020365608341|0|53|318|-80.837892|52|34.937113|SHREDDED/GRATED CHEESE|1.95|3|SARGENTO REDUCED FAT MOZZ|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|35.072594466811061|00046100000823|CHEESE|DAIRY|-80.994596|80.994609246917534|372|2
35.061685|f5eba5ea6c4a5803779f3369735f484ee0e8099b|3.95|2014-10-06 17:00:00|1.4132775322775095|2|4610000084|475|0.611941844547108|0|58|318|-80.994596|52|35.061685|SHREDDED/GRATED CHEESE|1.98|3|SARGENTO REDUCED FAT MOZZ|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00046100000823|CHEESE|DAIRY|-80.994596|1.4136223765226292|475|1
35.061685|af73890ee4bd4e44146029324e2779aaacd297f7|9.9|2014-09-28 08:30:00|1.4132775322775095|2|1780014597|475|0.611941844547108|0|58|154|-80.994596|24|35.061685|NFS-CAT FOOD WET|1.4000000000000004|1|ONE BRAISED CUTS CHICKN GRAVY|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00017800146029|PET FOOD/SUPPLIES|G1 GROCERY|-80.994596|1.4136223765226292|475|10
35.061685|b7a93670c951a305802de6a181d801ca8c6b99fe|5.39|2014-11-25 17:34:00|1.4132775322775095|2|7203000018|475|0.611941844547108|0|58|1685|-80.994596|385|35.061685|ENTENMANNS (SWEET GOODS)|2.7|14|ENT RICH FROSTED DONUTS PP|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00072030000183|SWEET GOODS|BAKERY|-80.994596|1.4136223765226292|475|1
35.061685|b3e13525b66818d67d48be5fb49cad3206633afd|2.25|2014-12-31 14:02:00|1.4132775322775095|2||475|0.611941844547108|0|58|1617|-80.994596|373|35.061685|ROLLS BULK|0.0|14|BULK ROLLS|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00072036955555|ROLLS|BAKERY|-80.994596|1.4136223765226292|475|3
35.061685|80c823b754002fa4e3ef768c137ff0aeda2fac40|1.49|2014-09-29 12:04:00|1.4132775322775095|2|2840002819|475|0.611941844547108|0|58|206|-80.994596|31|35.061685|FRONT END SNACKS|0.0|1|LAYS CLASSIC|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00028400027960|SNACKS|G1 GROCERY|-80.994596|1.4136223765226292|475|1
35.061685|0cdcaf2aa777db2624097f1a44c758f2b5a63689|6.98|2014-10-19 11:03:00|1.4132775322775095|2|2800000820|475|0.611941844547108|0|58|131|-80.994596|20|35.061685|GRAPE JUICE-SHELF|0.4|1|JUICY JUICE WHT GRAPE|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00028000108366|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.994596|1.4136223765226292|475|2
35.061685|e879307a60ef280826d79cf66252dcbbbe84f911|3.49|2015-01-10 11:05:00|1.4132775322775095|2|2840023981|475|0.611941844547108|0|58|203|-80.994596|31|35.061685|CHEESE SNACKS|0.0|1|CHEETOS CHEDDAR JALAPENO|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00028400239837|SNACKS|G1 GROCERY|-80.994596|1.4136223765226292|475|1
35.061685|f04786c7ced81590301e4e1f42961256ae36c2d6|15.99|2014-10-20 17:31:00|1.4132775322775095|2|87126000465|475|0.611941844547108|0|58|740|-80.994596|87|35.061685|NFS-ROSE BQT|0.0|9|DZ ROSE BQT 3 RED/5 COLOR  ELI|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00871260004653|FLORAL|FLORAL|-80.994596|1.4136223765226292|475|1
35.061685|55a40c6b4711c25accc0eebdbbce283d62b677ec|1.95|2015-02-25 15:01:00|80.994598860450068|2|76211103726|475|35.080020365608341|0|53|1599|-80.837892|370|34.937113|PASTRY|0.0|22|"SBUX ""LB"" MADELINES"|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|35.072594466811061|00762111037268|STARBUCKS|COFFEE SHOP|-80.994596|80.994609246917534|372|1
35.061685|820bc794e6dea31a814659fab95c9fe4c3f5cb44|6.79|2014-12-02 13:48:00|1.4132775322775095|2|1200080994|475|0.611941844547108|0|58|55|-80.994596|8|35.061685|REGULAR|1.8|23|MUG ROOT BEER FRIDGEMATE|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00012000810008|CARBONATED BEVERAGES|BEVERAGE|-80.994596|1.4136223765226292|475|1
35.061685|4c8785a4c5c1594d15b9b5d822958ce85b1604f4|5.98|2014-12-10 10:07:00|1.4132775322775095|2|1410009840|475|0.611941844547108|0|58|1256|-80.994596|13|35.061685|WHOLESOME CRACKERS|1.98|1|PP PF BAKED NATURALS 4 CHEESE|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00014100092308|CRACKERS|G1 GROCERY|-80.994596|1.4136223765226292|475|2
35.061685|14cc52bdf966c92fac069ac4478fc490a254c4ee|3.39|2014-11-12 20:07:00|1.4132775322775095|2|5000012734|475|0.611941844547108|0|58|341|-80.994596|57|35.061685|CREAMERS|0.89|3|COFFEEMATE SF FRENCH VANILLA|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00050000848119|MILK|DAIRY|-80.994596|1.4136223765226292|475|1
35.061685|eabff9b8d80ddf5756f5a6f80fc87e7602fbfa4a|6.49|2015-02-23 16:25:00|1.4132775322775095|2|4470006376|475|0.611941844547108|0|58|485|-80.994596|101|35.061685|PREMIUM WIENERS|3.25|19|OM SELECTS ANGUS BEEF FRANK|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00044700063774|WIENERS|CASE READY MEATS|-80.994596|1.4136223765226292|475|1
35.061685|73e0ec7fcea547f92b525426f20703ee49c0d664|3.59|2015-02-25 11:08:00|1.4132775322775095|2|1070051851|475|0.611941844547108|0|58|52|-80.994596|7|35.061685|PKG NON CHOC|0.0|1|JOLLY RANCHER ASTD ORIGINAL|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00010700518514|CANDY|G1 GROCERY|-80.994596|1.4136223765226292|475|1
35.061685|9db343218c75e8977cabb288ddf47509dd533e5b|3.59|2014-12-30 07:03:00|1.4132775322775095|2|1070051851|475|0.611941844547108|0|58|52|-80.994596|7|35.061685|PKG NON CHOC|0.0|1|JOLLY RANCHER ASTD ORIGINAL|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00010700518514|CANDY|G1 GROCERY|-80.994596|1.4136223765226292|475|1
35.061685|95fbe3bc5e9eea631f156d828bc251bccf21f405|3.59|2014-12-15 16:15:00|1.4132775322775095|2|1070051851|475|0.611941844547108|0|58|52|-80.994596|7|35.061685|PKG NON CHOC|0.0|1|JOLLY RANCHER ASTD ORIGINAL|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00010700518514|CANDY|G1 GROCERY|-80.994596|1.4136223765226292|475|1
35.061685|493fe3b2f233681610cc9b3671a994f32a6812fa|3.59|2015-01-05 10:26:00|1.4132775322775095|2|1070051851|475|0.611941844547108|0|58|52|-80.994596|7|35.061685|PKG NON CHOC|0.0|1|JOLLY RANCHER ASTD ORIGINAL|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00010700518514|CANDY|G1 GROCERY|-80.994596|1.4136223765226292|475|1
35.061685|d02dd13b2a7f5c0bc40a3563b318db8533a457b2|3.59|2014-11-28 13:41:00|1.4132775322775095|2|1070051851|475|0.611941844547108|0|58|52|-80.994596|7|35.061685|PKG NON CHOC|0.0|1|JOLLY RANCHER ASTD ORIGINAL|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00010700518514|CANDY|G1 GROCERY|-80.994596|1.4136223765226292|475|1
35.061685|aee3dd31e6b5e30c94ab15be3ed1962355825663|6.99|2014-11-07 17:23:00|1.4132775322775095|2|4400088032|475|0.611941844547108|0|58|1252|-80.994596|12|35.061685|LUNCH BOX COOKIES|1.0|1|NABISCO SS CHIPS AHOY MINI|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00044000020279|COOKIES|G1 GROCERY|-80.994596|1.4136223765226292|475|1
35.061685|72caabc01c8cd0e28910e98697e44ccabd00884f|6.98|2015-02-28 11:36:00|1.4132775322775095|2|7797503405|475|0.611941844547108|0|58|202|-80.994596|31|35.061685|PRETZELS|0.98|1|SNYDERS BUTTER SNAPS|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00077975034057|SNACKS|G1 GROCERY|-80.994596|1.4136223765226292|475|2
35.061685|28612b5066d31a2b6464c2e8d68c5f75f58fb724|6.98|2014-11-10 11:19:00|1.4132775322775095|2|7797503405|475|0.611941844547108|0|58|202|-80.994596|31|35.061685|PRETZELS|0.98|1|SNYDERS BUTTER SNAPS|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00077975034057|SNACKS|G1 GROCERY|-80.994596|1.4136223765226292|475|2
35.061685|4a3cc8d498066696364c20a98ab4398e3f028d6e|6.49|2015-01-06 16:07:00|1.4132775322775095|2|4242116019|475|0.611941844547108|0|58|1855|-80.994596|430|35.061685|BH SALAMI/CHUBBS|0.0|6|BH ANTI GENOA & PROVOLONE|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00042421160192|SPECIALTY MEAT|DELI|-80.994596|1.4136223765226292|475|1
35.061685|3df5088dd24275a0471c7e4dc67ca20e9b4a2e0b|0.29|2015-02-27 13:54:00|1.4132775322775095|2|4133507899|475|0.611941844547108|0|58|1984|-80.994596|480|35.061685|PC CONDIMENTS|0.0|6|KEN'S CAESAR DRESSING|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00041335082798|DRY GOODS|DELI|-80.994596|1.4136223765226292|475|1
35.061685|778f635ff36ebab66fa3f3fb0842318b8d92099f|1.19|2015-01-23 11:19:00|1.4132775322775095|2|7550000001|475|0.611941844547108|0|58|76|-80.994596|11|35.061685|MEAT SAUCES|0.0|1|TEXAS PETE HOT SAUCE 6|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00075500000010|CONDIMENTS|G1 GROCERY|-80.994596|1.4136223765226292|475|1
35.061685|f44ae374118e677704c274dd1608ecb399e45337|7.38|2015-01-12 15:41:00|80.994598860450068|2|5000030262|475|35.08002036854041|0|53|341|-80.97058|57|35.03469|CREAMERS|0.0|3|COFFEE MATE FAT FREE|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|35.072594466811061|00050000339525|MILK|DAIRY|-80.994596|80.994599868442151|82|2
35.061685|6ce7bc4fd097c17b5a2257eb1022b4b143db6979|2.91|2015-01-11 08:57:00|1.4132775322775095|2|7203698757|475|0.611941844547108|0|58|31|-80.994596|4|35.061685|NON CARBONATED WATER|0.0|1|HT DISTILLED WATER|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00072036360601|BOTTLED WATER|G1 GROCERY|-80.994596|1.4136223765226292|475|3
35.061685|a4ae5b630890af4f5d5dd2be2b1d2ef7e3220db1|9.38|2014-11-08 16:09:00|1.4132775322775095|2|20496000000|475|0.611941844547108|0|58|755|-80.994596|87|35.061685|NFS-BALLOONS|0.0|9|*BALLOONS|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00204960000005|FLORAL|FLORAL|-80.994596|1.4136223765226292|475|1
35.061685|dab97c5981a0fda1170d65c8b504fe5ba352e5dc|0.29|2015-02-24 13:42:00|1.4132775322775095|2|4133507899|475|0.611941844547108|0|58|1984|-80.994596|480|35.061685|PC CONDIMENTS|0.0|6|KEN'S LITE ITLIAN DRESSING|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00041335080190|DRY GOODS|DELI|-80.994596|1.4136223765226292|475|1
35.061685|2d1431caabf3675f031331aa974cd33019f4f6ec|0.29|2014-10-01 11:36:00|1.4132775322775095|2|4133507899|475|0.611941844547108|0|58|1984|-80.994596|480|35.061685|PC CONDIMENTS|0.0|6|KEN'S LITE ITLIAN DRESSING|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00041335080190|DRY GOODS|DELI|-80.994596|1.4136223765226292|475|1
35.061685|789e3f07618d122b531094f0f593b20e573cae1a|1.99|2015-02-13 18:00:00|1.4132775322775095|2||475|0.611941844547108|0|58|500|-80.994596|64|35.061685|FRESH APPLES|0.34|4|GOLD DEL APPLE EASTERN|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00204137000005|FRESH PRODUCE|PRODUCE|-80.994596|1.4136223765226292|475|1
35.061685|deefc0ec56a84b0ccf032a8cb1e2be242c5877f9|2.49|2014-12-01 14:41:00|1.4132775322775095|2|7279900861|475|0.611941844547108|0|58|50|-80.994596|7|35.061685|PEG CANDY|0.0|1|WERTHER'S ORIGINAL BUTTER TOFF|649a44bdab4cdb88c58d289550f53961a3249fef|1.2669297067003125|0.61177642288969325|00072799008611|CANDY|G1 GROCERY|-80.994596|1.4136223765226292|475|1
35.323246|43b8ba794672c509c28ee5a2f18e43f8138aa947|16.53|2015-02-16 16:41:00|1.4102725052409182|4|20188000000|166|0.6165069451919168|0|1|299|-80.945176|49|35.323246|ANGUS BEEF|0.0|2|ANGUS BEEF BNLS CHUCK ROAST|671ceca91db15d80a0c0e5acc89274eeefcbf927|0.8246694273071761|0.61833652052202714|00201880000009|BEEF|MEAT|-80.945176|1.4127598348062935|166|1
35.323246|812fb5de9fe7cc108dc866bd92eaf4728a5b55ef|17.39|2014-12-06 18:13:00|1.4102725052409182|4|27085500000|166|0.6165069451919168|0|1|973|-80.945176|201|35.323246|FRESH PERDUE CHICKEN|0.0|2|PERDUE OVEN STUFFER ROASTER|671ceca91db15d80a0c0e5acc89274eeefcbf927|0.8246694273071761|0.61833652052202714|00270855000009|POULTRY|MEAT|-80.945176|1.4127598348062935|166|1
35.323246|895a640a2482d283e610621cf3988a462b6db018|19.36|2014-12-06 18:15:00|1.4102725052409182|4|27085500000|166|0.6165069451919168|0|1|973|-80.945176|201|35.323246|FRESH PERDUE CHICKEN|0.0|2|PERDUE OVEN STUFFER ROASTER|671ceca91db15d80a0c0e5acc89274eeefcbf927|0.8246694273071761|0.61833652052202714|00270855000009|POULTRY|MEAT|-80.945176|1.4127598348062935|166|1
35.323246|5ea463b6c5b33397b9a6c2e434c6ed9772117d26|7.69|2015-01-16 15:42:00|1.4102725052409182|4|8087817730|166|0.6165069451919168|0|1|3503|-80.945176|1045|35.323246|CONDITIONER-PREMIUM|1.69|17|PANTENE COND DAM DETOX REBUILD|671ceca91db15d80a0c0e5acc89274eeefcbf927|0.8246694273071761|0.61833652052202714|00080878177301|HAIR & SCALP CARE|HBC|-80.945176|1.4127598348062935|166|1
35.323246|f2c021a7d4d84281f843c87da0363e4c1298e74c|5.98|2014-12-22 17:23:00|1.4102725052409182|4|4470036113|166|0.6165069451919168|0|1|659|-80.945176|103|35.323246|CHILDRENS LUNCH SNACKS|0.2|19|FUNPACK LUNCH TRKY/AMER STACK|671ceca91db15d80a0c0e5acc89274eeefcbf927|0.8246694273071761|0.61833652052202714|00044700006740|LUNCH SNACKS|CASE READY MEATS|-80.945176|1.4127598348062935|166|2
35.323246|5460960445e052c4ceb8f697d2d94dc393617259|1.19|2015-01-17 17:56:00|1.4102725052409182|4|1500007135|166|0.6165069451919168|0|1|6|-80.945176|1|35.323246|JARRED BABY FOOD|0.19|1|GERBER 1ST SWEET POTATOES|671ceca91db15d80a0c0e5acc89274eeefcbf927|0.8246694273071761|0.61833652052202714|00015000071189|BABY FOOD|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|860992e6d847d719bcaadbc86efa2baed9b083b3|35.88|2014-12-13 16:46:00|1.4102725052409182|4|20496100000|166|0.6165069451919168|0|1|754|-80.945176|87|35.323246|NFS-SGLE STEM CUT FLOWER|0.0|9|*SINGLE STEM CUT FLOWERS|671ceca91db15d80a0c0e5acc89274eeefcbf927|0.8246694273071761|0.61833652052202714|00204961000004|FLORAL|FLORAL|-80.945176|1.4127598348062935|166|2
35.323246|6bb5adc3ba6742b63cde43edfc720b33e1d5a544|28.99|2015-01-11 17:54:00|1.4102725052409182|4|5000011178|166|0.6165069451919168|0|1|1181|-80.945176|1|35.323246|BABY FORMULA - DRY|3.0|1|L GERBER GOODSTART GENTLE PWDR|671ceca91db15d80a0c0e5acc89274eeefcbf927|0.8246694273071761|0.61833652052202714|00050000111787|BABY FOOD|G1 GROCERY|-80.945176|1.4127598348062935|166|1
34.977331|267582f6720af6506193869fc1d6eb97292b3344|3.29|2014-12-19 16:29:00|1.41290891556208|3|2840004768|149|0.6104695895098807|0|33|202|-81.027334|31|34.977331|PRETZELS|0.29|1|ROLD GOLD PRETZEL CLASSIC THIN|67e73b6075b00299fbe43b733da4006ae51c2ec2|6.232193769327634|0.61055446569467375|00028400047678|SNACKS|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|aa75ddbaae7a36bb2ad9e00757d51ea927777195|6.58|2014-12-13 11:50:00|1.41290891556208|3|2840004768|149|0.6104695895098807|0|33|202|-81.027334|31|34.977331|PRETZELS|1.58|1|ROLD GOLD PRETZEL CLASSIC THIN|67e73b6075b00299fbe43b733da4006ae51c2ec2|6.232193769327634|0.61055446569467375|00028400047678|SNACKS|G1 GROCERY|-81.027334|1.4141937624131469|149|2
34.977331|14a7164b866968a01c259b003b07b6bf274f1b8e|9.7|2014-12-29 14:55:00|1.41290891556208|3|7790011553|149|0.6104695895098807|0|33|361|-81.027334|105|34.977331|BREAKFAST SAUSAGE|3.0300000000000002|19|JIMMY DEAN MILD SAUSAGE|67e73b6075b00299fbe43b733da4006ae51c2ec2|6.232193769327634|0.61055446569467375|00077900115530|BREAKFAST SAUSAGE|CASE READY MEATS|-81.027334|1.4141937624131469|149|2
34.977331|54a075a6589542d7c7f4daa968cd2a7aff2f8277|4.29|2014-12-26 16:43:00|1.41290891556208|3|4178000011|149|0.6104695895098807|0|33|201|-81.027334|31|34.977331|POTATO CHIPS|1.79|1|UTZ RED FAT SC & O RIPPLE CHIP|67e73b6075b00299fbe43b733da4006ae51c2ec2|6.232193769327634|0.61055446569467375|00041780000668|SNACKS|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|b5c5a33a9857ce2ba3b9bbb753d0025c43ef94d1|4.29|2014-09-12 12:35:00|1.41290891556208|3|4178000011|149|0.6104695895098807|0|33|201|-81.027334|31|34.977331|POTATO CHIPS|1.79|1|UTZ REGULAR POTATO CHIPS|67e73b6075b00299fbe43b733da4006ae51c2ec2|6.232193769327634|0.61055446569467375|00041780000118|SNACKS|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|717190fc49c21ebf862438abc0d543a3c2221e54|3.99|2015-02-03 20:21:00|1.41290891556208|3|7203670998|149|0.6104695895098807|0|33|31|-81.027334|4|34.977331|NON CARBONATED WATER|0.0|1|HT PURIFIED WATER 8 OZ 24PK|67e73b6075b00299fbe43b733da4006ae51c2ec2|6.232193769327634|0.61055446569467375|00072036709981|BOTTLED WATER|G1 GROCERY|-81.027334|1.4141937624131469|149|1
34.977331|9de23bc5d15fd345b613de799f88b786ff2b405c|36.99|2014-12-29 14:51:00|1.41290891556208|3|82061603122|149|0.6104695895098807|0|33|7287|-81.027334|1600|34.977331|CHRISTMAS PLUSH IMP|27.74|18|"I/O 15"" ROUND ANIMALS"|67e73b6075b00299fbe43b733da4006ae51c2ec2|6.232193769327634|0.61055446569467375|00820616031225|SEASONAL MERCHANDISE|GM|-81.027334|1.4141937624131469|149|1
34.977331|f2ae53f04d336eec968235ca15555bbff3a2fe67|36.99|2014-12-29 14:51:00|1.41290891556208|3|82061603122|149|0.6104695895098807|0|33|7287|-81.027334|1600|34.977331|CHRISTMAS PLUSH IMP|27.74|18|"I/O 15"" ROUND ANIMALS"|67e73b6075b00299fbe43b733da4006ae51c2ec2|6.232193769327634|0.61055446569467375|00820616031225|SEASONAL MERCHANDISE|GM|-81.027334|1.4141937624131469|149|1
34.977331|aabe35a8bbc83bc10885cdff8e76015ecbc58366|23.98|2014-12-31 17:20:00|1.41290891556208|3|2301286481|149|0.6104695895098807|0|33|1477|-81.027334|485|34.977331|SUSHI HYBRID|0.0|6|"CHEF SAMPLER ""A"""|67e73b6075b00299fbe43b733da4006ae51c2ec2|6.232193769327634|0.61055446569467375|00023012864811|SUSHI|DELI|-81.027334|1.4141937624131469|149|2
35.106477|811597fd640ef67ff48805778d61db8c5487a5e8|3.59|2014-11-24 12:10:00|80.806073375020532|2|7341003205|4|35.114108445221994|0|0|1029|-80.824767|162|35.116751|RYE/PUMP|0.0|7|ARN JEWISH RYE PLAIN PP|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00073410032008|SLICED BREAD|COMMERCIAL BAKERY|-80.806073|80.806073208986547|294|1
35.106477|3c7a1081dcdce0be4f00a83988d8b044901d4852|3.59|2014-09-19 18:22:00|80.806073375020532|2|7341016305|4|35.114108445221994|0|0|1035|-80.824767|163|35.116751|SANDWICH ROLL|0.6|7|ARN SELECT 100% WHEAT HAMS PP|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00073410161456|BUNS/ROLLS|COMMERCIAL BAKERY|-80.806073|80.806073208986547|294|1
35.106477|4bba72c768ad4af8a27f624033cb72277fff7c28|2.59|2015-03-06 17:42:00|80.806073375020532|2|7680853357|4|35.114108445221994|0|0|1208|-80.824767|23|35.116751|WHSE PASTA VALUE ADD|0.0|1|BARILLA PLUS SPAGHETTI|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00076808533576|PASTA|G1 GROCERY|-80.806073|80.806073208986547|294|1
35.106477|8e8a3d838710f3adeda41e0317d010a1c53f8c20|3.49|2015-02-20 17:36:00|80.806073375020532|2|7797509132|4|35.114108445221994|0|0|202|-80.824767|31|35.116751|PRETZELS|0.49|1|SOH POPPERS CINN SUGAR|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00077975091449|SNACKS|G1 GROCERY|-80.806073|80.806073208986547|294|1
35.106477|4d5dd74907e523eed16a03097165a64f1412cb3d|3.79|2015-01-16 18:24:00|80.806073375020532|2||4|35.114108445221994|0|0|539|-80.824767|64|35.116751|FRESH CAULIFLOWER|0.0|4|WHT CAULIFLOWER 12'S(RPC)|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00204079000002|FRESH PRODUCE|PRODUCE|-80.806073|80.806073208986547|294|1
35.106477|3ebc8f8213731d42f186035fadc100600cadb9af|3.0|2014-09-13 18:05:00|80.806073375020532|2||4|35.114108445221994|0|0|531|-80.824767|64|35.116751|FRESH CORN|0.2|4|COO YELLOW CORN|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00204078000003|FRESH PRODUCE|PRODUCE|-80.806073|80.806073208986547|294|5
35.106477|0d406489c57e15f7ef4116d2a76ffd86e325ef55|3.0|2014-09-26 16:14:00|80.806073375020532|2||4|35.114108445221994|0|0|531|-80.824767|64|35.116751|FRESH CORN|0.0|4|COO YELLOW CORN|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00204078000003|FRESH PRODUCE|PRODUCE|-80.806073|80.806073208986547|294|5
35.106477|5d434ec3d04a23b039e26767a655d458e4113f2d|3.0|2014-10-09 17:22:00|80.806073375020532|2||4|35.114108445221994|0|0|531|-80.824767|64|35.116751|FRESH CORN|0.0|4|COO YELLOW CORN|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00204078000003|FRESH PRODUCE|PRODUCE|-80.806073|80.806073208986547|294|5
35.106477|6b8ae430355246fa83678438959d5acc92733d21|3.0|2014-11-14 18:19:00|80.806073375020532|2||4|35.114108445221994|0|0|531|-80.824767|64|35.116751|FRESH CORN|0.0|4|COO YELLOW CORN|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00204078000003|FRESH PRODUCE|PRODUCE|-80.806073|80.806073208986547|294|5
35.106477|392a2fb299ae9306987ac19012d9f2886123c273|1.6|2015-01-30 17:53:00|80.806073375020532|2||4|35.114108445221994|0|0|531|-80.824767|64|35.116751|FRESH CORN|0.0|4|COO YELLOW CORN|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00204078000003|FRESH PRODUCE|PRODUCE|-80.806073|80.806073208986547|294|2
35.106477|eac17f9d5ac7bc8f5b58e1ae71d052ca3be424e9|3.2|2015-02-25 14:37:00|80.806073375020532|2||4|35.114108445221994|0|0|531|-80.824767|64|35.116751|FRESH CORN|0.0|4|COO YELLOW CORN|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00204078000003|FRESH PRODUCE|PRODUCE|-80.806073|80.806073208986547|294|4
35.106477|c20104875fdd1c7936a3fd88881b7276b02656c0|3.49|2015-02-28 17:46:00|80.806073375020532|2||4|35.114108445221994|0|0|539|-80.824767|64|35.116751|FRESH CAULIFLOWER|0.99|4|WHT CAULIFLOWER 12'S(RPC)|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00204079000002|FRESH PRODUCE|PRODUCE|-80.806073|80.806073208986547|294|1
35.106477|62655c9c35d4df206382aeffd62845423cfc8451|2.69|2015-01-24 14:36:00|80.806073375020532|2|7512800016|4|35.114108445221994|0|0|1273|-80.824767|50|35.116751|BAG VEG NON STEAM|0.7|5|SAVANNAH SWT CORN HUSHPUPPY|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00075128000126|VEGETABLES-FROZEN|FROZEN|-80.806073|80.806073208986547|294|1
35.106477|f9800d2d807aff242054754a45a66e79089d2438|3.49|2014-12-11 17:30:00|80.806073375020532|2|75733955555|4|35.114108445221994|0|0|68|-80.824767|11|35.116751|BARBECUE SAUCES|0.51|1|STICKY FNGR BBQ SC TENN WHISKY|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00757339777775|CONDIMENTS|G1 GROCERY|-80.806073|80.806073208986547|294|1
35.106477|b33e638a67fb20199752462c511c621745663467|3.49|2014-12-20 18:28:00|80.806073375020532|2|75733955555|4|35.114108445221994|0|0|68|-80.824767|11|35.116751|BARBECUE SAUCES|0.51|1|STICKY FNGR BBQ SC TENN WHISKY|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00757339777775|CONDIMENTS|G1 GROCERY|-80.806073|80.806073208986547|294|1
35.106477|acc162d5aeda964a5ab4a656366dd9287f2bb5d1|1.39|2014-11-21 18:11:00|80.806073375020532|2|5210094269|4|35.114108445221994|0|0|80|-80.824767|34|35.116751|SEASONING PACKETS|0.39|1|E  MC CHILI SEASONING MIX|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00052100091501|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.806073|80.806073208986547|294|1
35.106477|ea5f72926cc182c2aeb7aa897a69a692f4d18806|1.39|2014-10-03 14:36:00|80.806073375020532|2|5210094269|4|35.114108445221994|0|0|80|-80.824767|34|35.116751|SEASONING PACKETS|0.39|1|E  MC CHILI SEASONING MIX|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00052100091501|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.806073|80.806073208986547|294|1
35.106477|a5f55a61937ef90ddd13118d6438a98dbfae3e0d|12.0|2014-11-25 16:36:00|80.806073375020532|2|66440100015|4|35.114108445221994|0|0|1165|-80.824767|87|35.116751|NFS-FRESH CONSUMER BUNCH|0.0|9|BUNCH- HYPERIUCM ASST.|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00664401000153|FLORAL|FLORAL|-80.806073|80.806073208986547|294|3
35.106477|584ed5f8229c9ea132815879f9a9c898cfb63006|1.49|2015-01-02 18:23:00|80.806073375020532|2|7203653022|4|35.114108445221994|0|0|1273|-80.824767|50|35.116751|BAG VEG NON STEAM|0.5|5|HT CROWDER PEAS|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00072036530172|VEGETABLES-FROZEN|FROZEN|-80.806073|80.806073208986547|294|1
35.106477|cef51651e8b7ac307e49318997992f678343467e|15.98|2015-02-13 15:15:00|80.806073375020532|2|2840000288|4|35.114108445221994|0|0|205|-80.824767|31|35.116751|REMAINING SNACKS|4.0|1|FRITOLAY CLASSIC 20 CTN|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00028400002882|SNACKS|G1 GROCERY|-80.806073|80.806073208986547|294|2
35.106477|afd56572b2882e795c25bc19130f4ac6f39dfbac|1.89|2014-10-31 16:32:00|80.806073375020532|2|2700038249|4|35.114108445221994|0|0|70|-80.824767|11|35.116751|KETCHUP|0.0|1|HUNTS KETCHUP 24|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00027000382493|CONDIMENTS|G1 GROCERY|-80.806073|80.806073208986547|294|1
35.106477|fa71964046fefde830a68d261ea94f04a7cec7ed|10.99|2014-12-05 15:15:00|80.806073375020532|2|7203683001|4|35.114108445221994|0|0|352|-80.824767|110|35.116751|IQF CHICKEN|2.51|19|HT 2.5 LB CHICKEN TENDR BRST|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00072036830029|FROZEN CASE MEAT|CASE READY MEATS|-80.806073|80.806073208986547|294|1
35.106477|3d36baaf46870b990e2e339b898bb8dd5d41ea56|2.27|2015-02-07 17:04:00|80.806073375020532|2|7203656065|4|35.114108445221994|0|0|315|-80.824767|52|35.116751|CHEESE-PROCESSED-SLICED|0.0|3|HT 2% SINGLE WRAP CHEESE|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00072036600844|CHEESE|DAIRY|-80.806073|80.806073208986547|294|1
35.106477|95f1cd7dbdbe9bbed34283f4f534a859a2bb871f|2.27|2015-01-09 18:02:00|80.806073375020532|2|7203656065|4|35.114108445221994|0|0|315|-80.824767|52|35.116751|CHEESE-PROCESSED-SLICED|0.0|3|HT 2% SINGLE WRAP CHEESE|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00072036600844|CHEESE|DAIRY|-80.806073|80.806073208986547|294|1
35.106477|f3df5b27abb48b939403a78fe0a8f10f6f8ea6f3|4.49|2014-12-06 14:36:00|80.806073375020532|2|7824500008|4|35.114108445221994|0|0|184|-80.824767|28|35.116751|SALAD DRESSINGS-LIQUID|0.5|1|HENDRICK DRS VIN SWEET ITALIAN|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00078245000055|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.806073|80.806073208986547|294|1
35.106477|0558e22af46c73f80da2b03f6fafadb0f6de0334|6.98|2015-02-06 16:28:00|80.806073375020532|2|3760011544|4|35.114108445221994|0|0|175|-80.824767|27|35.116751|CANNED MEATS|1.98|1|SPAM LITE 12 OZ|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00037600175340|PREPARED FOODS-RTS|G1 GROCERY|-80.806073|80.806073208986547|294|2
35.106477|f6eaef67dd91b39e20998a7bf7afdb7b93060e08|3.99|2014-12-27 18:20:00|80.806073375020532|2||4|35.114108445221994|0|0|506|-80.824767|64|35.116751|FRESH MELONS|0.0|4|CANTALOUPES, JUMBO|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00204050000007|FRESH PRODUCE|PRODUCE|-80.806073|80.806073208986547|294|1
35.106477|050e3a688234349c48951b54265c36b166509b56|2.99|2014-10-15 15:47:00|80.806073375020532|2|8186420216|4|35.114108445221994|0|0|583|-80.824767|136|35.116751|NUTS|0.0|4|ROASTED PEANUTS IN-SHELL|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00081864222166|OTHER MERCHANDISE|PRODUCE|-80.806073|80.806073208986547|294|1
35.106477|e191f2ca1611e8ca997a3c1282b1689bf4914722|2.99|2014-10-07 17:07:00|1.4091206135396188|2|8186420216|4|0.6127236124256613|0|47|583|-80.806073|136|35.106477|NUTS|0.0|4|ROASTED PEANUTS IN-SHELL|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|0.61242566243833529|00081864222166|OTHER MERCHANDISE|PRODUCE|-80.806073|1.4103320294568917|4|1
35.106477|9a911e09affdfa1c0041adb1df7b6cd67d9c0d64|5.99|2014-11-11 16:42:00|80.806073375020532|2|7203688216|4|35.114108445221994|0|0|500|-80.824767|64|35.116751|FRESH APPLES|0.0|4|HT HONEYCRISP APPLE 3LB|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00072036882165|FRESH PRODUCE|PRODUCE|-80.806073|80.806073208986547|294|1
35.106477|f55b383b6317420f8ed89a19d7ff52d064f41b7d|2.31|2014-09-30 17:50:00|80.806073375020532|2||4|35.114108445221994|0|0|501|-80.824767|64|35.116751|FRESH PEARS|0.35|4|BOSC PEARS|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00204413000002|FRESH PRODUCE|PRODUCE|-80.806073|80.806073208986547|294|1
35.106477|36dedc24d45033023660dddc407d1f957b6efe73|5.69|2014-09-20 16:29:00|80.806073375020532|2|7756725423|4|35.114108445221994|0|0|252|-80.824767|45|35.116751|PREMIUM ICE CREAM|2.85|5|BREYER'S LACTOSE FREE VAN|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00077567227003|ICE CREAM|FROZEN|-80.806073|80.806073208986547|294|1
35.106477|3c841657deb45d48f98b8382a8bd527c7286ea79|4.99|2014-10-26 15:23:00|80.806073375020532|2|3338307764|4|35.114108445221994|0|0|500|-80.824767|64|35.116751|FRESH APPLES|0.0|4|GALA APPLES 3LB BAG|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00072036880314|FRESH PRODUCE|PRODUCE|-80.806073|80.806073208986547|294|1
35.106477|4bb94970de322c2ddb9b66cc42a7a65188104240|0.38|2014-12-03 17:42:00|80.806073375020532|2||4|35.114108445221994|0|0|502|-80.824767|64|35.116751|FRESH BANANAS|0.0|4|BANANAS, YELLOW|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00204011000008|FRESH PRODUCE|PRODUCE|-80.806073|80.806073208986547|294|1
35.106477|860d9bcdf838153fdae039a162333b513cad0305|0.73|2015-01-24 14:40:00|80.806073375020532|2||4|35.114108445221994|0|0|502|-80.824767|64|35.116751|FRESH BANANAS|0.0|4|BANANAS, YELLOW|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00204011000008|FRESH PRODUCE|PRODUCE|-80.806073|80.806073208986547|294|1
35.106477|0940f465d92af2ea53646e84e12cbe886c30ec25|1.1|2014-11-10 12:49:00|80.806073375020532|2||4|35.11410844522382|0|0|502|-80.78468|64|35.096737|FRESH BANANAS|0.0|4|BANANAS, YELLOW|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00204011000008|FRESH PRODUCE|PRODUCE|-80.806073|80.806073043302163|30|1
35.106477|548593c75f48734a2bcef542b0f3273eaf177482|1.25|2015-02-12 12:30:00|80.806073375020532|2|5100002421|4|35.114108445221994|0|0|214|-80.824767|33|35.116751|BROTH|0.0|1|SWANSON BROTH LOW SOD BEEF|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00051000142979|SOUP|G1 GROCERY|-80.806073|80.806073208986547|294|1
35.106477|cd53d089304e523f60d4376a76829845d31e0ea4|4.0|2014-12-05 15:25:00|80.806073375020532|2|4300000953|4|35.114108445221994|0|0|272|-80.824767|307|35.116751|TOPPINGS FROZEN|1.0|5|COOL WHIP WHIPPED TOPPING|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00043000009536|DESSERTS FROZEN|FROZEN|-80.806073|80.806073208986547|294|2
35.106477|e923fc52bf248fcd139caa30a85ef911e694a8f1|3.76|2015-02-03 16:27:00|80.806073375020532|2|20394300000|4|35.114108445221994|0|0|643|-80.824767|137|35.116751|PORK OFFALS-FROZEN|0.0|2|MORTY PRIDE SMOKED HOCKS|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00203943000001|PORK|MEAT|-80.806073|80.806073208986547|294|1
35.106477|9044f8a82380bc975239c42c9160c7eb9dff8647|11.14|2014-11-19 14:31:00|80.806073375020532|2|20194700000|4|35.114108445221994|0|0|299|-80.824767|49|35.116751|ANGUS BEEF|0.0|2|ANGUS BEEF BNLS SHOULDER ROAST|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00201947000003|BEEF|MEAT|-80.806073|80.806073208986547|294|1
35.106477|ae50a79f3decc6973477ee4c936d2cfb3b6d364e|8.95|2014-09-27 14:44:00|80.806073375020532|2|20194700000|4|35.114108445221994|0|0|299|-80.824767|49|35.116751|ANGUS BEEF|0.0|2|ANGUS BEEF BNLS SHOULDER ROAST|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00201947000003|BEEF|MEAT|-80.806073|80.806073208986547|294|1
35.106477|26e870394f9d7467a3eaa042583e1df702f75de3|9.94|2015-01-19 12:17:00|80.806073375020532|2|20194700000|4|35.114108445221994|0|0|299|-80.824767|49|35.116751|ANGUS BEEF|0.0|2|ANGUS BEEF BNLS SHOULDER ROAST|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00201947000003|BEEF|MEAT|-80.806073|80.806073208986547|294|1
35.106477|8f6baec7d21ae1e14d5d4616327d94f3fb3e259b|2.19|2014-11-20 13:28:00|80.806073375020532|2|1330018301|4|35.114108445221994|0|0|100|-80.824767|15|35.116751|CORN MEAL|0.0|1|MW BTTRMILK CORN MEAL MIX SR|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00013300183014|FLOUR|G1 GROCERY|-80.806073|80.806073208986547|294|1
35.106477|33aab79eeae28130c43747f36ca653d5d9114483|1.39|2014-12-24 13:37:00|80.806073375020532|2|3470001211|4|35.114108445221994|0|0|247|-80.824767|39|35.116751|VEGETABLES-FLANKER|0.0|1|ALLEN ITALIAN GREEN BEAN 15|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00034700012117|VEGETABLES-CAN/JAR|G1 GROCERY|-80.806073|80.806073208986547|294|1
35.106477|4332175bd3d1802c86ccf72fbcc574c0924eb6b0|1.13|2014-11-25 14:35:00|80.806073375020532|2||4|35.11410844522382|0|0|522|-80.78468|64|35.096737|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00204664000004|FRESH PRODUCE|PRODUCE|-80.806073|80.806073043302163|30|1
35.106477|ab911457fecb5697de3c39016b477102b6be0dae|1.79|2014-12-16 17:46:00|80.806073375020532|2|7203663220|4|35.114108445221994|0|0|330|-80.824767|55|35.116751|EGGS|0.0|3|HT GRADE A    LARGE EGGS|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00072036632203|EGGS FRESH|DAIRY|-80.806073|80.806073208986547|294|1
35.106477|20eb4cf893ae3608e56993aa0dd3e180e64e6920|5.91|2014-12-10 14:20:00|80.806073375020532|2|20579000000|4|35.114108445162479|0|0|1824|-80.85753|410|35.116638|BH LOAVES|0.0|6|BOARS HEAD LOWER SODIUM BOLGNA|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00205790000005|BH MEAT|DELI|-80.806073|80.806074183674468|204|1
35.106477|ba7364e3ac6ad5b5c342421234df01ee1c4399be|2.99|2014-12-05 17:45:00|80.806073375020532|2|4069503007|4|35.114108445221994|0|0|555|-80.824767|64|35.116751|PACKAGED SALADS|0.0|4|ROMIANE HEARTS|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00033383651620|FRESH PRODUCE|PRODUCE|-80.806073|80.806073208986547|294|1
35.106477|bcb52b2639f8042e9e6e98fdab0c57ced4a893b8|5.99|2014-12-16 17:03:00|80.806073375020532|2|20496400000|4|35.114108445162479|0|0|756|-80.85753|87|35.116638|NFS-FLORAL ACCESSORIES|0.0|9|*ACCESSORIES|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00204964000001|FLORAL|FLORAL|-80.806073|80.806074183674468|204|1
35.106477|e6db8062e620f2503a355bb944f0cd479708defa|3.19|2015-01-12 17:26:00|80.806073375020532|2|4060034500|4|35.114108445221994|0|0|313|-80.824767|51|35.116751|MARGARINE|0.0|3|ICBINB COOKING AND BAKING STIC|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00040600034166|BUTTER & MARGARINE|DAIRY|-80.806073|80.806073208986547|294|1
35.106477|e86b44d81b726eac10c3a30de3fde9cb5311a6ee|3.19|2014-11-26 17:56:00|80.806073375020532|2|4060034500|4|35.114108445221994|0|0|313|-80.824767|51|35.116751|MARGARINE|0.0|3|ICBINB COOKING AND BAKING STIC|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00040600034166|BUTTER & MARGARINE|DAIRY|-80.806073|80.806073208986547|294|1
35.106477|28ad3725f01df90415dbe074385e0b510dece5d6|2.65|2014-09-20 16:09:00|80.806073375020532|2|4530000549|4|35.114108445162479|0|0|125|-80.85753|19|35.116638|PEANUT BUTTER|0.0|1|PETER PAN RF CREAMY PBUTTER|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00045300005447|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.806073|80.806074183674468|204|1
35.106477|d1e9a854a9368b1d1bcc8c9708d847de50d751a3|3.15|2015-02-10 17:34:00|80.806073375020532|2|7225003712|4|35.114108445221994|0|0|1026|-80.824767|162|35.116751|WHEAT|0.0|7|NATOWN 100% WHEAT BRD|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00072250037129|SLICED BREAD|COMMERCIAL BAKERY|-80.806073|80.806073208986547|294|1
35.106477|6305d1db2601fc564af505718b324e0001d9e527|6.3|2014-11-12 16:19:00|80.806073375020532|2|7225003712|4|35.114108445221994|0|0|1026|-80.824767|162|35.116751|WHEAT|1.57|7|NATOWN 100% WHEAT BRD|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00072250037129|SLICED BREAD|COMMERCIAL BAKERY|-80.806073|80.806073208986547|294|2
35.106477|d6502c409ca2fce509f0adf376b18d614baabbbd|1.39|2014-09-15 15:22:00|80.806073375020532|2|7020001063|4|35.114108445221994|0|0|22|-80.824767|28|35.116751|CROUTONS|0.0|1|TEXAS CROUTON SEASONED|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00070200010659|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.806073|80.806073208986547|294|1
35.106477|fdbe4971ab4bde15a1c51eac4c5ee79e8a113f5a|35.22|2014-12-13 14:18:00|1.4091206135396188|2|20165900000|4|0.6127236124256613|0|47|297|-80.806073|49|35.106477|GROUND BEEF|0.0|2|GROUND BEEF 93% LEAN|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|0.61242566243833529|00201659000001|BEEF|MEAT|-80.806073|1.4103320294568917|4|6
35.106477|a82965a39991bccc04437f0e2b9b29d90d725c6f|2.59|2014-09-24 12:53:00|80.806073375020532|2|5100017520|4|35.114108445221994|0|0|1201|-80.824767|33|35.116751|RTS CANNED|1.09|1|CAM HOMESTYLE HR WG PSTA FAGIO|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00051000195692|SOUP|G1 GROCERY|-80.806073|80.806073208986547|294|1
35.106477|309813732e48fccc0cde0ec220e61d1481139595|0.97|2015-02-20 18:32:00|80.806073375020532|2|7203698757|4|35.114108445221994|0|0|31|-80.824767|4|35.116751|NON CARBONATED WATER|0.0|1|HT DISTILLED WATER|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00072036360601|BOTTLED WATER|G1 GROCERY|-80.806073|80.806073208986547|294|1
35.106477|4a97c9dd21d34dea7736d47881184c351a0256bc|2.35|2014-10-30 16:44:00|80.806073375020532|2||4|35.114108445221994|0|0|536|-80.824767|64|35.116751|FRESH SQUASH|0.0|4|COO ZUCCHINI SQUASH, FANCY|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00204067000007|FRESH PRODUCE|PRODUCE|-80.806073|80.806073208986547|294|1
35.106477|e4f1b3d9276d36483e8734c38185247b8b508282|4.99|2014-12-11 17:40:00|80.806073375020532|2|7244010400|4|35.114108445221994|0|0|6787|-80.824767|1568|35.116751|MAGAZINES MONTHLY|0.0|18|SOUTHERN LIVING|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00072440104006|MAGAZINES|GM|-80.806073|80.806073208986547|294|1
35.106477|77d68aae79196002cb5a32416f19ce75bea37993|3.69|2014-11-26 21:07:00|80.806073375020532|2|1258700020|4|35.114108445221994|0|0|444|-80.824767|76|35.116751|NFS-PLASTIC WRAPS|0.69|1|GLAD WRAP|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00012587000205|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.806073|80.806073208986547|294|1
35.106477|4a8088a3c180e2752b8aa3755ac97af43b7eaf19|6.99|2014-10-28 15:08:00|80.806073375020532|2||4|35.114108445221994|0|0|1347|-80.824767|64|35.116751|PUMPKINS|1.99|4|CARVING PUMPKINS, LARGE|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00204737000009|FRESH PRODUCE|PRODUCE|-80.806073|80.806073208986547|294|1
35.106477|9ad0cc5e4dd81901f668ce6a89cf2105fc23f6cd|2.85|2014-11-16 17:08:00|80.806073375020532|2|7203656061|4|35.114108445221994|0|0|320|-80.824767|53|35.116751|COTTAGE CHEESE|0.35|3|HT LOW FAT COTTAGE CHEESE|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00072036560636|CULTURES|DAIRY|-80.806073|80.806073208986547|294|1
35.106477|44a67143dfc10107c56aa2e08c6c66df7033246a|3.29|2015-02-11 12:46:00|80.806073375020532|2|7225000486|4|35.11410844302619|0|0|1034|-80.80146|163|35.17739|HOT DOG|0.0|7|NATOWN 100% WHEAT HD BUNS|68e685d2c1e6c0fed622e098ebc72efc70f7af28|0.5273144356914982|35.114108445179689|00072250004862|BUNS/ROLLS|COMMERCIAL BAKERY|-80.806073|80.806080079877972|208|1
35.04711|8b780306d7bad1b9a5c9c81e8a4cdd704e1e9f35|1.79|2014-12-22 18:01:00|80.648225123995502|4||129|35.075900011657374|0|30|502|-80.709466|64|35.124987|FRESH BANANAS|0.0|4|BANANAS, YELLOW|6ebb35822a525b11870b63f1fce58381f329f69b|1.9893205637554092|35.078006462436761|00204011000008|FRESH PRODUCE|PRODUCE|-80.64817|80.648188781722752|157|1
35.04711|75234cbad7a05fe84fec9148a1541d74ab3f9bb2|1.18|2014-11-15 18:39:00|80.648225123995502|4||129|35.075900011657374|0|30|502|-80.709466|64|35.124987|FRESH BANANAS|0.0|4|BANANAS, YELLOW|6ebb35822a525b11870b63f1fce58381f329f69b|1.9893205637554092|35.078006462436761|00204011000008|FRESH PRODUCE|PRODUCE|-80.64817|80.648188781722752|157|1
35.04711|4571042310954932d957883e33cfe9e3edf625de|6.49|2014-10-26 18:03:00|1.4091206135396188|4|7203688056|129|0.6116874628086298|0|47|562|-80.64817|64|35.04711|FRESH CUT FRUIT|0.0|4|HT MIXED FRUIT CHUNKS 32OZ|6ebb35822a525b11870b63f1fce58381f329f69b|1.9893205637554092|0.61242566243833529|00072036880567|FRESH PRODUCE|PRODUCE|-80.64817|1.407576102208115|129|1
35.04711|51efdc17d3e911c54954a53c2c81259013f8e3b7|9.98|2014-10-26 18:04:00|1.4091206135396188|4|71575620002|129|0.6116874628086298|0|47|504|-80.64817|64|35.04711|FRESH BERRIES|2.5|4|STRAWBERRIES 1LB CLAM|6ebb35822a525b11870b63f1fce58381f329f69b|1.9893205637554092|0.61242566243833529|00071430007525|FRESH PRODUCE|PRODUCE|-80.64817|1.407576102208115|129|2
35.172688|d6bd8c149a11fea38479289b0b496a51cf5bb287|2.29|2014-11-20 15:49:00|80.632521683083056|4|7203695175|474|35.200890600085224|0|39|1607|-80.66939|371|35.28326|FROZEN DOUGH (BREAD)|0.0|14|FRESH LRG FRENCH BREAD|732d336cb2f5ae52a0796a84326f295a7900162a|1.9487327675272896|35.177497916598789|00072036951755|BREAD|BAKERY|-80.661096|80.661134430684854|46|1
35.172688|467dde7cd430f1679df04aedcf14e1ab696a9c1f|6.85|2014-11-28 09:39:00|1.4094857484078087|4|7192147763|474|0.6138792123766993|0|26|284|-80.661096|892|35.172688|SUPER PREMIUM PIZZA|0.0|5|12in CPK TC MARGHERITA PIZZA|732d336cb2f5ae52a0796a84326f295a7900162a|1.9487327675272896|0.61471665291522548|00071921290535|FROZEN PIZZA|FROZEN|-80.661096|1.407801703467228|474|1
35.172688|5e3dd67066a3c10a6a5bcbfe4ff7372bcf52feb2|2.19|2014-09-29 18:13:00|80.632521683083056|4|1200000230|474|35.200890616948811|0|39|55|-80.70901|8|35.17335|REGULAR|0.69|23|MT DEW CODE RED  2 LTR|732d336cb2f5ae52a0796a84326f295a7900162a|1.9487327675272896|35.177497916598789|00012000105425|CARBONATED BEVERAGES|BEVERAGE|-80.661096|80.661103269991628|174|1
35.444064|2ceaf84a10b4acbd55296ab16f9ddf0604054480|3.69|2015-01-20 15:31:00|1.4102725052409182|2|7518500700|121|0.6186156170875914|0|1|1030|-80.995484|162|35.444064|SLICED BREAD POTATO|0.0|7|MARTINS POTATO BREAD|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00075185007007|SLICED BREAD|COMMERCIAL BAKERY|-80.995484|1.413637875046387|121|1
35.444064|7d3de575c7c858dbd8bdcd008e75aa4f724c4a34|3.69|2014-11-12 16:39:00|1.4102725052409182|2|7518500700|121|0.6186156170875914|0|1|1030|-80.995484|162|35.444064|SLICED BREAD POTATO|0.0|7|MARTINS POTATO BREAD|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00075185007007|SLICED BREAD|COMMERCIAL BAKERY|-80.995484|1.413637875046387|121|1
35.444064|3852a54c90d7fe3a765e00bdd651347dfedacb46|1.49|2015-02-12 10:29:00|1.4102725052409182|2|8265733412|121|0.6186156170875914|0|1|31|-80.995484|4|35.444064|NON CARBONATED WATER|0.24|1|DEER PARK WATER 3LT|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00082657334127|BOTTLED WATER|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|4b374b417b7446ffaf6af6e0687da5983fb7cb55|5.49|2015-03-05 14:00:00|1.4102725052409182|2|8298800006|121|0.6186156170875914|0|1|1276|-80.995484|279|35.444064|FROZEN SANDWICHES|0.0|5|WHITE CASTLE M/W CHEESEBURGER|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00082988010066|FROZEN SANDWICH AND SNACKS|FROZEN|-80.995484|1.413637875046387|121|1
35.444064|031a215061502fd1fde1243d2f058afc33a41fe2|4.83|2015-01-19 12:29:00|1.4102725052409182|2|20165500000|121|0.6186156170875914|0|1|297|-80.995484|49|35.444064|GROUND BEEF|0.0|2|HT PREMIUM GRND BEEF 80% LEAN|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00201655000005|BEEF|MEAT|-80.995484|1.413637875046387|121|1
35.444064|66d2c094b9f1637fcf558550102c2c79a296b5a2|5.96|2015-01-12 09:54:00|1.4102725052409182|2|8265733412|121|0.6186156170875914|0|1|31|-80.995484|4|35.444064|NON CARBONATED WATER|0.96|1|DEER PARK WATER 3LT|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00082657334127|BOTTLED WATER|G1 GROCERY|-80.995484|1.413637875046387|121|4
35.444064|9bd6b2a63910e1f70b25f3e5b8d6e47cf8618be2|5.49|2014-12-08 09:43:00|1.4102725052409182|2|8298800006|121|0.6186156170875914|0|1|1276|-80.995484|279|35.444064|FROZEN SANDWICHES|0.0|5|WHITE CASTLE M/W CHEESEBURGER|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00082988010066|FROZEN SANDWICH AND SNACKS|FROZEN|-80.995484|1.413637875046387|121|1
35.444064|819821d2216a75803e917a30afa1bc58f261b0a2|1.78|2015-01-02 17:39:00|1.4102725052409182|2||121|0.6186156170875914|0|1|532|-80.995484|64|35.444064|FRESH CUCUMBERS|0.0|4|COO CUCUMBERS S/S|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00204062000002|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|2
35.444064|19b937f387ac1b54ee7b6b05223c00863cacb131|3.83|2014-12-18 18:12:00|1.4102725052409182|2|20165500000|121|0.6186156170875914|0|1|297|-80.995484|49|35.444064|GROUND BEEF|0.0|2|HT PREMIUM GRND BEEF 80% LEAN|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00201655000005|BEEF|MEAT|-80.995484|1.413637875046387|121|1
35.444064|8e10f323bf7a63fd2290432e15b8281cb18808aa|7.99|2014-10-15 13:22:00|1.4102725052409182|2|2100061161|121|0.6186156170875914|0|1|314|-80.995484|52|35.444064|CHEESE-PROCESSED-OTHER|0.0|3|KRAFT VELVEETA CHEESE|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00021000611614|CHEESE|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|d259056492f5b2c569889fd1c38a1731d02bcf70|7.99|2014-12-27 19:04:00|1.4102725052409182|2|1820000956|121|0.6186156170875914|0|1|457|-80.995484|82|35.444064|DOMESTIC SINGLES/SIX PACKS|0.0|16|MICHELOB LIGHT 6PK 12OZ BOTTLE|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00018200009563|DOMESTIC BEER|BEER|-80.995484|1.413637875046387|121|1
35.444064|9b6bc15f1a27cf077ff15a1faafd7e25a35a662f|4.99|2014-11-24 09:31:00|1.4102725052409182|2|2100061526|121|0.6186156170875914|0|1|315|-80.995484|52|35.444064|CHEESE-PROCESSED-SLICED|0.0|3|KRAFT SINGLE WRAP CHS|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00021000615261|CHEESE|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|ddf8802eb9633f5eb904df89d0b7458028ed11c4|3.39|2014-11-05 08:43:00|1.4102725052409182|2|1312000286|121|0.6186156170875914|0|1|1469|-80.995484|278|35.444064|REGULAR CUT FRIES|0.0|5|ORE-IDA CTRY STYLE HASH BROWNS|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00013120008337|FROZEN POTATO|FROZEN|-80.995484|1.413637875046387|121|1
35.444064|158ceeaa46d04e932457594298d0e4ce6afdc33a|3.99|2015-01-14 19:02:00|1.4102725052409182|2|4470003050|121|0.6186156170875914|0|1|840|-80.995484|102|35.444064|TUBS|0.49|19|OM DELI FRESH HONEY HAM|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00044700030547|LUNCHMEATS|CASE READY MEATS|-80.995484|1.413637875046387|121|1
35.444064|6e8d1a2995731228caf61786b88c52e9d9e844c1|3.59|2014-10-28 15:01:00|1.4102725052409182|2|4127100970|121|0.6186156170875914|0|1|341|-80.995484|57|35.444064|CREAMERS|0.3|3|I/O ITNAT'L PUMPKIN PIE SPICE|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00041271009705|MILK|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|12b282e1021a3d65704839e4b4f8ad1c77a05400|3.15|2014-09-12 13:06:00|1.4102725052409182|2|4127102564|121|0.6186156170875914|0|1|341|-80.995484|57|35.444064|CREAMERS|0.0|3|ITNAT'L FRENCH VANILLA|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00041271025644|MILK|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|77a681cbce38584bc6c73b57372d95d8e7cabc8e|3.25|2015-01-30 08:45:00|1.4102725052409182|2|4127102564|121|0.6186156170875914|0|1|341|-80.995484|57|35.444064|CREAMERS|0.48|3|ITNAT'L FRENCH VANILLA|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00041271025644|MILK|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|4528f79a43c007af32398e8aceeabe897b28b589|3.25|2015-02-24 14:56:00|1.4102725052409182|2|4127102564|121|0.6186156170875914|0|1|341|-80.995484|57|35.444064|CREAMERS|0.25|3|ITNAT'L FRENCH VANILLA|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00041271025644|MILK|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|5cdce94a05311b15dcd172dde26b0be4f117e6d9|3.49|2014-10-07 17:06:00|1.4102725052409182|2|4127102564|121|0.6186156170875914|0|1|341|-80.995484|57|35.444064|CREAMERS|0.49|3|ITNAT'L FRENCH VANILLA|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00041271025644|MILK|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|b90b985b9c4673984b5dbc73bb0fd3146ff563f1|3.25|2014-11-03 18:20:00|1.4102725052409182|2|4127102564|121|0.6186156170875914|0|1|341|-80.995484|57|35.444064|CREAMERS|0.25|3|ITNAT'L FRENCH VANILLA|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00041271025644|MILK|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|6ff4855da7609b89b6efa3b01324fa816aa063ec|3.25|2014-11-17 11:07:00|1.4102725052409182|2|4127102564|121|0.6186156170875914|0|1|341|-80.995484|57|35.444064|CREAMERS|0.0|3|ITNAT'L FRENCH VANILLA|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00041271025644|MILK|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|210b85c167027fc6573f85015616c7ae27369337|23.98|2014-11-20 12:03:00|1.4102725052409182|2|4300004648|121|0.6186156170875914|0|1|66|-80.995484|10|35.444064|GROUND CAN|6.0|1|MAXWELL HOUSE MASTER BLEND|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00043000046500|COFFEE|G1 GROCERY|-80.995484|1.413637875046387|121|2
35.444064|97586537c0467087601c5cf796f4bcbf09006d37|7.78|2014-09-19 15:46:00|1.4102725052409182|2|3800039125|121|0.6186156170875914|0|1|81|-80.995484|9|35.444064|RTE CEREAL KIDS|1.8|1|KELLOGG APPLE JACKS 8.7|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00038000391323|CEREAL|G1 GROCERY|-80.995484|1.413637875046387|121|2
35.444064|ae497b1e02319f16d5e09c49cc00497724cb5ea3|2.89|2014-11-13 14:06:00|1.4102725052409182|2|7203663102|121|0.6186156170875914|0|1|339|-80.995484|57|35.444064|EGGNOGS/DRINKS|0.39|3|I/O HARRIS TEETER EGG NOG|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00072036631022|MILK|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|2790c2bd1671870382e60cf96262027c6b036c5d|1.79|2015-01-07 17:05:00|1.4102725052409182|2|1800000261|121|0.6186156170875914|0|1|325|-80.995484|54|35.444064|BISCUITS-REFRIGERATED|0.0|3|GRANDS BUTTERMILK BISCUITS|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00018000001873|DOUGH PRODUCTS|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|5d21aba921bd1e27c0653306cb2faa3404c81445|2.69|2014-12-05 15:17:00|1.4102725052409182|2|7008506010|121|0.6186156170875914|0|1|1277|-80.995484|279|35.444064|FROZEN SNACKS|0.0|5|BAGEL BITES CHEESE & PEPP|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00070085060121|FROZEN SANDWICH AND SNACKS|FROZEN|-80.995484|1.413637875046387|121|1
35.444064|9bf9045d65c36afcb2129a81d44dc0f86111b5bf|7.99|2015-02-05 08:58:00|1.4102725052409182|2|2840000288|121|0.6186156170875914|0|1|205|-80.995484|31|35.444064|REMAINING SNACKS|1.0|1|FRITOLAY CLASSIC 20 CTN|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00028400002882|SNACKS|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.444064|3b2ea4247cae081e8fd24ef39fcdeb90ce6b5e73|12.99|2015-03-01 13:34:00|1.4102725052409182|2|7023666062|121|0.6186156170875914|0|1|751|-80.995484|87|35.444064|NFS-BOUQUETS|0.0|9|$12.99 SWEET SURPRIZE BOUQUET|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00070236660620|FLORAL|FLORAL|-80.995484|1.413637875046387|121|1
35.444064|ebed0d223d1bf88f69abdeaef56f95b048bfe736|3.58|2014-10-03 11:19:00|1.4102725052409182|2|5210003850|121|0.6186156170875914|0|1|80|-80.995484|34|35.444064|SEASONING PACKETS|0.0|1|MC BEEF STROGANOFF|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00052100038506|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.995484|1.413637875046387|121|2
35.444064|f5a218692bcb3fa1491611dc715c332fcf5f6a99|5.49|2014-10-10 14:27:00|1.4102725052409182|2|4900000548|121|0.6186156170875914|0|1|55|-80.995484|8|35.444064|REGULAR|1.32|23|CLASSIC COKE12OZ PET8PK FRDGPK|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00049000005486|CARBONATED BEVERAGES|BEVERAGE|-80.995484|1.413637875046387|121|1
35.444064|3fd68d6cce543c1c961169a9936991ef103a7005|5.99|2014-10-24 17:33:00|1.4102725052409182|2|7778200787|121|0.6186156170875914|0|1|355|-80.995484|104|35.444064|FRESH GRILLING SAUSAGE|0.0|19|JOHNSONVILLE BEER'N BRATWURST|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00077782007978|DINNER SAUSAGE|CASE READY MEATS|-80.995484|1.413637875046387|121|1
35.444064|5953db337d0571ccc25b86d893d27ba54c3434b7|0.99|2014-12-29 13:46:00|1.4102725052409182|2||121|0.6186156170875914|0|1|540|-80.995484|64|35.444064|FRESH CELERY|0.0|4|COO CELERY (RPC) 24'S|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00204070000001|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|2df2dc690b6fc584096b1bb4fe93027ab74096f9|1.99|2014-10-27 10:26:00|1.4102725052409182|2||121|0.6186156170875914|0|1|540|-80.995484|64|35.444064|FRESH CELERY|0.3|4|COO CELERY (RPC) 24'S|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00204070000001|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|efdb350ae1f2796d590fff27459b76de082d35fb|14.07|2014-09-24 17:14:00|1.4102725052409182|2|20332600000|121|0.6186156170875914|0|1|641|-80.995484|137|35.444064|PREMIUM PORK|2.03|2|VALUE PK BONE-IN PORK CHOPS|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00203326000000|PORK|MEAT|-80.995484|1.413637875046387|121|1
35.444064|0e0cde038401491224e4ebbbc71a160188c76ea5|1.37|2014-10-30 19:37:00|1.4102725052409182|2|7203626061|121|0.6186156170875914|0|1|719|-80.995484|10|35.444064|NFS-COFFEE FILTERS|0.0|1|HT 12 CUP BASKET FILTERS|74274279a5c20ba457e583b929cab76eddd12342|0.4026674255336212|0.61833652052202714|00072036260611|COFFEE|G1 GROCERY|-80.995484|1.413637875046387|121|1
35.06858|6c22ad972b5038cf9ddd35c9db7ac777acd022e6|3.99|2015-01-26 13:50:00|1.4091206135396188|1|75166677005|273|0.612062184999033|0|47|522|-80.7007|64|35.06858|FRESH TOMATOES|0.0|4|NATURESWEET CHERUBS 10.5 OZ|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00751666770058|FRESH PRODUCE|PRODUCE|-80.7007|1.4084929236641879|273|1
35.06858|3b8fe528a6aa8f1cbeae1ce2397db3bfd7c8bdab|1.0|2014-09-27 11:05:00|1.4091206135396188|1|78352054321|273|0.612062184999033|0|47|8598|-80.7007|1792|35.06858|NEWSPAPERS|0.0|18|DAILY  CHARLOTTE OBSERVER|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00783520543218|NEWSPAPERS|GM|-80.7007|1.4084929236641879|273|1
35.06858|6918b88dfe0b0b64a8913685c80c89f467e718f3|4.59|2015-02-13 15:09:00|1.4091206135396188|1|1600027569|273|0.612062184999033|0|47|81|-80.7007|9|35.06858|RTE CEREAL KIDS|1.59|1|GM LUCKY CHARMS 16OZ|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00016000275690|CEREAL|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|7cfb942e165979ad919c4ff1d76e0cf6f34c3498|2.99|2015-02-20 18:17:00|1.4091206135396188|1|7357529500|273|0.612062184999033|0|47|82|-80.7007|11|35.06858|VINEGAR|0.0|1|NAKANO VINEGAR RICE SEASONED|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00073575295003|CONDIMENTS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|bb805eabcef3cf146a4b04e6a7e94a39d21c99e4|8.45|2014-10-25 11:50:00|1.4091206135396188|1|7680828073|273|0.612062184999033|0|47|149|-80.7007|23|35.06858|WHSE PASTA CORE|0.0|1|BARILLA PASTA PENNE RIGATE|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00076808280739|PASTA|G1 GROCERY|-80.7007|1.4084929236641879|273|5
35.06858|928e25887120654020afe5479be6113edc5bd0ed|5.99|2014-12-29 17:35:00|80.700248323638462|1|9955508534|273|35.101654671114375|0|7|37|-80.732725|10|35.082768|PODS/CUPS/SINGLES|0.0|1|DONUT HOUSE DECAF K-CUPS|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|35.096297298232479|00099555089349|COFFEE|G1 GROCERY|-80.7007|80.700700114358924|147|1
35.06858|26779c787c58c9885aff60dbb925454e2333dfb5|5.99|2015-01-10 11:12:00|1.4091206135396188|1|9955508534|273|0.612062184999033|0|47|37|-80.7007|10|35.06858|PODS/CUPS/SINGLES|0.0|1|DONUT HOUSE DECAF K-CUPS|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00099555089349|COFFEE|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|e04d4c23b35a7686e2bb7507c3fdf7b03722d254|6.49|2015-01-31 10:55:00|1.4091206135396188|1|9955508534|273|0.612062184999033|0|47|37|-80.7007|10|35.06858|PODS/CUPS/SINGLES|0.0|1|DONUT HOUSE DECAF K-CUPS|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00099555089349|COFFEE|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|d4e29513b8a80ea6860d425e40d028f0c0472cc7|23.96|2014-12-13 11:08:00|1.4091206135396188|1|9955508534|273|0.612062184999033|0|47|37|-80.7007|10|35.06858|PODS/CUPS/SINGLES|0.0|1|DONUT HOUSE DECAF K-CUPS|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00099555089349|COFFEE|G1 GROCERY|-80.7007|1.4084929236641879|273|4
35.06858|127085a4056450029db1bd6f3c4208633444119a|5.97|2015-02-28 10:06:00|1.4091206135396188|1|2400016717|273|0.612062184999033|0|47|110|-80.7007|16|35.06858|FRUIT-CORE|0.97|1|DEL MONTE CHERRY MXD FRT LS.|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00024000019091|FRUIT-CAN/JAR|G1 GROCERY|-80.7007|1.4084929236641879|273|3
35.06858|67cc02c2753cead8d65c43b26155de56753761b8|5.19|2014-12-21 14:02:00|80.700248323638462|1|1980012738|273|35.101654671104228|0|7|724|-80.562829|69|35.006282|NFS-DRAIN CLEANER/OPENER|0.0|1|DRANO FOAMING LIQUID|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|35.096297298232479|00019800127381|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.7007|80.7007010071423|60|1
35.06858|fc7e472de6a983e415058a59efdff2e2bbe7a0d7|14.07|2014-11-20 17:29:00|1.4091206135396188|1|4900002468|273|0.612062184999033|0|47|55|-80.7007|8|35.06858|REGULAR|0.0|23|CLASSIC COKE .5 LITER/6 PK.|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00049000024685|CARBONATED BEVERAGES|BEVERAGE|-80.7007|1.4084929236641879|273|3
35.06858|3b94914333c67f8c696f9626546bc8766637df17|3.0|2014-11-30 20:27:00|1.4091206135396188|1|4023217761|273|0.612062184999033|0|47|8598|-80.7007|1792|35.06858|NEWSPAPERS|0.0|18|CHARLOTTE OBSERVER THANKGIVING|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00040232177613|NEWSPAPERS|GM|-80.7007|1.4084929236641879|273|1
35.06858|076ce2281c1dd48d4ecc9a693d3d3136c07bef65|1.79|2015-03-01 13:52:00|1.4091206135396188|1||273|0.612062184999033|0|47|540|-80.7007|64|35.06858|FRESH CELERY|0.0|4|COO CELERY (RPC) 24'S|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00204070000001|FRESH PRODUCE|PRODUCE|-80.7007|1.4084929236641879|273|1
35.06858|4718bd23434b492dbcc07fd9d86d72b00cd05b9e|6.98|2015-01-17 10:06:00|1.4091206135396188|1|20455000000|273|0.612062184999033|0|47|542|-80.7007|64|35.06858|FRESH VEGETABLES REMAIN|0.0|4|BRUSSEL SPROUTS 1LB (RPC)|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00094922577160|FRESH PRODUCE|PRODUCE|-80.7007|1.4084929236641879|273|2
35.06858|2734cf6d60bfc836a6c59207c60cb36903d66327|7.12|2014-11-01 11:01:00|1.4091206135396188|1|7740012733|273|0.612062184999033|0|47|838|-80.7007|102|35.06858|PEGS|0.0|19|CARL BUDDIG ORIGINAL HONEY HAM|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00077400128535|LUNCHMEATS|CASE READY MEATS|-80.7007|1.4084929236641879|273|8
35.06858|076cb97dc0cf826a4fabae0663f9d6674fb9ae08|7.12|2014-11-08 11:48:00|1.4091206135396188|1|7740012733|273|0.612062184999033|0|47|838|-80.7007|102|35.06858|PEGS|0.0|19|CARL BUDDIG ORIGINAL HONEY HAM|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00077400128535|LUNCHMEATS|CASE READY MEATS|-80.7007|1.4084929236641879|273|8
35.06858|1e8221a111a5c97219766a6fcd9b781bb88ad41c|4.59|2014-11-10 15:20:00|1.4091206135396188|1|2059300020|273|0.612062184999033|0|47|1459|-80.7007|40|35.06858|FROZEN BISCUITS|0.0|5|MARY B'S 20CT BUTRMILK BISCUIT|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00020593000201|FROZEN DOUGH|FROZEN|-80.7007|1.4084929236641879|273|1
35.06858|b6d181e36656187b77a200a2c01fa4f180e94127|2.89|2014-10-17 19:42:00|1.4091206135396188|1|7203697887|273|0.612062184999033|0|47|74|-80.7007|9|35.06858|RTE CEREAL ALL FAMILY|0.92|1|HT CER OATS & MORE HONEY|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036978875|CEREAL|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|bba82c168eadbd2f04570cb5a8a3da519d45d5a1|7.0|2014-10-31 15:23:00|1.4091206135396188|1|7203698425|273|0.612062184999033|0|47|254|-80.7007|892|35.06858|PREMIUM PIZZA|0.0|5|HT THIN CRUST PEPP/SAUS PIZZA|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036984265|FROZEN PIZZA|FROZEN|-80.7007|1.4084929236641879|273|2
35.06858|128c5c696c0fef4995fc2e53b0d02bbcfc982980|3.99|2014-11-01 19:17:00|1.4091206135396188|1|7203663995|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HARRIS TEETER 1% MILK|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036631275|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|d902d96ae9637061dede6cc0fe6d354a45a9f9b9|3.99|2014-10-21 18:51:00|1.4091206135396188|1|7203663995|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HARRIS TEETER 1% MILK|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036631275|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|050da14b5c588940b46da2eb1603d256806bbafd|3.99|2014-10-12 08:52:00|1.4091206135396188|1|7203663995|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|1.02|3|HARRIS TEETER 1% MILK|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036631275|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|742d5167e83ed83bb8d65cde52958bb18627e40b|3.49|2015-02-26 19:36:00|1.4091206135396188|1|7203663995|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HARRIS TEETER 1/2% MILK GALL|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036632012|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|d720d085b3cecfbe87aa40318e4a2447c2a5c14c|3.99|2014-09-25 17:00:00|1.4091206135396188|1|7203663995|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HARRIS TEETER 1% MILK|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036631275|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|d21009c3a786a5d9f8f78b81354aa37286328e7b|3.99|2014-12-09 18:55:00|1.4091206135396188|1|7203663995|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HARRIS TEETER 1% MILK|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036631275|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|fb64395244f60c366c9e3f13b9a11db5e7018fe3|11.97|2014-12-02 16:43:00|1.4091206135396188|1|7203663995|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|1.52|3|HARRIS TEETER 1% MILK|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036631275|MILK|DAIRY|-80.7007|1.4084929236641879|273|3
35.06858|00061d40b890c83260a0a5ed8fdae78a02b6b625|3.99|2014-09-13 10:14:00|1.4091206135396188|1|7203663995|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HARRIS TEETER 1% MILK|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036631275|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|141fe26c6f1e9ed102f84b909257885e5b0a1351|3.99|2014-11-14 19:37:00|1.4091206135396188|1|7203663995|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HARRIS TEETER 1% MILK|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036631275|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|b4edcbeab1eed2c16aef25461dc5f0688e67be68|3.99|2014-12-29 16:47:00|1.4091206135396188|1|7203663995|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HARRIS TEETER 1% MILK|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036631275|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|92db944d6447e68232ff2163ce62f5e705940d85|3.99|2014-11-20 07:45:00|1.4091206135396188|1|7203663995|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HARRIS TEETER 1% MILK|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036631275|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|81d02d24dcdcbbc93687c325ce4d80e60709ffcc|3.99|2014-09-28 17:36:00|1.4091206135396188|1|7203663995|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HARRIS TEETER 1% MILK|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036631275|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|9a2d9842baeddccf30457c43286164597187a6d1|3.49|2015-03-05 19:30:00|1.4091206135396188|1|7203663995|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HARRIS TEETER 1/2% MILK GALL|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036632012|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|e0312fc6ebd8394cb175b89f1eb0f90d22697128|3.99|2014-10-28 09:17:00|1.4091206135396188|1|7203663995|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HARRIS TEETER 1% MILK|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036631275|MILK|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|229a866c1f2fa82461ab8799cbb976105c8cfa94|3.99|2014-12-21 16:31:00|80.700248323638462|1|7203663995|273|35.101654671114375|0|7|342|-80.732725|57|35.082768|FRESH MILK|0.0|3|HARRIS TEETER 1% MILK|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|35.096297298232479|00072036631275|MILK|DAIRY|-80.7007|80.700700114358924|147|1
35.06858|452606350279c0b2ad668f984701fa14202b57c8|3.33|2015-02-28 22:21:00|1.4091206135396188|1|7203643010|273|0.612062184999033|0|47|252|-80.7007|45|35.06858|PREMIUM ICE CREAM|0.33|5|HT PREM PEANUT BUTTER CUP IC|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036430250|ICE CREAM|FROZEN|-80.7007|1.4084929236641879|273|1
35.06858|591c49742d7f94aad31538f4eb14c6e668a8d104|2.69|2014-12-07 14:08:00|1.4091206135396188|1|7294570544|273|0.612062184999033|0|47|1025|-80.7007|162|35.06858|WHITE|0.2|7|SL S&S  W.G. WHITE BREAD|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072945705449|SLICED BREAD|COMMERCIAL BAKERY|-80.7007|1.4084929236641879|273|1
35.06858|4bdfe28315823a9bdb8e71343860ae91da3f3e0b|2.19|2014-11-15 17:37:00|1.4091206135396188|1|1330018301|273|0.612062184999033|0|47|100|-80.7007|15|35.06858|CORN MEAL|0.0|1|MW BTTRMILK CORN MEAL MIX SR|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00013300183014|FLOUR|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|d589c96a5d165d27d71c71eb99f101228c3d644b|2.19|2014-10-17 17:38:00|1.4091206135396188|1|1330018301|273|0.612062184999033|0|47|100|-80.7007|15|35.06858|CORN MEAL|0.0|1|MW BTTRMILK CORN MEAL MIX SR|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00013300183014|FLOUR|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|69bd0f92fc831eee8b931ed75d2b2ec649b1b86d|7.78|2014-12-01 17:49:00|80.700248323638462|1|3700081114|273|35.101654671114375|0|7|4181|-80.732725|1085|35.082768|MISC TRIAL SIZE ITEM|0.9|17|(FE) FEBREEZE CAR CHECKSTAND|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|35.096297298232479|00037000865889|TRIAL SIZE|HBC|-80.7007|80.700700114358924|147|2
35.06858|688f9dd97b75dec7bfde079d6169729711d85b61|5.97|2015-02-16 17:18:00|1.4091206135396188|1|7203697992|273|0.612062184999033|0|47|273|-80.7007|43|35.06858|PREMIUM NOVELTIES|0.0|5|HT ICE CREAM SANDWICH-24PK|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036979926|FROZEN NOVELTIES|FROZEN|-80.7007|1.4084929236641879|273|1
35.06858|bfe3abc9da6d6e89b64790bb57f284cc36533015|2.99|2014-09-19 17:51:00|1.4091206135396188|1|7203608990|273|0.612062184999033|0|47|82|-80.7007|11|35.06858|VINEGAR|0.0|1|HT VINEGAR BALSAMIC|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036089908|CONDIMENTS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|8f64a1a659fdd17081647c622143bb67d422bde9|4.29|2015-01-31 15:02:00|1.4091206135396188|1|4178000011|273|0.612062184999033|0|47|201|-80.7007|31|35.06858|POTATO CHIPS|2.14|1|UTZ RIPPLE POTATO CHIPS|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00041780000910|SNACKS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|08b8e0cf9162e85d7b119a649de17ea8d8eba1fa|3.0|2014-09-14 13:58:00|1.4091206135396188|1||273|0.612062184999033|0|47|531|-80.7007|64|35.06858|FRESH CORN|0.2|4|COO YELLOW CORN|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00204078000003|FRESH PRODUCE|PRODUCE|-80.7007|1.4084929236641879|273|5
35.06858|fa9b1dbb647c5b99d7552d99649bea5ab3ef669f|6.3|2014-10-22 18:45:00|1.4091206135396188|1|7105200009|273|0.612062184999033|0|47|1461|-80.7007|40|35.06858|FROZEN GARLIC TOAST AND BRD|1.57|5|COLE'S GARLIC TOAST|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00071052000478|FROZEN DOUGH|FROZEN|-80.7007|1.4084929236641879|273|2
35.06858|3f36fb5d11d486ba046c14009f7ee5162a70473b|3.49|2014-10-19 17:25:00|1.4091206135396188|1|664|273|0.612062184999033|0|47|1639|-80.7007|377|35.06858|BULK (DONUTS)|0.0|14|PICK 6  DONUTS|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00000000006640|DONUTS|BAKERY|-80.7007|1.4084929236641879|273|1
35.06858|0d1a26e522f37a4c133202b339f08f8c6c93acc5|3.49|2015-02-19 17:41:00|1.4091206135396188|1|664|273|0.612062184999033|0|47|1639|-80.7007|377|35.06858|BULK (DONUTS)|0.0|14|PICK 6  DONUTS|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00000000006640|DONUTS|BAKERY|-80.7007|1.4084929236641879|273|1
35.06858|91c4f042d50eee485d0df763ab23042d3a445aeb|3.49|2015-01-04 09:09:00|1.4091206135396188|1|664|273|0.612062184999033|0|47|1639|-80.7007|377|35.06858|BULK (DONUTS)|0.0|14|PICK 6  DONUTS|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00000000006640|DONUTS|BAKERY|-80.7007|1.4084929236641879|273|1
35.06858|31913296361ec13d95230e4d10abefac6ce87004|3.99|2015-02-25 19:14:00|1.4091206135396188|1|7203688076|273|0.612062184999033|0|47|523|-80.7007|64|35.06858|FRESH POTATOES|0.99|4|HT RUSSET POTATO 5LB BAG|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036880765|FRESH PRODUCE|PRODUCE|-80.7007|1.4084929236641879|273|1
35.06858|a4eecc6c94e2dd0c611d6b07f63f8242eb7a7bdf|3.49|2014-10-30 15:19:00|1.4091206135396188|1|7203659049|273|0.612062184999033|0|47|313|-80.7007|51|35.06858|MARGARINE|0.5|3|HT MARGARINE SPREAD|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036590497|BUTTER & MARGARINE|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|a84ef51156c392d33ac69951126a9ae91956a9b1|3.49|2015-02-06 12:15:00|1.4091206135396188|1|7203659049|273|0.612062184999033|0|47|313|-80.7007|51|35.06858|MARGARINE|0.5|3|HT MARGARINE SPREAD|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036590497|BUTTER & MARGARINE|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|1560fe08088d695ff1b39a7ab26a421049098ef9|3.49|2014-12-11 16:41:00|1.4091206135396188|1|7203659049|273|0.612062184999033|0|47|313|-80.7007|51|35.06858|MARGARINE|0.5|3|HT MARGARINE SPREAD|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036590497|BUTTER & MARGARINE|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|8b6257ecc1bcf525a23441320fbc963c0df6d99a|3.97|2015-02-22 17:51:00|1.4091206135396188|1|7203663053|273|0.612062184999033|0|47|335|-80.7007|56|35.06858|ORANGE JUICE-REGRIGERATED|0.0|3|HT ORANGE JUICE GALLON|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036630537|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|99ac816ad0b2019afcbdf3c23af144e344b4effa|3.79|2014-10-26 12:35:00|1.4091206135396188|1|2500005542|273|0.612062184999033|0|47|335|-80.7007|56|35.06858|ORANGE JUICE-REGRIGERATED|0.79|3|SIMPLY ORANGE GROVE MADE|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00025000055447|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|b3c9c047f78ee866decbc384ecad8d45649d2c15|3.96|2014-10-13 17:28:00|1.4091206135396188|1|3400000031|273|0.612062184999033|0|47|47|-80.7007|7|35.06858|REGISTER BARS|0.5|1|HEATH BAR ORIGINAL|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00010700060808|CANDY|G1 GROCERY|-80.7007|1.4084929236641879|273|4
35.06858|253bf6dfc72aa7c49626269df08a51db15d8a404|3.69|2014-12-28 13:41:00|1.4091206135396188|1|61144334026|273|0.612062184999033|0|47|214|-80.7007|33|35.06858|BROTH|0.9|1|KITCHEN BASICS STOCK VEGETABLE|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00611443340211|SOUP|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|cc2104d48538db14ddaddb31c54535011723fcbd|1.94|2015-03-01 16:08:00|1.4091206135396188|1|7203637031|273|0.612062184999033|0|47|212|-80.7007|33|35.06858|CONDENSED SOUP|0.0|1|HT SP RS CRM MUSHROOM|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036978547|SOUP|G1 GROCERY|-80.7007|1.4084929236641879|273|2
35.06858|a9bfde5c25afacfe396965b36ace99fc93aee3c0|0.97|2015-03-03 17:18:00|1.4091206135396188|1|7203637031|273|0.612062184999033|0|47|212|-80.7007|33|35.06858|CONDENSED SOUP|0.0|1|HT SP RS CRM MUSHROOM|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036978547|SOUP|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|05a8760029f6f21844a9a874cfa1b22c9ad6a605|3.79|2014-12-22 10:52:00|1.4091206135396188|1|4850002013|273|0.612062184999033|0|47|335|-80.7007|56|35.06858|ORANGE JUICE-REGRIGERATED|0.79|3|TROPICANA PP GROVESTAND|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00048500304143|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|f0d0aa22414d360d5a9f65b08665ccc74c6e875c|1.49|2014-12-12 18:41:00|1.4091206135396188|1|20406100000|273|0.612062184999033|0|47|525|-80.7007|64|35.06858|FRESH LETTUCE|0.0|4|ICEBERG LETTUCE|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00033383650203|FRESH PRODUCE|PRODUCE|-80.7007|1.4084929236641879|273|1
35.06858|471ea9080809ca2decc7eee699ec03ca4e999878|12.77|2015-03-08 17:07:00|1.4091206135396188|1|20319700000|273|0.612062184999033|0|47|641|-80.7007|137|35.06858|PREMIUM PORK|6.58|2|VALUE PK PORK BUTT CNTRY RIB|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00203197000000|PORK|MEAT|-80.7007|1.4084929236641879|273|1
35.06858|e04bb2de218aa98388e0c15418132d3c6ac73ba1|5.49|2015-01-24 18:50:00|1.4091206135396188|1|4400003327|273|0.612062184999033|0|47|1248|-80.7007|12|35.06858|SANDWICH COOKIES|1.0|1|OREO FAMILY SIZED|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00044000033279|COOKIES|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|524f2d00257cd0ed694f0fa1c61db37a0b8e05f3|8.58|2014-12-31 15:40:00|1.4091206135396188|1|2840016014|273|0.612062184999033|0|47|201|-80.7007|31|35.06858|POTATO CHIPS|2.14|1|LAYS BBQ|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00028400160131|SNACKS|G1 GROCERY|-80.7007|1.4084929236641879|273|2
35.06858|6be74116eb23a8224edef2402ec611b26389d872|1.77|2015-01-25 10:26:00|1.4091206135396188|1|7203639031|273|0.612062184999033|0|47|228|-80.7007|36|35.06858|TABLE SYRUP|0.1|1|HT LITE BUTTER FLAVORED SYRUP|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036390349|TABLE SYRUPS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|558df7d629cd4a707f210b9e5ce30e298ec4988a|1.17|2014-10-18 17:09:00|1.4091206135396188|1|7294012570|273|0.612062184999033|0|47|70|-80.7007|11|35.06858|KETCHUP|0.0|1|VINE RIPE KETCHUP 24|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072940125709|CONDIMENTS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|2b6112988632f3fb3537c0fcc953319e58a12e17|2.19|2014-09-18 09:07:00|1.4091206135396188|1|84981900002|273|0.612062184999033|0|47|55|-80.7007|8|35.06858|REGULAR|1.2|23|NATURES TWIST LEMONADE 2L|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00849819000029|CARBONATED BEVERAGES|BEVERAGE|-80.7007|1.4084929236641879|273|1
35.06858|e5f20c56efac69f8ed17b926f35214998a81fbf3|2.19|2014-10-29 20:00:00|1.4091206135396188|1|4900005010|273|0.612062184999033|0|47|55|-80.7007|8|35.06858|REGULAR|0.2|23|CLASSIC COKE 2 LT CONTOUR|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00049000050103|CARBONATED BEVERAGES|BEVERAGE|-80.7007|1.4084929236641879|273|1
35.06858|6103d58b91e81702e674e02f4ccd1c7dfad8d2d8|2.69|2015-02-04 20:26:00|1.4091206135396188|1|3000016900|273|0.612062184999033|0|47|721|-80.7007|31|35.06858|RICE SNACKS|0.0|1|QUAKER OATS CARAMEL CORN CAKES|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00030000169100|SNACKS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|f42dc007385c52843f6e21ed8599b0217c90f62d|13.99|2014-09-26 14:47:00|1.4091206135396188|1|1820014990|273|0.612062184999033|0|47|461|-80.7007|84|35.06858|FLAVORED MALT BEVERAGE|0.0|16|BUD LIGHT LIME 12PK LNNR|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00018200149900|SPECIALTY|BEER|-80.7007|1.4084929236641879|273|1
35.06858|cd40591ea0b38664521fa56f709c071ac0669786|13.99|2014-12-20 17:46:00|1.4091206135396188|1|1820014990|273|0.612062184999033|0|47|461|-80.7007|84|35.06858|FLAVORED MALT BEVERAGE|0.0|16|BUD LIGHT LIME 12PK LNNR|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00018200149900|SPECIALTY|BEER|-80.7007|1.4084929236641879|273|1
35.06858|ab02ace257651d8973f251d445d195aa8121909c|5.98|2015-01-17 14:12:00|1.4091206135396188|1|7433610102|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HIGHLAND CREST 2% REDUCE FAT|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00074336101021|MILK|DAIRY|-80.7007|1.4084929236641879|273|2
35.06858|234a739bac57b33ab8e8b0d91156f47e011126a5|5.98|2015-01-11 18:36:00|1.4091206135396188|1|7433610102|273|0.612062184999033|0|47|342|-80.7007|57|35.06858|FRESH MILK|0.0|3|HIGHLAND CREST 2% REDUCE FAT|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00074336101021|MILK|DAIRY|-80.7007|1.4084929236641879|273|2
35.06858|cccd7fe8fb3b9860f9a39410ef4019cc15a09784|1.17|2014-10-03 14:34:00|1.4091206135396188|1|7203690020|273|0.612062184999033|0|47|1034|-80.7007|163|35.06858|HOT DOG|0.2|7|H T HOT DOG BUNS|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036900203|BUNS/ROLLS|COMMERCIAL BAKERY|-80.7007|1.4084929236641879|273|1
35.06858|dfafba13692854e26f09e53233b3e0efc6317743|1.94|2014-10-08 19:53:00|1.4091206135396188|1|7203690010|273|0.612062184999033|0|47|1025|-80.7007|162|35.06858|WHITE|0.0|7|H T SANDWICH BREAD|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036900104|SLICED BREAD|COMMERCIAL BAKERY|-80.7007|1.4084929236641879|273|2
35.06858|17c3d1a686f38cb04481117cee36d1cd71a1889c|1.17|2014-10-22 12:44:00|1.4091206135396188|1|7203690020|273|0.612062184999033|0|47|1034|-80.7007|163|35.06858|HOT DOG|0.0|7|H T HOT DOG BUNS|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036900203|BUNS/ROLLS|COMMERCIAL BAKERY|-80.7007|1.4084929236641879|273|1
35.06858|315cfb5a7c62cb2207167175448ca0167847bac2|1.94|2014-12-27 19:04:00|1.4091206135396188|1|7203690010|273|0.612062184999033|0|47|1025|-80.7007|162|35.06858|WHITE|0.0|7|H T SANDWICH BREAD|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036900104|SLICED BREAD|COMMERCIAL BAKERY|-80.7007|1.4084929236641879|273|2
35.06858|4afa6336f09dc6a810f8b3b6fe607a66b0105273|3.98|2014-10-11 16:42:00|1.4091206135396188|1|7203671215|273|0.612062184999033|0|47|225|-80.7007|35|35.06858|SUGAR-GRANULATED|0.0|1|HT GRANULATED SUGAR|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036712158|SUGAR/SUBSTITUTES|G1 GROCERY|-80.7007|1.4084929236641879|273|2
35.06858|6750a1b1c3c8af10a3f3f94539114e7df058ba93|2.29|2015-01-07 15:19:00|1.4091206135396188|1|1800000260|273|0.612062184999033|0|47|325|-80.7007|54|35.06858|BISCUITS-REFRIGERATED|1.29|3|GRANDS BUTTERMILK BISCUITS|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00018000001828|DOUGH PRODUCTS|DAIRY|-80.7007|1.4084929236641879|273|1
35.06858|91fa2f3fc19e127e959df5d6538f7642b819e428|2.5|2014-09-29 16:40:00|1.4091206135396188|1|7203697755|273|0.612062184999033|0|47|81|-80.7007|9|35.06858|RTE CEREAL KIDS|0.53|1|HT CER FRUIT O'S|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036979919|CEREAL|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|271c8d26e6ddab263c5a0455b58782e38607ccbf|10.0|2014-12-13 09:59:00|1.4091206135396188|1|7203697755|273|0.612062184999033|0|47|81|-80.7007|9|35.06858|RTE CEREAL KIDS|2.12|1|HT CER FRUIT O'S|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036979919|CEREAL|G1 GROCERY|-80.7007|1.4084929236641879|273|4
35.06858|7212d904567161810812b7389da61c3214679e32|2.5|2015-02-14 20:27:00|1.4091206135396188|1|7203697755|273|0.612062184999033|0|47|81|-80.7007|9|35.06858|RTE CEREAL KIDS|0.53|1|HT CER FRUIT O'S|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036979919|CEREAL|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|f1cb052adc5de47e315055847eb9c28b2ca0f9c0|1.87|2014-11-30 14:55:00|1.4091206135396188|1|7203642061|273|0.612062184999033|0|47|236|-80.7007|38|35.06858|DRY BEANS|0.0|1|HT BEANS DRY PINTO 32|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036420619|RICE GRAINS AND BEANS|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|5488fbf4c61d04fc13bb1d7787deec711e0727e5|2.37|2015-03-09 19:34:00|1.4091206135396188|1|7203632024|273|0.612062184999033|0|47|195|-80.7007|30|35.06858|SALAD & COOKING OIL|0.0|1|HT CORN OIL|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00072036320247|SHORTENING/OIL|G1 GROCERY|-80.7007|1.4084929236641879|273|1
35.06858|f274bbde78d11c22fbb382a429e80fbb7fe483f0|3.94|2014-10-20 12:04:00|1.4091206135396188|1|5420004053|273|0.612062184999033|0|47|416|-80.7007|71|35.06858|NFS-BLEACH|0.0|1|101 REGULAR BLEACH|74a263b33df2b570128af55aac4be269997e9efe|2.2853799015412375|0.61242566243833529|00054200040533|LAUNDRY SUPPLIES|G1 GROCERY|-80.7007|1.4084929236641879|273|2
35.28326|9c6e8c0de4f4a8dc8fe75d61c0b363eec0723d35|1.99|2014-11-09 11:17:00|1.4094857484078087|1|5100017520|46|0.6158090578372145|0|26|1201|-80.66939|33|35.28326|RTS CANNED|0.49|1|CAM HOMESTYLE CREOLE CHICKEN|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00051000195647|SOUP|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|9080a2ba3f7a8f07fbbef5d0f9cd12b73fdf597a|3.98|2015-01-03 12:50:00|1.4094857484078087|1|5100000524|46|0.6158090578372145|0|26|1201|-80.66939|33|35.28326|RTS CANNED|0.98|1|CHUNKY HR SIRLOIN BURGER|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00051000180346|SOUP|G1 GROCERY|-80.66939|1.4079464610753885|46|2
35.28326|fcf591e0da64f49df73a8b2584693ea520efddec|4.58|2014-10-05 19:39:00|1.4094857484078087|1|5100000524|46|0.6158090578372145|0|26|1201|-80.66939|33|35.28326|RTS CANNED|1.58|1|CHUNKY HR SIRLOIN BURGER|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00051000180346|SOUP|G1 GROCERY|-80.66939|1.4079464610753885|46|2
35.28326|604f00e69993c3352b666bf0f7d23cbda6ebca36|6.79|2014-11-16 11:38:00|1.4094857484078087|1|4900002890|46|0.6158090578372145|0|26|54|-80.66939|8|35.28326|DIET|6.79|23|DT SPRITE ZERO 12PK FRIDGEPKCN|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00049000037111|CARBONATED BEVERAGES|BEVERAGE|-80.66939|1.4079464610753885|46|1
35.28326|4f1b3f97fef840eef224a280000f7aedbfd80d05|2.89|2015-03-08 09:19:00|1.4094857484078087|1|3760007060|46|0.6158090578372145|0|26|714|-80.66939|274|35.28326|MICROWAVE MEALS|0.39|1|HORMEL CMPL TURKEY DRESSING|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00037600369183|PREP FOODS DINNERS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|009f5685dc30fb51a1479abfa18d585954d2bf2b|2.89|2015-01-06 18:05:00|1.4094857484078087|1|3760007060|46|0.6158090578372145|0|26|714|-80.66939|274|35.28326|MICROWAVE MEALS|0.39|1|HORMEL CMPL TURKEY DRESSING|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00037600369183|PREP FOODS DINNERS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|e9f30f6c647fd18dbe236014eb345a37f8723c9e|2.29|2014-10-15 17:46:00|1.4094857484078087|1|7357013000|46|0.6158090578372145|0|26|1267|-80.66939|53|35.28326|DIPS AND SPREADS|0.79|3|HELUVA GOOD FRENCH ONION DIP|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00073570130002|CULTURES|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|1905a30bb932f9d2137662a12b22204295adee4e|2.58|2014-11-28 09:50:00|1.4094857484078087|1|7205861029|46|0.6158090578372145|0|26|1147|-80.66939|229|35.28326|HOT COCOA MIX|1.2|1|I/O LD O LK CAPP AMARETTO|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00072058610289|COCOAS CREAMERS SYRUPS|G1 GROCERY|-80.66939|1.4079464610753885|46|2
35.28326|a0dd47b083526ba29f249817c1c018727d42387a|5.49|2014-10-19 18:22:00|1.4094857484078087|1|7403006610|46|0.6158090578372145|0|26|332|-80.66939|52|35.28326|STRING/SNACK|2.49|3|SORRENTO CHEDDAR STICKSTERS|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00074030069207|CHEESE|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|aabf1376f05613e19d002150c0ca4e807b4bc785|3.59|2014-12-22 19:10:00|1.4094857484078087|1|4150022020|46|0.6158090578372145|0|26|164|-80.66939|39|35.28326|VEGETABLES-SPECIALTY|0.6|1|FRENCHS FRIED ONION 6 OZ|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00041500220208|VEGETABLES-CAN/JAR|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|11ec9c8c3a3957c6afd8fc6d8b62f9fa794196af|3.39|2015-01-12 18:19:00|1.4094857484078087|1|2100012382|46|0.6158090578372145|0|26|320|-80.66939|53|35.28326|COTTAGE CHEESE|0.89|3|BREAKSTONE 2% L/F COTTAGE CHS|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00021000123827|CULTURES|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|c36f3614196d8a4bf6b99e121a790ff68ad0a7e7|3.39|2015-03-07 21:01:00|1.4094857484078087|1|2100012382|46|0.6158090578372145|0|26|320|-80.66939|53|35.28326|COTTAGE CHEESE|0.89|3|BREAKSTONE 2% L/F COTTAGE CHS|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00021000123827|CULTURES|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|ce0003959089d3962e3093554feff8a4de8c4179|11.99|2014-12-20 13:17:00|1.4094857484078087|1|3700088206|46|0.6158090578372145|0|26|426|-80.66939|72|35.28326|NFS-PAPER TOWELS|2.0|1|BOUNTY TOWEL 6 RL WHITE|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00037000882060|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|d734dc59a877a65141664e574dbed747dbd92e11|3.89|2014-11-25 13:49:00|80.669414401537693|1|3700042728|46|35.302041710208115|0|19|4074|-80.737839|1080|35.297134|TOOTHPASTE-CHILD|0.9|17|CREST NEAT SQZ KID|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|35.305725790410776|00037000003380|ORAL HYGIENE|HBC|-80.66939|80.669393843943624|258|1
35.28326|f5619f7356e745604c65ce14f877aef3312671bd|2.19|2015-01-18 14:49:00|80.669414401537693|1|3760003895|46|35.302041710208115|0|19|659|-80.737839|103|35.297134|CHILDRENS LUNCH SNACKS|0.19|19|HORMEL REV ITALIAN WRAP|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|35.305725790410776|00037600676076|LUNCH SNACKS|CASE READY MEATS|-80.66939|80.669393843943624|258|1
35.28326|2272966152b5067bec66cb51d10fabce147e6f7e|1.57|2014-11-25 13:53:00|80.669414401537693|1|7009030410|46|35.302041710208115|0|19|225|-80.737839|35|35.297134|SUGAR-GRANULATED|0.0|1|CRYSTAL FINE GRANULATED SUGAR|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|35.305725790410776|00070090304104|SUGAR/SUBSTITUTES|G1 GROCERY|-80.66939|80.669393843943624|258|1
35.28326|0eaf6d461bff34cd79d413e638eb468d35018abd|3.39|2015-02-09 18:52:00|1.4094857484078087|1|5100020472|46|0.6158090578372145|0|26|1261|-80.66939|274|35.28326|MEAL STARTERS|0.0|1|CAMP SLOWCOOK TAVERN POT ROAST|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00051000204721|PREP FOODS DINNERS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|b5eb42cf4248034905ea76b6f646bfaa78bec794|6.99|2014-10-18 11:33:00|1.4094857484078087|1|7116967062|46|0.6158090578372145|0|26|7248|-80.66939|1600|35.28326|HALLOWEEN ACCESSORIES IMP|1.0|18|PUMPKIN CARVING KIT|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00071169670625|SEASONAL MERCHANDISE|GM|-80.66939|1.4079464610753885|46|1
35.28326|a23880b980034536ac05b450ce59e2480922bd91|7.54|2014-12-13 11:21:00|1.4094857484078087|1|7203603040|46|0.6158090578372145|0|26|217|-80.66939|34|35.28326|EXTRACTS FOOD COLORING|0.0|1|HT VANILLA EXTRACT|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00072036030405|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.66939|1.4079464610753885|46|2
35.28326|bbc59e1ebe5254dfe6bfa58b707cdef857d78b8d|13.99|2014-10-10 17:06:00|80.669414401537693|1|9256710537|46|35.302041678522976|0|19|6790|-80.605588|1568|35.43259|MAGAZINES SEMI ANNUAL|0.0|18|LIFE SPECIAL|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|35.305725790410776|00092567105373|MAGAZINES|GM|-80.66939|80.669432442000655|202|1
35.28326|3957c803e29d27e3016646fdc6bbb27fdbb6f39b|3.59|2015-01-24 13:41:00|1.4094857484078087|1|4116400022|46|0.6158090578372145|0|26|1469|-80.66939|278|35.28326|REGULAR CUT FRIES|0.59|5|MRS T'S POTATO CHDR PIEROGIES|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00041164000222|FROZEN POTATO|FROZEN|-80.66939|1.4079464610753885|46|1
35.28326|2b8dc7cee0039c130828fead92724c9d00b17209|3.79|2014-10-19 10:47:00|1.4094857484078087|1|4470000857|46|0.6158090578372145|0|26|839|-80.66939|102|35.28326|STACK PACKS|0.0|19|OSCAR MAYER BOLOGNA|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00044700008577|LUNCHMEATS|CASE READY MEATS|-80.66939|1.4079464610753885|46|1
35.28326|290c92e37c3f66673dc0d134a86a7237b6a05a5a|24.99|2015-02-07 16:44:00|1.4094857484078087|1|72760005980|46|0.6158090578372145|0|26|1509|-80.66939|87|35.28326|FLOR-FLORAL-CANDY ARANGEMENT|0.0|9|MIXED CHOCOLATE VASE  VALENTIN|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00727600059800|FLORAL|FLORAL|-80.66939|1.4079464610753885|46|1
35.28326|476f9a09ad1a962f526099391b1ac8e6b46b4b7e|10.96|2015-02-01 13:05:00|1.4094857484078087|1||46|0.6158090578372145|0|26|503|-80.66939|64|35.28326|FRESH GRAPES|1.57|4|RED GRAPES,SEEDLESS 12/16|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00204023000003|FRESH PRODUCE|PRODUCE|-80.66939|1.4079464610753885|46|1
35.28326|715ffe79af8a7ed39b6d1b31d578c244a27cadc1|2.19|2014-10-11 16:12:00|80.669414401537693|1|7203656071|46|35.302041710208115|0|19|316|-80.737839|52|35.297134|CREAM CHEESE|0.0|3|HT HONEY NUT SOFT CREAM CHEESE|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|35.305725790410776|00072036600837|CHEESE|DAIRY|-80.66939|80.669393843943624|258|1
35.28326|9c21c9d4fd58746e567cf7be7cc57488a6ad6e14|4.89|2014-12-26 14:53:00|1.4094857484078087|1|1600048366|46|0.6158090578372145|0|26|74|-80.66939|9|35.28326|RTE CEREAL ALL FAMILY|0.0|1|GM CHEERIOS HONEY NUT 21.6|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00016000483668|CEREAL|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|21787d9ae5ddd8209b6cec33b827f4a6f147dc24|2.69|2014-09-23 17:24:00|80.669414401537693|1|7203663996|46|35.302041710208115|0|19|342|-80.737839|57|35.297134|FRESH MILK|0.0|3|HARRIS TEETER 2%   MILK|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|35.305725790410776|00072036639998|MILK|DAIRY|-80.66939|80.669393843943624|258|1
35.28326|9430f0658ba388db4c83911ee552f40b51d93e1b|4.29|2014-09-26 19:07:00|80.669414401537693|1|2840015636|46|35.302041678522976|0|19|204|-80.605588|31|35.43259|TORTILLA CHIPS|2.15|1|DORTIOS NACHO CHEESE|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|35.305725790410776|00028400156363|SNACKS|G1 GROCERY|-80.66939|80.669432442000655|202|1
35.28326|6e4cdb1326252965368286b254d3b9d05a12711a|2.3|2014-12-31 16:17:00|80.669414401537693|1|2700050006|46|35.302041710208115|0|19|1221|-80.737839|275|35.297134|PASTA SC VALUE|0.0|1|HUNTS SC SPAG GARLIC HERB|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|35.305725790410776|00027000500118|PASTA SAUCES|G1 GROCERY|-80.66939|80.669393843943624|258|2
35.28326|277861b1f62a14399e9378845dad533a6f5dee8d|1.15|2015-02-18 13:07:00|80.669414401537693|1|2700050006|46|35.302041694565766|0|19|1221|-80.810056|275|35.219587|PASTA SC VALUE|0.15|1|HUNTS SC SPAG GARLIC HERB|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|35.305725790410776|00027000500118|PASTA SAUCES|G1 GROCERY|-80.66939|80.669419945960428|401|1
35.28326|20d5e1cb6546ad6e668a1e44db2d4cdbc1a9779b|3.65|2014-11-24 12:07:00|80.669414401537693|1|3010067264|46|35.302041710208115|0|19|91|-80.737839|13|35.297134|SPRAYED BUTTER CRACKERS|1.15|1|TOWN HOUSE PRETZEL THINS PARMS|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|35.305725790410776|00030100102335|CRACKERS|G1 GROCERY|-80.66939|80.669393843943624|258|1
35.28326|f32db38c24c89d4ad3ed7a6b394ab825d6303710|0.72|2014-09-21 10:17:00|1.4094857484078087|1||46|0.6158090578372145|0|26|502|-80.66939|64|35.28326|FRESH BANANAS|0.0|4|BANANAS, YELLOW|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00204011000008|FRESH PRODUCE|PRODUCE|-80.66939|1.4079464610753885|46|1
35.28326|acf2fe149f5635768a1cde29c25704ac336eabd4|3.99|2015-02-12 17:07:00|1.4094857484078087|1|3760039885|46|0.6158090578372145|0|26|362|-80.66939|102|35.28326|PEPPERONIS|0.0|19|HORMEL PEPPERONI MINIS|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00037600591829|LUNCHMEATS|CASE READY MEATS|-80.66939|1.4079464610753885|46|1
35.28326|13f1fff5f24c9d4e980b2159ff9a7dca37b3d339|3.35|2014-09-22 17:34:00|1.4094857484078087|1|7203656080|46|0.6158090578372145|0|26|318|-80.66939|52|35.28326|SHREDDED/GRATED CHEESE|1.35|3|HT FANCY SHRED SHARP CHED CHE|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00072036550262|CHEESE|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|bfbd23d7f079d741881281b3b79e55f26624c6f4|1.79|2015-02-15 08:11:00|1.4094857484078087|1|1800000261|46|0.6158090578372145|0|26|325|-80.66939|54|35.28326|BISCUITS-REFRIGERATED|0.29|3|GRANDS FLAKY BISCUITS|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00018000002610|DOUGH PRODUCTS|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|fc990d618dd62b547dc95fb7cea5d312378fe6a9|11.16|2014-11-28 13:36:00|1.4094857484078087|1|7203698417|46|0.6158090578372145|0|26|423|-80.66939|72|35.28326|NFS-DISPOSE PLATES/BOWLS|1.16|1|YH ELEGWARE BOWL 20 OZ|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00072036984180|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.66939|1.4079464610753885|46|4
35.28326|2cec69f64db69f83f25b5cf52083d01361398fb5|5.98|2014-10-25 09:48:00|1.4094857484078087|1|8186422116|46|0.6158090578372145|0|26|583|-80.66939|136|35.28326|NUTS|0.98|4|SALTED PEANUTS IN-SHELL|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00081864221169|OTHER MERCHANDISE|PRODUCE|-80.66939|1.4079464610753885|46|2
35.28326|c9ba0e5ce75207d1c501c7ee2c2e316822a0f912|19.99|2014-09-14 18:30:00|80.669414401537693|1|8281597780|46|35.302041678522976|0|19|6851|-80.605588|1578|35.43259|UMBRELLAS|0.0|18|"62"" DBL CANOPY GOLF UMBRELLA"|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|35.305725790410776|00082815977807|UMBRELLAS|GM|-80.66939|80.669432442000655|202|1
35.28326|20837ae9dd02e70191c930425734cc84bc13e295|1.77|2015-02-23 16:40:00|1.4094857484078087|1|7203657031|46|0.6158090578372145|0|26|322|-80.66939|53|35.28326|SOUR CREAM|0.0|3|HT SOUR CREAM|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00072036570314|CULTURES|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|38d87ead2d8d0f33a99af7c33a9ffadc16789d51|1.99|2014-11-08 17:02:00|1.4094857484078087|1|7127915101|46|0.6158090578372145|0|26|555|-80.66939|64|35.28326|PACKAGED SALADS|0.0|4|F.E. SHREDS|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00071279151014|FRESH PRODUCE|PRODUCE|-80.66939|1.4079464610753885|46|1
35.28326|8e6d3a8c34c8c6f65a95028e9e31aeffae3662d5|3.99|2015-01-17 17:28:00|1.4094857484078087|1|5929057322|46|0.6158090578372145|0|26|92|-80.66939|13|35.28326|REMAINING CRACKERS|0.99|1|CARRS CRACK PEPPER TABLE CRACK|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00059290575927|CRACKERS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|7ededb4c27617350d2205e95866110c8bb96a414|12.99|2014-12-24 10:08:00|1.4094857484078087|1|8470409132|46|0.6158090578372145|0|26|9983|-80.66939|889|35.28326|NFS-SPARKLING|0.0|13|CB-KORBEL BRUT|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00084704091328|SPARKLING|WINE|-80.66939|1.4079464610753885|46|1
35.28326|888556d754ae390764174859931d239dbe6f0fa4|2.99|2015-02-25 21:25:00|80.669414401537693|1|67791671646|46|35.302041678522976|0|19|7002|-80.605588|1600|35.43259|VALENTINE PARTY GOOD/DECORTN|2.24|18|I/O 4PC GLITTER HEART CUTOUTS|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|35.305725790410776|00677916716464|SEASONAL MERCHANDISE|GM|-80.66939|80.669432442000655|202|1
35.28326|928fbe84814499f3e9fbe890c7bd8bdeb232661a|3.99|2015-02-22 16:52:00|1.4094857484078087|1|1520125907|46|0.6158090578372145|0|26|7071|-80.66939|1600|35.28326|EASTER EGGS/NOVELTIES|1.0|18|I/OKRAZY MASN JAR W/DAISY STRW|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00015201259072|SEASONAL MERCHANDISE|GM|-80.66939|1.4079464610753885|46|1
35.28326|099ac4b87c74e467050d857f50b07046e24999af|3.19|2014-10-30 16:35:00|80.669414401537693|1|82951530146|46|35.302041694001396|0|19|205|-80.70901|31|35.17335|REMAINING SNACKS|1.6|1|SENSBL PORT VEG CHIPS LT SALT|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|35.305725790410776|00829515301460|SNACKS|G1 GROCERY|-80.66939|80.669420472648255|174|1
35.28326|5871d798279d00ebe893adbe80e7ccb181915a5b|3.49|2014-12-29 17:41:00|1.4094857484078087|1|7080003720|46|0.6158090578372145|0|26|839|-80.66939|102|35.28326|STACK PACKS|0.0|19|SMITHFIELD CUBED HAM|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00070800037209|LUNCHMEATS|CASE READY MEATS|-80.66939|1.4079464610753885|46|1
35.28326|64735d3320dd1610ca15cd6a07cad72f12794df2|5.49|2014-11-07 13:01:00|80.669414401537693|1|7192196143|46|35.302041710208115|0|19|254|-80.737839|892|35.297134|PREMIUM PIZZA|1.5|5|DIGIORNO TC SPINACH & GARLC|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|35.305725790410776|00071921451431|FROZEN PIZZA|FROZEN|-80.66939|80.669393843943624|258|1
35.28326|09bb18d8ddb29f0562aa762afd502715e2e1655c|16.99|2014-09-27 15:29:00|1.4094857484078087|1|79837312125|46|0.6158090578372145|0|26|458|-80.66939|82|35.28326|CRAFT BEER|0.0|16|MAGIC HAT THIS & THAT 12PK|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00798373121254|DOMESTIC BEER|BEER|-80.66939|1.4079464610753885|46|1
35.28326|83279396826872ff0c59fe58d6ab8a46f7ac8400|10.09|2015-01-10 18:07:00|1.4094857484078087|1||46|0.6158090578372145|0|26|566|-80.66939|64|35.28326|SERVICE BAR|0.71|4|HT 7 LAYER MEXICAN BEAN DIP|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00204506000001|FRESH PRODUCE|PRODUCE|-80.66939|1.4079464610753885|46|2
35.28326|a8bd7601c2cd8ba1d9cdb0297c091ba3e72b9d7b|35.95|2014-12-31 17:58:00|80.669414401537693|1|7080004118|46|35.302041678522976|0|19|358|-80.605588|100|35.43259|REGULAR BACON|0.0|19|SMITHFIELD PREMIUM BACON|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|35.305725790410776|00070800041183|BACON|CASE READY MEATS|-80.66939|80.669432442000655|202|5
35.28326|b45255a3fe366100ade73d2f9ab266a0ebd103cd|3.49|2015-02-16 17:30:00|1.4094857484078087|1|4610000107|46|0.6158090578372145|0|26|331|-80.66939|52|35.28326|NATURAL SLICED|0.0|3|SARGENTO DELI STYLE PROVOLNE|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00046100001233|CHEESE|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|c5f0b796002a58236736c42e0712dbbb3c7aee78|3.99|2014-11-28 15:46:00|1.4094857484078087|1|7110021094|46|0.6158090578372145|0|26|182|-80.66939|28|35.28326|MAYO|0.0|1|D HVR SNDWICH SPREAD GARLIC PA|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00071100210958|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|5a113a0136519f4ea95d166cf391984a00876717|2.75|2014-11-02 13:47:00|1.4094857484078087|1|5100012573|46|0.6158090578372145|0|26|137|-80.66939|20|35.28326|TOMATO & VEGETABLE JUICE|0.25|1|V8 SPLASH APPLE MEDLEY|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00051000203465|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|b814982373051d26b955125dde6046e3e8985468|2.19|2014-10-18 17:59:00|80.669414401537693|1|7800008246|46|35.302041678522976|0|19|54|-80.605588|8|35.43259|DIET|0.2|23|DIET DR PEPPER 2 LITER|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|35.305725790410776|00078000083460|CARBONATED BEVERAGES|BEVERAGE|-80.66939|80.669432442000655|202|1
35.28326|3146b90ef844f939480b8de8096a8b1a7077ad45|1.99|2014-11-01 12:23:00|1.4094857484078087|1|7130904547|46|0.6158090578372145|0|26|1025|-80.66939|162|35.28326|WHITE|0.0|7|SUNBEAM OLD FASHION BREAD|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00071309045474|SLICED BREAD|COMMERCIAL BAKERY|-80.66939|1.4079464610753885|46|1
35.28326|fbc573dbcf908927c92e55574305385f75821fe8|2.89|2014-10-25 09:57:00|1.4094857484078087|1|5150000162|46|0.6158090578372145|0|26|123|-80.66939|19|35.28326|JELLY/JAMS|0.89|1|SMUCKER GRAPE JELLY|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00051500001622|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|24083801270c93eecd934bc97c5c91e59e633eb2|3.49|2014-11-27 07:18:00|80.669414401537693|1|7080003719|46|35.302041710208115|0|19|839|-80.737839|102|35.297134|STACK PACKS|0.99|19|SMITHFIELD DICED HAM|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|35.305725790410776|00070800037193|LUNCHMEATS|CASE READY MEATS|-80.66939|80.669393843943624|258|1
35.28326|af8256ff402c819377e8382fb453dc278420a2b1|3.79|2015-01-17 17:50:00|80.669414401537693|1|7203684009|46|35.302041707803518|0|19|5777|-80.784334|1530|35.384824|HOME BREWING|0.0|18|SAFALE #S-04 ALE YEAST|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|35.305725790410776|00072036840097|201 CENTRAL|GM|-80.66939|80.6694022620281|476|1
35.28326|5e428fa36e515440d7fd5eaa62d2f620430c9227|8.99|2014-12-07 15:49:00|1.4094857484078087|1|31254770153|46|0.6158090578372145|0|26|4030|-80.66939|1080|35.28326|ORAL RINSE-ANTISEPTIC|2.0|17|LISTERINE COOL MINT-42755|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00312547427555|ORAL HYGIENE|HBC|-80.66939|1.4079464610753885|46|1
35.28326|70055ba5050ac05d6a347af52ad72670c8cc8dfe|12.99|2015-02-07 18:52:00|1.4094857484078087|1|8378322200|46|0.6158090578372145|0|26|458|-80.66939|82|35.28326|CRAFT BEER|0.0|16|SIERRA NEVADA PALE ALE 12PK|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00083783222005|DOMESTIC BEER|BEER|-80.66939|1.4079464610753885|46|1
35.28326|32bf8e133476e9ba26a275d8de8fd78d991ef0eb|3.99|2014-12-30 13:26:00|1.4094857484078087|1|7203663995|46|0.6158090578372145|0|26|342|-80.66939|57|35.28326|FRESH MILK|0.0|3|HARRIS TEETER 2% MILK|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00072036639981|MILK|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|4d60d74de69ae8cace0ee94fbf8e0389af93a19f|9.58|2014-09-11 17:05:00|80.669414401537693|1|74759961702|46|35.302041708907709|0|19|16|-80.782849|3|35.372142|BAKING CHOCOLATE/CHIPS/MORSELS|0.0|1|GHIRADELLI SWEET BAKING COCOA|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|35.305725790410776|00747599617027|BAKING SUPPLIES|G1 GROCERY|-80.66939|80.66939938605897|122|2
35.28326|900aa30e117cd6d016aacc6261cf684ed39969ef|6.79|2015-02-12 07:25:00|80.669414401537693|1|30085075605|46|35.302041694565766|0|19|4243|-80.810056|1200|35.219587|NASAL PRODUCT-ADULT|0.0|17|AFRIN SINUS NASAL SPRAY-11201|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|35.305725790410776|00300854112011|COUGH/COLD/SINUS|HBC|-80.66939|80.669419945960428|401|1
35.28326|3876832ecc0a78fe19d4f49af4063dc6bd268e73|3.49|2015-02-01 13:01:00|1.4094857484078087|1|8265750080|46|0.6158090578372145|0|26|31|-80.66939|4|35.28326|NON CARBONATED WATER|0.0|1|DEER PARK 2.5 GAL SPRING WATER|74ca696e4baeaf4415a169f9a1a39fa51ec73b7b|1.297770837281219|0.61471665291522548|00082657500805|BOTTLED WATER|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.585842|6cd304534c9853592c958aa9ac5dfa57d8a174d8|2.39|2014-12-31 15:45:00|1.4102725052409182|4|73639310300|99|0.6210901099944839|0|1|247|-80.875654|39|35.585842|VEGETABLES-FLANKER|0.39|1|GLORY SND 27 GREENS COLLARD|78aaefff7d92885b541ecc1f31e1970add6d9de1|9.271796484786439|0.61833652052202714|00736393103003|VEGETABLES-CAN/JAR|G1 GROCERY|-80.875654|1.411546447003722|99|1
35.082768|7fa04168cf87313cf8d573167984ae396c84468a|5.59|2014-10-05 09:00:00|80.732732175546019|4||147|35.086815466033769|0|35|503|-80.850065|64|35.030252|FRESH GRAPES|0.37|4|RED GRAPES,SEEDLESS 12/16|7e8d1925740b0e396e4e859399c5273c09c311f3|0.27967029097388546|35.101032182271901|00204023000003|FRESH PRODUCE|PRODUCE|-80.732725|80.732730329036855|470|1
35.082768|7e85952a9fa1942af303a081d100cecabf27d384|2.27|2014-12-31 13:39:00|80.732732175546019|4|7203656065|147|35.086815466033769|0|35|315|-80.850065|52|35.030252|CHEESE-PROCESSED-SLICED|0.0|3|HT 2% SINGLE WRAP CHEESE|7e8d1925740b0e396e4e859399c5273c09c311f3|0.27967029097388546|35.101032182271901|00072036600844|CHEESE|DAIRY|-80.732725|80.732730329036855|470|1
35.082768|bf2f848041870f777578e6954f84f6641add2120|2.59|2015-02-25 17:00:00|80.732732175546019|4|7203652035|147|35.086815466033769|0|35|74|-80.850065|9|35.030252|RTE CEREAL ALL FAMILY|0.32|1|HT CER TOASTED OATS|7e8d1925740b0e396e4e859399c5273c09c311f3|0.27967029097388546|35.101032182271901|00072036520357|CEREAL|G1 GROCERY|-80.732725|80.732730329036855|470|1
35.082768|f768391781cd7c38e505a0fc1942176493543128|8.38|2014-11-01 11:03:00|80.732732175546019|4|4812110208|147|35.086815465818994|0|35|1037|-80.847383|164|35.024464|ENGLISH MUFFINS|2.09|7|THOMAS ENG MUFFN ORIG 6 PK PP|7e8d1925740b0e396e4e859399c5273c09c311f3|0.27967029097388546|35.101032182271901|00048121102081|BREAKFAST|COMMERCIAL BAKERY|-80.732725|80.73273056732836|317|2
35.082768|c09919026dfb82bbfa7abe18a274a3e62d6ebec3|7.49|2014-11-02 08:41:00|80.732732175546019|4|88133400051|147|35.086815466033769|0|35|36|-80.850065|10|35.030252|PREMIUM GROUND|0.0|1|DUNKIN'D ORIGNAL GROUND|7e8d1925740b0e396e4e859399c5273c09c311f3|0.27967029097388546|35.101032182271901|00881334000467|COFFEE|G1 GROCERY|-80.732725|80.732730329036855|470|1
35.082768|fae038017f151cad4ddd9951860be8b09b40f5d4|7.49|2015-01-06 12:56:00|80.732732175546019|4|88133400051|147|35.086815466033769|0|35|36|-80.850065|10|35.030252|PREMIUM GROUND|0.0|1|DUNKIN'D ORIGNAL GROUND|7e8d1925740b0e396e4e859399c5273c09c311f3|0.27967029097388546|35.101032182271901|00881334000467|COFFEE|G1 GROCERY|-80.732725|80.732730329036855|470|1
35.082768|da2f08db3ab071baa6c36e5dad228ac89cfcfa33|5.99|2014-12-26 10:33:00|80.732732175546019|4|7203688215|147|35.086815466033769|0|35|500|-80.850065|64|35.030252|FRESH APPLES|0.0|4|HT GALA APPLE 5LB|7e8d1925740b0e396e4e859399c5273c09c311f3|0.27967029097388546|35.101032182271901|00072036882158|FRESH PRODUCE|PRODUCE|-80.732725|80.732730329036855|470|1
35.082768|5f86b77429b924eea247f454c3d845829f498960|0.57|2014-10-16 16:56:00|80.732732175546019|4||147|35.086815466033769|0|35|502|-80.850065|64|35.030252|FRESH BANANAS|0.0|4|BANANAS, YELLOW|7e8d1925740b0e396e4e859399c5273c09c311f3|0.27967029097388546|35.101032182271901|00204011000008|FRESH PRODUCE|PRODUCE|-80.732725|80.732730329036855|470|1
35.082768|23ee053517ae8d1b206090cc0754c991601916ae|3.0|2014-11-22 10:12:00|80.732732175546019|4|7203608990|147|35.086815466033769|0|35|82|-80.850065|11|35.030252|VINEGAR|0.5|1|HT VINEGAR BALSAMIC|7e8d1925740b0e396e4e859399c5273c09c311f3|0.27967029097388546|35.101032182271901|00072036089908|CONDIMENTS|G1 GROCERY|-80.732725|80.732730329036855|470|1
35.082768|bdc8dced58ef5876a34d7ce8ba67d206f5ed1e6d|0.54|2015-01-11 09:55:00|80.732732175546019|4||147|35.086815466033769|0|35|502|-80.850065|64|35.030252|FRESH BANANAS|0.0|4|BANANAS, YELLOW|7e8d1925740b0e396e4e859399c5273c09c311f3|0.27967029097388546|35.101032182271901|00204011000008|FRESH PRODUCE|PRODUCE|-80.732725|80.732730329036855|470|1
35.082768|9d6fd11d76220c689df9fbd1516615bb95c5c09c|3.69|2014-09-20 09:45:00|80.732732175546019|4|7518500003|147|35.086815467613945|0|35|1033|-80.816172|163|35.059823|HAMBURGER|0.0|7|MARTIN'S POTATO SANDWICH ROLLS|7e8d1925740b0e396e4e859399c5273c09c311f3|0.27967029097388546|35.101032182271901|00075185000039|BUNS/ROLLS|COMMERCIAL BAKERY|-80.732725|80.732728048954272|66|1
35.082768|ce89907f176815ab870ae9190d1303a3bc5d7a01|3.69|2014-12-20 14:09:00|80.732732175546019|4|7518500003|147|35.086815466033769|0|35|1033|-80.850065|163|35.030252|HAMBURGER|0.0|7|MARTIN'S POTATO SANDWICH ROLLS|7e8d1925740b0e396e4e859399c5273c09c311f3|0.27967029097388546|35.101032182271901|00075185000039|BUNS/ROLLS|COMMERCIAL BAKERY|-80.732725|80.732730329036855|470|1
35.082768|11e6d9abe8641384c470c3fb2d495542790f6991|2.99|2014-12-21 09:46:00|80.732732175546019|4|81204900640|147|35.086815466033769|0|35|504|-80.850065|64|35.030252|FRESH BERRIES|0.0|4|BLUEBERRIES 6 OZ|7e8d1925740b0e396e4e859399c5273c09c311f3|0.27967029097388546|35.101032182271901|00817621010109|FRESH PRODUCE|PRODUCE|-80.732725|80.732730329036855|470|1
35.082768|c89322429813d6f12744ddc664cecc46396ab065|4.45|2014-12-06 11:10:00|80.732732175546019|4||147|35.086815466033769|0|35|507|-80.850065|64|35.030252|FRESH ORANGES|0.29|4|NAVEL ORANGE, LRG|7e8d1925740b0e396e4e859399c5273c09c311f3|0.27967029097388546|35.101032182271901|00233107000004|FRESH PRODUCE|PRODUCE|-80.732725|80.732730329036855|470|5
35.082768|fa6d64efd8f7132231d2565c4f889273db51a9b4|4.45|2014-12-07 08:59:00|80.732732175546019|4||147|35.086815466033769|0|35|507|-80.850065|64|35.030252|FRESH ORANGES|0.29|4|NAVEL ORANGE, LRG|7e8d1925740b0e396e4e859399c5273c09c311f3|0.27967029097388546|35.101032182271901|00233107000004|FRESH PRODUCE|PRODUCE|-80.732725|80.732730329036855|470|5
35.082768|818c418224a293582e73b92dfa1dd558d5331aa4|5.0|2014-11-26 11:11:00|80.732732175546019|4|7203698557|147|35.086815466033769|0|35|424|-80.850065|72|35.030252|NFS-FACIAL TISSUE|0.0|1|HT FACIAL TISSUE LOTION|7e8d1925740b0e396e4e859399c5273c09c311f3|0.27967029097388546|35.101032182271901|00072036985583|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.732725|80.732730329036855|470|4
35.082768|fe055b08827bff360bad24beb2df27a297c73dc9|3.59|2014-10-19 09:19:00|80.732732175546019|4|7433610102|147|35.086815466033769|0|35|342|-80.850065|57|35.030252|FRESH MILK|0.0|3|HIGHLAND CREST 2% REDUCE FAT|7e8d1925740b0e396e4e859399c5273c09c311f3|0.27967029097388546|35.101032182271901|00074336101021|MILK|DAIRY|-80.732725|80.732730329036855|470|1
35.082768|f352ca4b45f8aa2a56ebe128746eebeff3edf785|7.99|2015-03-04 16:53:00|80.732732175546019|4|68954408301|147|35.086815465818994|0|35|685|-80.847383|61|35.024464|GREEK|0.0|3|FAGE TOTAL 2%|7e8d1925740b0e396e4e859399c5273c09c311f3|0.27967029097388546|35.101032182271901|00689544083023|YOGURT|DAIRY|-80.732725|80.73273056732836|317|1
35.082768|460a6ecca5c48a9107628fe6efe7426ed3c7ac91|3.98|2014-11-29 11:05:00|80.732732175546019|4|88596708120|147|35.086815466033769|0|35|422|-80.850065|71|35.030252|NFS-REMAIN LAUNDRY SUPPL|0.0|1|NIAGARA STARCH|7e8d1925740b0e396e4e859399c5273c09c311f3|0.27967029097388546|35.101032182271901|00885967081206|LAUNDRY SUPPLIES|G1 GROCERY|-80.732725|80.732730329036855|470|2
35.082768|3d162a0397d17caae64d42a841a5f73519ac3c58|1.97|2015-01-29 15:57:00|80.732732175546019|4|7203603118|147|35.086815465818994|0|35|209|-80.847383|20|35.024464|POWDERED SOFT DRINKS|0.0|1|HT DRINK MIX FRUIT PUNCH QT|7e8d1925740b0e396e4e859399c5273c09c311f3|0.27967029097388546|35.101032182271901|00072036031181|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.732725|80.73273056732836|317|1
35.40953|2e83cf428c90740f35e94fb5a3f1cb88f89966a9|8.99|2015-03-08 18:43:00|80.89430079996653|2|61278110261|209|35.422821403014979|0|32|265|-80.995484|307|35.444064|FROZEN PIES|2.0|5|M CALLENDER CHERRY CRUNCH PIE|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|35.45572462568753|00612781101359|DESSERTS FROZEN|FROZEN|-80.86175|80.861754060610338|121|1
35.40953|e83a61c8b489077f6e8438ef945ec99921aa50cb|8.99|2014-12-14 15:54:00|1.4102725052409182|2|61278110261|209|0.6180128850837077|0|1|265|-80.86175|307|35.40953|FROZEN PIES|4.5|5|M CALLENDER CHERRY CRUNCH PIE|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00612781101359|DESSERTS FROZEN|FROZEN|-80.86175|1.4113037764245249|209|1
35.40953|00a09784724241ee42b39fa5c824e5cc4a449742|2.39|2015-01-25 16:16:00|80.89430079996653|2|7203695175|209|35.422821403014979|0|32|1607|-80.995484|371|35.444064|FROZEN DOUGH (BREAD)|0.9|14|FRESH LRG FRENCH BREAD|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|35.45572462568753|00072036951755|BREAD|BAKERY|-80.86175|80.861754060610338|121|1
35.40953|716926ee5dc7ad50c2ff1baf605a9f110bb547a1|2.58|2014-11-01 17:12:00|80.89430079996653|2|4920005675|209|35.422821403014979|0|32|224|-80.995484|35|35.444064|SUGAR-BROWN|0.6|1|DOMINO LT BRWN SUGAR-BOX|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|35.45572462568753|00049200056752|SUGAR/SUBSTITUTES|G1 GROCERY|-80.86175|80.861754060610338|121|2
35.40953|4084dccacec527ffdc289c819a7231c0c9b68216|1.89|2015-03-03 14:03:00|80.89430079996653|2|7203663214|209|35.422821402542247|0|32|330|-80.861571|55|35.444615|EGGS|0.0|3|HT GRADE A    EX-LARGE EGGS|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|35.45572462568753|00072036632142|EGGS FRESH|DAIRY|-80.86175|80.861755950576324|340|1
35.40953|8a9051239fc8cd9b66955f6679068caebf342735|1.89|2015-01-18 15:56:00|80.89430079996653|2|7203663214|209|35.422821402542247|0|32|330|-80.861571|55|35.444615|EGGS|0.0|3|HT GRADE A    EX-LARGE EGGS|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|35.45572462568753|00072036632142|EGGS FRESH|DAIRY|-80.86175|80.861755950576324|340|1
35.40953|dd2209c23be20d6cd874faeb149b9732a31ff9d0|31.92|2014-12-07 17:53:00|1.4102725052409182|2|7203661016|209|0.6180128850837077|0|1|297|-80.86175|49|35.40953|GROUND BEEF|3.04|2|GROUND CHUCK 80% LEAN 2 LB|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00072036610164|BEEF|MEAT|-80.86175|1.4113037764245249|209|4
35.40953|2d1e2f7256ec6fd87272d58707cb40b9388f1a49|7.99|2014-12-05 20:12:00|80.89430079996653|2|4100032816|209|35.422821402542247|0|32|1247|-80.861571|37|35.444615|SINGLES PODS CUPS TEA|1.99|1|LIPTON K-CUP TEA INDULGE BLACK|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|35.45572462568753|00041000328527|TEA|G1 GROCERY|-80.86175|80.861755950576324|340|1
35.40953|0eba8b269022c258a94011992aea155a70a6d085|2.99|2015-01-09 20:24:00|80.89430079996653|2|4144900210|209|35.422821402542247|0|32|231|-80.861571|37|35.444615|INSTANT TEA|1.5|1|ALPINE SPICED CIDER REGULAR|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|35.45572462568753|00041449002101|TEA|G1 GROCERY|-80.86175|80.861755950576324|340|1
35.40953|8ca092672a740b8175423d3e823adc89b3991202|7.99|2014-12-05 20:11:00|80.89430079996653|2|4100032816|209|35.422821402542247|0|32|1247|-80.861571|37|35.444615|SINGLES PODS CUPS TEA|1.0|1|LIPTON K-CUP TEA INDULGE BLACK|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|35.45572462568753|00041000328527|TEA|G1 GROCERY|-80.86175|80.861755950576324|340|1
35.40953|07c9d6f426f65e8ccee2ace04be6596e84e4cfba|3.85|2014-09-20 18:54:00|1.4102725052409182|2|3800001611|209|0.6180128850837077|0|1|61|-80.86175|9|35.40953|RTE CEREAL ADULT|1.36|1|KELLOGG SPECIAL K MULTI GRAIN|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00038000915567|CEREAL|G1 GROCERY|-80.86175|1.4113037764245249|209|1
35.40953|038ad563473d47b804de88e54617b116e4ea6d75|3.99|2015-02-22 14:10:00|1.4102725052409182|2|4400002854|209|0.6180128850837077|0|1|1248|-80.86175|12|35.40953|SANDWICH COOKIES|1.49|1|OREO GOLDEN DOUBLE STUF|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00044000025403|COOKIES|G1 GROCERY|-80.86175|1.4113037764245249|209|1
35.40953|1cabdd2234071ca491704f5cace0707e3349f7c7|3.99|2014-09-28 18:36:00|1.4102725052409182|2|4400002854|209|0.6180128850837077|0|1|1248|-80.86175|12|35.40953|SANDWICH COOKIES|1.49|1|OREO GOLDEN DOUBLE STUF|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00044000025403|COOKIES|G1 GROCERY|-80.86175|1.4113037764245249|209|1
35.40953|b23f3b197b0c8eb52b270b414118563c7404dffd|5.94|2014-12-31 18:05:00|1.4102725052409182|2|4173600180|209|0.6180128850837077|0|1|194|-80.86175|30|35.40953|OLIVE OIL|4.0|1|FILIPPO BERIO PURE OLIVE OIL|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00041736001800|SHORTENING/OIL|G1 GROCERY|-80.86175|1.4113037764245249|209|2
35.40953|3af49e90a7c8f3f26d1866590625ac563c247de3|9.38|2014-12-02 18:56:00|1.4102725052409182|2|4900002468|209|0.6180128850837077|0|1|54|-80.86175|8|35.40953|DIET|2.72|23|DIET COKE .5 LITER/6 PK.|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.86175|1.4113037764245249|209|2
35.40953|06892b69a58243e259ec4a4d1ee18c3cb4811ce5|3.65|2014-11-09 17:11:00|1.4102725052409182|2|4610000012|209|0.6180128850837077|0|1|318|-80.86175|52|35.40953|SHREDDED/GRATED CHEESE|1.15|3|SARGENTO OTB 4 CHSE MEX FINE C|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00046100000922|CHEESE|DAIRY|-80.86175|1.4113037764245249|209|1
35.40953|dacb54b1447272563faaabfcedd1fcd7012e3450|3.95|2014-10-05 17:50:00|1.4102725052409182|2|4610000012|209|0.6180128850837077|0|1|318|-80.86175|52|35.40953|SHREDDED/GRATED CHEESE|1.97|3|SARGENTO OTB 4 CHSE MEX FINE C|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00046100000922|CHEESE|DAIRY|-80.86175|1.4113037764245249|209|1
35.40953|d15448232faab3a30445055b040a1b9c9a264a1b|9.7|2014-12-20 18:33:00|1.4102725052409182|2|7790011553|209|0.6180128850837077|0|1|361|-80.86175|105|35.40953|BREAKFAST SAUSAGE|3.04|19|JIMMY DEAN MILD SAUSAGE|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00077900115530|BREAKFAST SAUSAGE|CASE READY MEATS|-80.86175|1.4113037764245249|209|2
35.40953|2fe0c203ed0e9df82414c8bfe203b8be082231c9|19.38|2014-10-17 18:15:00|1.4102725052409182|2|88133400051|209|0.6180128850837077|0|1|36|-80.86175|10|35.40953|PREMIUM GROUND|7.4|1|DUNKIN'D ORIGNAL GROUND|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00881334000467|COFFEE|G1 GROCERY|-80.86175|1.4113037764245249|209|2
35.40953|8bcb2339ffd926c86d5b82f67273c28745d75483|3.19|2014-11-26 15:41:00|1.4102725052409182|2|7225002910|209|0.6180128850837077|0|1|1039|-80.86175|166|35.40953|DINNER ROLLS|0.7|7|MERITA 24CT DINNER ROLLS|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00072250029100|MEAL ACCOMPANIMENT|COMMERCIAL BAKERY|-80.86175|1.4113037764245249|209|1
35.40953|8805807178e43a1bb2699c99ccd2697ee79950d7|6.99|2015-02-01 13:58:00|80.89430079996653|2|7203695357|209|35.422821403014979|0|32|1295|-80.995484|383|35.444064|PIES PASTRY CASE TAX|3.02|14|"9"" KEY LIME PIE"|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|35.45572462568753|00072036953575|PASTRY CASE|BAKERY|-80.86175|80.861754060610338|121|1
35.40953|4e32329f1d902425c5cd0344e62934ef4f680062|11.32|2015-02-09 16:34:00|1.4102725052409182|2|20598400000|209|0.6180128850837077|0|1|1822|-80.86175|410|35.40953|BH CHICKEN|2.06|6|BOARS HEAD EVERROAST CKN BRST|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00205984000002|BH MEAT|DELI|-80.86175|1.4113037764245249|209|1
35.40953|8c0c7957f755930b8ecc88cb420989ab609cea9b|5.82|2015-01-04 18:37:00|1.4102725052409182|2|20598400000|209|0.6180128850837077|0|1|1822|-80.86175|410|35.40953|BH CHICKEN|0.0|6|BOARS HEAD EVERROAST CKN BRST|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00205984000002|BH MEAT|DELI|-80.86175|1.4113037764245249|209|1
35.40953|809121069dcd7d2b9fd00c8ca4b3900abecdabc7|4.19|2015-02-15 17:08:00|1.4102725052409182|2|4812110208|209|0.6180128850837077|0|1|1037|-80.86175|164|35.40953|ENGLISH MUFFINS|2.1|7|THOMAS ENG MUFFN ORIG 6 PK PP|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00048121102081|BREAKFAST|COMMERCIAL BAKERY|-80.86175|1.4113037764245249|209|1
35.40953|38a6ec479041d95d97b895caaff5f3e778f9c0ff|8.38|2015-01-17 18:21:00|80.89430079996653|2|4812110208|209|35.422821399255355|0|32|1037|-80.762919|164|35.442529|ENGLISH MUFFINS|2.1|7|THOMAS ENG MUFFN ORIG 6 PK PP|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|35.45572462568753|00048121102081|BREAKFAST|COMMERCIAL BAKERY|-80.86175|80.861762921485493|471|2
35.40953|b65e59ad43cbe68fbadbdf46bc4e881614abf0a5|7.98|2014-12-22 14:58:00|1.4102725052409182|2|2850010245|209|0.6180128850837077|0|1|112|-80.86175|14|35.40953|PIE & PASTRY FILLING|2.98|1|LUCKY LF PREM CHERRY PIE FILL|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00028500102451|DESSERTS/GELS/SYRUPS|G1 GROCERY|-80.86175|1.4113037764245249|209|2
35.40953|6f11b4fa4867655d65f2fd1ea5ecb4f658a12d65|19.99|2014-11-16 15:48:00|1.4102725052409182|2|20641300000|209|0.6180128850837077|0|1|1653|-80.86175|381|35.40953|CELEBRATION CAKES|0.0|14|SPEC ORDER MARB 1/4 SHT CAKE|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00206413000006|CAKES|BAKERY|-80.86175|1.4113037764245249|209|1
35.40953|e6ec3956cf582501a07b32e6dae16dccfa01b40b|5.79|2014-10-19 14:42:00|80.89430079996653|2|20165500000|209|35.422821403014979|0|32|297|-80.995484|49|35.444064|GROUND BEEF|0.73|2|HT PREMIUM GRND BEEF 80% LEAN|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|35.45572462568753|00201655000005|BEEF|MEAT|-80.86175|80.861754060610338|121|1
35.40953|44a72b8fce286fec955e41d6127e17431feb6d90|0.79|2014-10-03 14:53:00|1.4102725052409182|2||209|0.6180128850837077|0|1|532|-80.86175|64|35.40953|FRESH CUCUMBERS|0.1|4|COO CUCUMBERS S/S|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00204062000002|FRESH PRODUCE|PRODUCE|-80.86175|1.4113037764245249|209|1
35.40953|651afe0d36e2052cca478f207a4f6964de7b9796|25.07|2015-02-02 19:11:00|1.4102725052409182|2|20165500000|209|0.6180128850837077|0|1|297|-80.86175|49|35.40953|GROUND BEEF|0.71|2|HT PREMIUM GRND BEEF 80% LEAN|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00201655000005|BEEF|MEAT|-80.86175|1.4113037764245249|209|5
35.40953|83ce0df9cfbf7a161c36e5898d1de4122d5d7cc3|3.99|2014-09-23 17:54:00|1.4102725052409182|2|7203663995|209|0.6180128850837077|0|1|342|-80.86175|57|35.40953|FRESH MILK|0.0|3|HARRIS TEETER 1% MILK|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00072036631275|MILK|DAIRY|-80.86175|1.4113037764245249|209|1
35.40953|74449feb8a612f582372c6bc1343294c3301a3ee|3.49|2015-02-07 18:28:00|1.4102725052409182|2|7203663995|209|0.6180128850837077|0|1|342|-80.86175|57|35.40953|FRESH MILK|1.72|3|HARRIS TEETER 1% MILK|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00072036631275|MILK|DAIRY|-80.86175|1.4113037764245249|209|1
35.40953|f85a0e37bee7e8a1364c944de51f67a092558c6a|3.99|2014-10-26 20:11:00|1.4102725052409182|2|7203663995|209|0.6180128850837077|0|1|342|-80.86175|57|35.40953|FRESH MILK|0.0|3|HARRIS TEETER 1% MILK|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00072036631275|MILK|DAIRY|-80.86175|1.4113037764245249|209|1
35.40953|9c018fbe3c7a105e39b9d4448411c5d4484140eb|3.29|2014-09-18 16:27:00|1.4102725052409182|2|20668800000|209|0.6180128850837077|0|1|1830|-80.86175|415|35.40953|FFM SLICING CHEESE|0.0|6|HT WHITE AMERICAN|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00206688000008|SLICING CHEESE|DELI|-80.86175|1.4113037764245249|209|1
35.40953|ae84325e6535982f184ca39ad389d17510aad380|3.99|2014-10-18 10:13:00|1.4102725052409182|2|4000015140|209|0.6180128850837077|0|1|46|-80.86175|7|35.40953|PKG CHOC|0.49|1|3 MUSKETEER FUN SIZE|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00040000151227|CANDY|G1 GROCERY|-80.86175|1.4113037764245249|209|1
35.40953|b6c827475db37e8848f7927275b65a6192ddbc9a|19.98|2014-09-15 19:13:00|1.4102725052409182|2|4200044517|209|0.6180128850837077|0|1|426|-80.86175|72|35.40953|NFS-PAPER TOWELS|6.0|1|BRAWNY 6 BIG ROLL PICK A SIZE|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00042000445177|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.86175|1.4113037764245249|209|2
35.40953|13a50a4a5d3e53ef10056ac487bc119aedaaf8dd|4.78|2015-01-10 14:44:00|1.4102725052409182|2|1340934115|209|0.6180128850837077|0|1|68|-80.86175|11|35.40953|BARBECUE SAUCES|1.02|1|SWEET BABY RAY BBQ SC HONEY|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00013409341155|CONDIMENTS|G1 GROCERY|-80.86175|1.4113037764245249|209|2
35.40953|b5cf5bd79375e8b96ed1841fbc39cc397925a53a|4.0|2014-12-23 17:24:00|1.4102725052409182|2|4300000953|209|0.6180128850837077|0|1|272|-80.86175|307|35.40953|TOPPINGS FROZEN|2.02|5|COOL WHIP EXTRA CREAMY|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00043000002742|DESSERTS FROZEN|FROZEN|-80.86175|1.4113037764245249|209|2
35.40953|9c14be5ff1ac2c402f947dea119d22e8dd10fd25|7.08|2014-11-20 19:24:00|1.4102725052409182|2|3800001611|209|0.6180128850837077|0|1|61|-80.86175|9|35.40953|RTE CEREAL ADULT|0.0|1|KELLOGG SPECIAL K FRUIT YOGURT|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00038000787119|CEREAL|G1 GROCERY|-80.86175|1.4113037764245249|209|4
35.40953|90568182d79fdf85ccd7094ca0d2e649dceb0c6f|5.29|2014-11-03 19:27:00|1.4102725052409182|2|7203670704|209|0.6180128850837077|0|1|252|-80.86175|45|35.40953|PREMIUM ICE CREAM|1.3|5|I/OHT ALL NATURAL PEPP BARK IC|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00072036707055|ICE CREAM|FROZEN|-80.86175|1.4113037764245249|209|1
35.40953|31eb549e6293a778a80a27da6d2ebe897a0ef703|8.9|2014-09-11 18:42:00|80.89430079996653|2|20543600000|209|35.422821403014979|0|32|1832|-80.995484|415|35.444064|BH SLICING CHEESE|0.0|6|BOARS HEAD MONTEREY JACK CHSE|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|35.45572462568753|00205436000000|SLICING CHEESE|DELI|-80.86175|80.861754060610338|121|1
35.40953|e1d6bb7f5f02563ae78a35f02a0a4e25cf2ee502|2.5|2014-11-25 15:05:00|80.89430079996653|2|4900005537|209|35.422821402542247|0|32|54|-80.861571|8|35.444615|DIET|0.52|23|COKE ZERO 1.25 LITER BOTTLE|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|35.45572462568753|00049000055412|CARBONATED BEVERAGES|BEVERAGE|-80.86175|80.861755950576324|340|2
35.40953|ffbd833891131b84aa0da1c2a65d65a749de580e|0.99|2014-12-09 15:38:00|1.4102725052409182|2||209|0.6180128850837077|0|1|535|-80.86175|64|35.40953|FRESH GREENS|0.0|4|COO KALE, BULK|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00204627000003|FRESH PRODUCE|PRODUCE|-80.86175|1.4113037764245249|209|1
35.40953|9200c473aede2eb812fcc8b18897c697971c6ee9|7.38|2015-01-11 12:52:00|1.4102725052409182|2|4400001570|209|0.6180128850837077|0|1|1256|-80.86175|13|35.40953|WHOLESOME CRACKERS|1.38|1|TOASTED CHIPS ORIGINAL|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00044000015596|CRACKERS|G1 GROCERY|-80.86175|1.4113037764245249|209|2
35.40953|cf751a95fb9e7c554737d486a9754f6e61fc06e4|4.58|2015-01-06 19:26:00|1.4102725052409182|2|7203663996|209|0.6180128850837077|0|1|342|-80.86175|57|35.40953|FRESH MILK|0.82|3|HARRIS TEETER 1%  MILK|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00072036631305|MILK|DAIRY|-80.86175|1.4113037764245249|209|2
35.40953|fe3e01e1c899ce6473e05378dc4139dd65339ea7|3.75|2014-11-16 13:19:00|1.4102725052409182|2|2400016286|209|0.6180128850837077|0|1|245|-80.86175|39|35.40953|VEGETABLES-CORE|1.25|1|DEL MONTE GRN BEANS FRENCH|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|0.61833652052202714|00024000162896|VEGETABLES-CAN/JAR|G1 GROCERY|-80.86175|1.4113037764245249|209|3
35.40953|94e0837825e72dd15293afd2af56ed58fad486db|1.55|2014-10-30 14:21:00|80.89430079996653|2|2920000212|209|35.422821402542247|0|32|149|-80.861571|23|35.444615|WHSE PASTA CORE|0.55|1|MUELLER THIN SPAGHETTI|8131f3cc069286da8e26ed029571c46fa675cee4|0.9184038792115339|35.45572462568753|00029200002140|PASTA|G1 GROCERY|-80.86175|80.861755950576324|340|1
35.140781|a853c71d4886f55a92ef4b72f55142a0833705a0|1.57|2014-11-03 15:45:00|80.632521683083056|3||39|35.192060774618689|0|39|502|-80.661096|64|35.172688|FRESH BANANAS|0.0|4|BANANAS, YELLOW|8459144dc4eb4f006173021c7c08de3acdc7eb55|3.5433086357791366|35.177497916598789|00204011000008|FRESH PRODUCE|PRODUCE|-80.62331|80.623320091295128|474|1
35.140781|9683b9b33b8bb8902f9e8c33e8aaa866846fe6e0|1.55|2015-01-24 14:21:00|80.632521683083056|3||39|35.192060774618689|0|39|502|-80.661096|64|35.172688|FRESH BANANAS|0.0|4|BANANAS, YELLOW|8459144dc4eb4f006173021c7c08de3acdc7eb55|3.5433086357791366|35.177497916598789|00204011000008|FRESH PRODUCE|PRODUCE|-80.62331|80.623320091295128|474|1
35.140781|79971c8276e7ab7178fa1b84fe855fdeafc6f407|1.86|2014-10-03 16:01:00|80.632521683083056|3||39|35.192060774618689|0|39|502|-80.661096|64|35.172688|FRESH BANANAS|0.0|4|BANANAS, YELLOW|8459144dc4eb4f006173021c7c08de3acdc7eb55|3.5433086357791366|35.177497916598789|00204011000008|FRESH PRODUCE|PRODUCE|-80.62331|80.623320091295128|474|1
35.140781|8dfede50e1327429bfae3f5b87499ee0fd049b2e|4.13|2014-09-25 14:32:00|80.632521683083056|3|20165700000|39|35.192060774618689|0|39|297|-80.661096|49|35.172688|GROUND BEEF|0.92|2|HT GROUND BEEF CHUCK 80% LEAN|8459144dc4eb4f006173021c7c08de3acdc7eb55|3.5433086357791366|35.177497916598789|00201657000003|BEEF|MEAT|-80.62331|80.623320091295128|474|1
35.140781|bb2308696e597260aa4bf194208e3c7e99bef77e|6.79|2015-02-09 17:30:00|80.632521683083056|3|9113135067|39|35.192060774618689|0|39|84|-80.661096|11|35.172688|CONDIMENTS-DSD VENDORS|0.0|1|BEE CITY HONEY BEARS|8459144dc4eb4f006173021c7c08de3acdc7eb55|3.5433086357791366|35.177497916598789|00091131350676|CONDIMENTS|G1 GROCERY|-80.62331|80.623320091295128|474|1
35.140781|be0761ee278896f5446b2679ecafde033bc209be|11.98|2015-01-04 13:43:00|80.632521683083056|3|76401420805|39|35.192060774618689|0|39|356|-80.661096|104|35.172688|GOURMET SAUSAGE|0.0|19|AIDELLS CAJUN ANDOUILLE SAUSAG|8459144dc4eb4f006173021c7c08de3acdc7eb55|3.5433086357791366|35.177497916598789|00764014458058|DINNER SAUSAGE|CASE READY MEATS|-80.62331|80.623320091295128|474|2
35.082768|a188ea3cb506f1fc8e4c192714e145007365debd|0.45|2014-12-24 13:05:00|1.4091206135396188|4||147|0.6123098123133061|0|47|524|-80.732725|64|35.082768|FRESH PROD FRESH ONIONS|0.0|4|COO YELLOW ONIONS, LRG|88adc9b2431567ae3a9d0afeec18f19f851e83a1|1.0450148292139363|0.61242566243833529|00204665000003|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|1
35.082768|5813c24689666594451b979f6b6916f4ebd6ac48|53.940000000000005|2014-12-22 12:18:00|1.4091206135396188|4|8072000062|147|0.6123098123133061|0|47|9927|-80.732725|884|35.082768|NFS FV CHARDONNAY|0.0|13|GLEN ELLEN CHAARD RES|88adc9b2431567ae3a9d0afeec18f19f851e83a1|1.0450148292139363|0.61242566243833529|00080720000627|FIGHTING VARIETL($0-$3.99)|WINE|-80.732725|1.409051865357139|147|6
35.082768|868489446f5d162103e61752489c5815689a1007|19.98|2015-02-16 11:40:00|1.4091206135396188|4|8072000062|147|0.6123098123133061|0|47|9927|-80.732725|884|35.082768|NFS FV CHARDONNAY|0.0|13|GLEN ELLEN CHAARD RES|88adc9b2431567ae3a9d0afeec18f19f851e83a1|1.0450148292139363|0.61242566243833529|00080720000627|FIGHTING VARIETL($0-$3.99)|WINE|-80.732725|1.409051865357139|147|2
35.082768|6c39bc2d5714a8eae7e58d5b3d34d9d84d12708a|19.98|2015-01-22 12:26:00|1.4091206135396188|4|8072000062|147|0.6123098123133061|0|47|9927|-80.732725|884|35.082768|NFS FV CHARDONNAY|0.0|13|GLEN ELLEN CHAARD RES|88adc9b2431567ae3a9d0afeec18f19f851e83a1|1.0450148292139363|0.61242566243833529|00080720000627|FIGHTING VARIETL($0-$3.99)|WINE|-80.732725|1.409051865357139|147|2
35.082768|6dae1c7167ed727e749ba0c1cd4f62ba9893cba3|2.0100000000000002|2015-02-25 11:58:00|1.4091206135396188|4|7203641111|147|0.6123098123133061|0|47|242|-80.732725|39|35.082768|CANNED BEANS|0.0|1|HT BEANS PINTO|88adc9b2431567ae3a9d0afeec18f19f851e83a1|1.0450148292139363|0.61242566243833529|00072036411112|VEGETABLES-CAN/JAR|G1 GROCERY|-80.732725|1.409051865357139|147|3
35.082768|a90b2d0bfcd32ef3985ff2a410e6244313a7c56c|2.78|2015-02-01 14:22:00|1.4091206135396188|4|5210094269|147|0.6123098123133061|0|47|80|-80.732725|34|35.082768|SEASONING PACKETS|0.78|1|E  MC CHILI SEASONING MIX|88adc9b2431567ae3a9d0afeec18f19f851e83a1|1.0450148292139363|0.61242566243833529|00052100091501|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.732725|1.409051865357139|147|2
35.082768|3633b6c73c4afb319a8638e08308caf562789f6c|6.0|2015-03-06 13:44:00|1.4091206135396188|4|7203698062|147|0.6123098123133061|0|47|54|-80.732725|8|35.082768|DIET|0.0|23|HT DIET TONIC WATER 2 LTR|88adc9b2431567ae3a9d0afeec18f19f851e83a1|1.0450148292139363|0.61242566243833529|00072036980625|CARBONATED BEVERAGES|BEVERAGE|-80.732725|1.409051865357139|147|4
35.082768|898f75d6a5ed42c4333992dd45692ffd3e0c0db7|7.08|2014-12-28 11:53:00|80.732732175546019|4|7203657031|147|35.09789175327596|0|35|322|-80.562829|53|35.006282|SOUR CREAM|0.0|3|HT SOUR CREAM|88adc9b2431567ae3a9d0afeec18f19f851e83a1|1.0450148292139363|35.101032182271901|00072036570314|CULTURES|DAIRY|-80.732725|80.732725512795|60|4
35.082768|885bf833f561ab6f238f8e711776eb88b4ad8e41|13.37|2015-02-12 12:31:00|1.4091206135396188|4|20331300000|147|0.6123098123133061|0|47|641|-80.732725|137|35.082768|PREMIUM PORK|0.0|2|PORK LOIN CHOPS BONE-IN CUSTOM|88adc9b2431567ae3a9d0afeec18f19f851e83a1|1.0450148292139363|0.61242566243833529|00203314000005|PORK|MEAT|-80.732725|1.409051865357139|147|1
35.082768|80eeff42539d54aba830b07125399e4e48603176|47.85|2014-12-23 17:18:00|80.732732175546019|4|20396000000|147|35.097891753221013|0|35|978|-80.78468|202|35.096737|SMOKED MEATS|9.59|2|SMFD SPIRAL CRUNCHY GLAZED HAM|88adc9b2431567ae3a9d0afeec18f19f851e83a1|1.0450148292139363|35.101032182271901|00203960000008|SMOKED HAMS|MEAT|-80.732725|80.732726656903608|30|1
35.082768|2e46fcfc14f8179d7080dae79229495075b71cb6|3.99|2015-01-16 18:08:00|1.4091206135396188|4|4470003050|147|0.6123098123133061|0|47|840|-80.732725|102|35.082768|TUBS|0.49|19|OM DELI FRESH ROTISSERE CHCKEN|88adc9b2431567ae3a9d0afeec18f19f851e83a1|1.0450148292139363|0.61242566243833529|00044700030998|LUNCHMEATS|CASE READY MEATS|-80.732725|1.409051865357139|147|1
35.082768|4f904743f8022b1698c79c55087777785a1f5be9|8.98|2015-01-07 13:20:00|1.4091206135396188|4|4470003050|147|0.6123098123133061|0|47|840|-80.732725|102|35.082768|TUBS|1.98|19|OM BOLD ITALIAN HERB TURKEY|88adc9b2431567ae3a9d0afeec18f19f851e83a1|1.0450148292139363|0.61242566243833529|00044700072820|LUNCHMEATS|CASE READY MEATS|-80.732725|1.409051865357139|147|2
35.082768|5a9fe7c900f2cca6c687c254a61007891a4d284c|4.99|2015-01-29 14:15:00|1.4091206135396188|4|4082201114|147|0.6123098123133061|0|47|1878|-80.732725|435|35.082768|HUMMUS|2.5|6|ROASTED RED PEPPER HUMMUS|88adc9b2431567ae3a9d0afeec18f19f851e83a1|1.0450148292139363|0.61242566243833529|00040822011549|SALADS|DELI|-80.732725|1.409051865357139|147|1
35.082768|81f500eb0ad99d890e562b3cb0b61dd81d37a28b|13.99|2015-02-22 16:27:00|1.4091206135396188|4|8066095787|147|0.6123098123133061|0|47|459|-80.732725|83|35.082768|IMPORT BEER|0.0|16|NEGRA MODELO 12PK BOTTLES|88adc9b2431567ae3a9d0afeec18f19f851e83a1|1.0450148292139363|0.61242566243833529|00080660957876|IMPORT BEER|BEER|-80.732725|1.409051865357139|147|1
35.082768|616153d6499159041140a4dd2726548a42dc8b0e|15.99|2015-03-01 17:12:00|1.4091206135396188|4|8066095787|147|0.6123098123133061|0|47|459|-80.732725|83|35.082768|IMPORT BEER|0.0|16|NEGRA MODELO 12PK BOTTLES|88adc9b2431567ae3a9d0afeec18f19f851e83a1|1.0450148292139363|0.61242566243833529|00080660957876|IMPORT BEER|BEER|-80.732725|1.409051865357139|147|1
35.082768|d847bdb0e29e687f36ae4bffbb93f3625d54337a|13.99|2015-01-10 18:30:00|1.4091206135396188|4|8066095787|147|0.6123098123133061|0|47|459|-80.732725|83|35.082768|IMPORT BEER|0.0|16|NEGRA MODELO 12PK BOTTLES|88adc9b2431567ae3a9d0afeec18f19f851e83a1|1.0450148292139363|0.61242566243833529|00080660957876|IMPORT BEER|BEER|-80.732725|1.409051865357139|147|1
35.082768|1d1237e291294c24a649cc239048b3a7cd8f8bee|2.57|2015-01-25 18:48:00|80.732732175546019|4|7203698634|147|35.097891752380185|0|35|425|-80.771677|72|35.066546|NFS-PAPER NAPKINS|0.0|1|YH NAPKINS 500 CT|88adc9b2431567ae3a9d0afeec18f19f851e83a1|1.0450148292139363|35.101032182271901|00072036986344|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.732725|80.732731382141537|45|1
35.082768|027b25e2dac0e279457b3f0c6993ef29d9d7aabf|2.57|2015-03-04 18:48:00|80.732732175546019|4|7203698634|147|35.097891752380185|0|35|425|-80.771677|72|35.066546|NFS-PAPER NAPKINS|0.0|1|YH NAPKINS 500 CT|88adc9b2431567ae3a9d0afeec18f19f851e83a1|1.0450148292139363|35.101032182271901|00072036986344|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.732725|80.732731382141537|45|1
35.082768|da1dfe5ea2acdf2f7c537932828a13d65b7aa208|2.35|2015-01-20 14:44:00|1.4091206135396188|4|4112907700|147|0.6123098123133061|0|47|1219|-80.732725|275|35.082768|PASTA SC CORE|0.0|1|CLASSICO SC SAUSAGE PEPPER ON|88adc9b2431567ae3a9d0afeec18f19f851e83a1|1.0450148292139363|0.61242566243833529|00041129077023|PASTA SAUCES|G1 GROCERY|-80.732725|1.409051865357139|147|1
35.082768|4d2c62773ba12932dd1e62ff2a04452dc1643050|0.85|2015-01-04 18:12:00|1.4091206135396188|4|7203636026|147|0.6123098123133061|0|47|54|-80.732725|8|35.082768|DIET|0.35|23|HT DIET TONIC WITH QUININE|88adc9b2431567ae3a9d0afeec18f19f851e83a1|1.0450148292139363|0.61242566243833529|00072036360410|CARBONATED BEVERAGES|BEVERAGE|-80.732725|1.409051865357139|147|1
35.082768|ba500ca64ad428c1be0053d4a491b8a0b5935720|1.7|2014-12-28 11:51:00|80.732732175546019|4|7203636026|147|35.09789175327596|0|35|54|-80.562829|8|35.006282|DIET|0.7|23|HT DIET TONIC WITH QUININE|88adc9b2431567ae3a9d0afeec18f19f851e83a1|1.0450148292139363|35.101032182271901|00072036360410|CARBONATED BEVERAGES|BEVERAGE|-80.732725|80.732725512795|60|2
35.082768|b9b2f384e7e4b3a68b5aac43610db5d4bd3fd989|1.7|2015-01-15 18:08:00|1.4091206135396188|4|7203636026|147|0.6123098123133061|0|47|54|-80.732725|8|35.082768|DIET|0.0|23|HT DIET TONIC WITH QUININE|88adc9b2431567ae3a9d0afeec18f19f851e83a1|1.0450148292139363|0.61242566243833529|00072036360410|CARBONATED BEVERAGES|BEVERAGE|-80.732725|1.409051865357139|147|2
35.140781|935ad3d93eabdb81c333f92bdb5c23a0bc5a9749|6.87|2014-12-07 12:06:00|1.4091206135396188|2|7225100105|39|0.6133223301722653|0|47|238|-80.62331|38|35.140781|RICE FLAVORED|1.87|1|NEAR EAST RICE PILAF|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00072251001051|RICE GRAINS AND BEANS|G1 GROCERY|-80.62331|1.4071422133560694|39|3
35.140781|dc4e403d0c585b49887ce07636c32c45be4799fd|131.88|2014-12-14 15:34:00|1.4091206135396188|2|8500001163|39|0.6133223301722653|0|47|9972|-80.62331|888|35.140781|NFS-U/PREM-CAB SAUVIGNON|0.0|13|LOUIS MARTINI CAB SAUV SONOMA|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00085000011638|ULTRA PREMIUM ($15-$19.99)|WINE|-80.62331|1.4071422133560694|39|12
35.140781|0749adfee2183e3687312b540ebc4c4596f2a0e9|21.98|2014-12-13 12:50:00|1.4091206135396188|2|8500001163|39|0.6133223301722653|0|47|9972|-80.62331|888|35.140781|NFS-U/PREM-CAB SAUVIGNON|0.0|13|LOUIS MARTINI CAB SAUV SONOMA|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00085000011638|ULTRA PREMIUM ($15-$19.99)|WINE|-80.62331|1.4071422133560694|39|2
35.140781|c5bc78b6e2a306c5799a885f4fd6e9ae26ec640d|12.99|2015-02-01 18:00:00|80.632521683083056|2|8500001163|39|35.153385273571423|0|39|9972|-80.709466|888|35.124987|NFS-U/PREM-CAB SAUVIGNON|0.0|13|LOUIS MARTINI CAB SAUV SONOMA|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|35.177497916598789|00085000011638|ULTRA PREMIUM ($15-$19.99)|WINE|-80.62331|80.623318564773399|157|1
35.140781|645844f147849197be66c8973bfd926f5141fc30|10.99|2014-10-06 18:31:00|1.4091206135396188|2|8500001163|39|0.6133223301722653|0|47|9972|-80.62331|888|35.140781|NFS-U/PREM-CAB SAUVIGNON|0.0|13|LOUIS MARTINI CAB SAUV SONOMA|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00085000011638|ULTRA PREMIUM ($15-$19.99)|WINE|-80.62331|1.4071422133560694|39|1
35.140781|9b6538826958377059783d4e141720099359fa5e|21.98|2014-10-03 18:27:00|80.632521683083056|2|8500001163|39|35.153385274882744|0|39|9972|-80.654118|888|35.123768|NFS-U/PREM-CAB SAUVIGNON|0.0|13|LOUIS MARTINI CAB SAUV SONOMA|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|35.177497916598789|00085000011638|ULTRA PREMIUM ($15-$19.99)|WINE|-80.62331|80.623314890179671|473|2
35.140781|4f3f749d0d44f168b925550537196f256d9ae8c9|12.99|2015-01-11 13:27:00|1.4091206135396188|2|8500001163|39|0.6133223301722653|0|47|9972|-80.62331|888|35.140781|NFS-U/PREM-CAB SAUVIGNON|0.0|13|LOUIS MARTINI CAB SAUV SONOMA|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00085000011638|ULTRA PREMIUM ($15-$19.99)|WINE|-80.62331|1.4071422133560694|39|1
35.140781|5a6ef95bd9fce77e382979d12a93a418a8bb5f2b|0.72|2014-12-31 14:07:00|80.632521683083056|2||39|35.153385274882744|0|39|502|-80.654118|64|35.123768|FRESH BANANAS|0.0|4|BANANAS, YELLOW|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|35.177497916598789|00204011000008|FRESH PRODUCE|PRODUCE|-80.62331|80.623314890179671|473|1
35.140781|e37e3fe5948ca1fc82ce7f669ee100a4269ec97e|0.7|2014-11-16 10:50:00|1.4091206135396188|2||39|0.6133223301722653|0|47|502|-80.62331|64|35.140781|FRESH BANANAS|0.0|4|BANANAS, YELLOW|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00204011000008|FRESH PRODUCE|PRODUCE|-80.62331|1.4071422133560694|39|1
35.140781|2d703a1ba8a0d22ee141bb48377754673aff31db|0.98|2014-10-23 17:56:00|80.632521683083056|2||39|35.153385274882744|0|39|502|-80.654118|64|35.123768|FRESH BANANAS|0.0|4|BANANAS, YELLOW|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|35.177497916598789|00204011000008|FRESH PRODUCE|PRODUCE|-80.62331|80.623314890179671|473|1
35.140781|4c06f40481613f70e663b7927073b57c821be084|3.99|2014-10-13 17:18:00|80.632521683083056|2|20405400000|39|35.153385274882744|0|39|504|-80.654118|64|35.123768|FRESH BERRIES|0.2|4|RED RASPBERRIES 6 OZ|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|35.177497916598789|00812049004402|FRESH PRODUCE|PRODUCE|-80.62331|80.623314890179671|473|1
35.140781|7fa3258f902efd36bf5eca81bc1153e01f665318|1.59|2014-09-21 10:31:00|1.4091206135396188|2|1090000383|39|0.6133223301722653|0|47|428|-80.62331|3|35.140781|NFS-BAKING CUPS|0.0|1|REYNOLDS FOIL BAKE CUPS|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00010900003834|BAKING SUPPLIES|G1 GROCERY|-80.62331|1.4071422133560694|39|1
35.140781|06bed06f57dd33ca9af91ee16064317a929f29c7|4.0|2014-09-14 18:12:00|1.4091206135396188|2|66440177739|39|0.6133223301722653|0|47|1165|-80.62331|87|35.140781|NFS-FRESH CONSUMER BUNCH|0.0|9|BUNCH- JUMBO SUNFLOWER 3 ST|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00664401777390|FLORAL|FLORAL|-80.62331|1.4071422133560694|39|1
35.140781|e003f994987fb5e268350d341bb16c8f7ba6c5ca|4.19|2014-10-02 19:55:00|80.632521683083056|2|4812127620|39|35.153385274882744|0|39|1037|-80.654118|164|35.123768|ENGLISH MUFFINS|0.0|7|THOMAS 100% WHEAT ENG MUFN PP|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|35.177497916598789|00048121184070|BREAKFAST|COMMERCIAL BAKERY|-80.62331|80.623314890179671|473|1
35.140781|470fc8f116175f736fce0d60b1a7f5810652dfef|3.49|2014-11-08 17:45:00|1.4091206135396188|2|4812127620|39|0.6133223301722653|0|47|1037|-80.62331|164|35.140781|ENGLISH MUFFINS|1.75|7|THOMAS 100% WHEAT ENG MUFN PP|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00048121184070|BREAKFAST|COMMERCIAL BAKERY|-80.62331|1.4071422133560694|39|1
35.140781|3b62a3cf3523d84d9e2b19aa6ca0df6812aa7d11|4.49|2015-01-18 17:23:00|80.632521683083056|2|2840009217|39|35.153385274882744|0|39|1981|-80.654118|480|35.123768|CHIPS|0.0|6|STACY'S PITA CHIPS NAKED|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|35.177497916598789|00028400092173|DRY GOODS|DELI|-80.62331|80.623314890179671|473|1
35.140781|42e4a9de3baa43d967252176cf2f643bca37ea90|5.25|2014-11-08 11:09:00|1.4091206135396188|2|7203633086|39|0.6133223301722653|0|47|1148|-80.62331|21|35.140781|ALMONDS|1.75|1|HT ROASTED ALMONDS LIGHT SALT|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00072036979537|NUTS|G1 GROCERY|-80.62331|1.4071422133560694|39|1
35.140781|a0d616e9b761630caddcf072fb18cf42d1a8edff|6.99|2014-11-03 18:22:00|1.4091206135396188|2|8143450009|39|0.6133223301722653|0|47|9948|-80.62331|886|35.140781|NFS-PREM-CAB SAUVIGNON|0.0|13|BLACKSTONE CAB SAUV|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00081434500090|PREMIUM ($8-$10.99)|WINE|-80.62331|1.4071422133560694|39|1
35.140781|437fd4582661c140b679f75853e2714c459bdbe1|6.99|2015-01-20 16:44:00|80.632521683083056|2|8143450009|39|35.153385274882744|0|39|9948|-80.654118|886|35.123768|NFS-PREM-CAB SAUVIGNON|0.0|13|BLACKSTONE CAB SAUV|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|35.177497916598789|00081434500090|PREMIUM ($8-$10.99)|WINE|-80.62331|80.623314890179671|473|1
35.140781|c49eb637617da1aa4339c403de6039c3d318e32f|13.98|2014-10-31 21:18:00|1.4091206135396188|2|8143450009|39|0.6133223301722653|0|47|9948|-80.62331|886|35.140781|NFS-PREM-CAB SAUVIGNON|0.0|13|BLACKSTONE CAB SAUV|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00081434500090|PREMIUM ($8-$10.99)|WINE|-80.62331|1.4071422133560694|39|2
35.140781|fafa1cb2154fcfae0f80bc8e4bf807bb3ba1211c|0.99|2015-02-06 13:09:00|1.4091206135396188|2|7252104965|39|0.6133223301722653|0|47|30|-80.62331|4|35.140781|CARBONATED WATER|0.0|1|VINTAGE SELTZER RASPBERRY 1LT|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00072521049769|BOTTLED WATER|G1 GROCERY|-80.62331|1.4071422133560694|39|1
35.140781|5173d77202ed62cb8d80047952bc198c8c201162|9.98|2014-12-20 10:23:00|1.4091206135396188|2|4650062248|39|0.6133223301722653|0|47|422|-80.62331|71|35.140781|NFS-REMAIN LAUNDRY SUPPL|0.0|1|SHOUT COLOR CATCHER|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00046500622489|LAUNDRY SUPPLIES|G1 GROCERY|-80.62331|1.4071422133560694|39|2
35.140781|63ec93300ed301a78bdb3826289dca9e2ae95c43|3.59|2014-11-02 11:54:00|80.632521683083056|2|5210004780|39|35.153385274882744|0|39|18|-80.654118|3|35.123768|CAKE DECORATIONS & ICING|1.59|1|MC RED ICING|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|35.177497916598789|00052100048406|BAKING SUPPLIES|G1 GROCERY|-80.62331|80.623314890179671|473|1
35.140781|3c346eaf577e801df4481b8b01b54ab7835bc880|3.99|2014-09-26 17:59:00|1.4091206135396188|2|4525511880|39|0.6133223301722653|0|47|523|-80.62331|64|35.140781|FRESH POTATOES|0.0|4|DUTCH YELLOW POTATO 24 OZ|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00045255118803|FRESH PRODUCE|PRODUCE|-80.62331|1.4071422133560694|39|1
35.140781|d4d72b3d7c813d2483580212ac579b4a4220b985|1.79|2015-02-28 20:22:00|1.4091206135396188|2|3660082801|39|0.6133223301722653|0|47|4237|-80.62331|1200|35.140781|MEDICATED LIP CARE|0.0|17|(PPL)CHAP STICK MST BALM|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00036600828010|COUGH/COLD/SINUS|HBC|-80.62331|1.4071422133560694|39|1
35.140781|4ea39eb5c0f153d9bb8113f3effba617415ec619|3.78|2015-02-09 14:33:00|80.632521683083056|2|5480003077|39|35.153385274882744|0|39|138|-80.654118|38|35.123768|RICE MICROWAVE|0.0|1|UNCLE BEN RR JASMINE|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|35.177497916598789|00054800344468|RICE GRAINS AND BEANS|G1 GROCERY|-80.62331|80.623314890179671|473|2
35.140781|b068201488fb8f870644e09bef8e34e1e3b2d6e2|1.57|2014-09-28 17:45:00|1.4091206135396188|2|7009030410|39|0.6133223301722653|0|47|225|-80.62331|35|35.140781|SUGAR-GRANULATED|0.07|1|CRYSTAL FINE GRANULATED SUGAR|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00070090304104|SUGAR/SUBSTITUTES|G1 GROCERY|-80.62331|1.4071422133560694|39|1
35.140781|04142fabfa0ff53293210f8258cc0a165a9587d1|1.99|2015-01-12 18:43:00|1.4091206135396188|2|7203670829|39|0.6133223301722653|0|47|257|-80.62331|39|35.140781|TOMATOES|0.0|1|HTT TOMATO PLUM CRUSHED|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00072036708298|VEGETABLES-CAN/JAR|G1 GROCERY|-80.62331|1.4071422133560694|39|1
35.140781|be0c8fe856589a80a6011f6323f0b063f1818979|5.99|2014-09-10 16:47:00|1.4091206135396188|2|1834175101|39|0.6133223301722653|0|47|9935|-80.62331|885|35.140781|NFS POP CAB SAUV|0.0|13|BAREFOOT CAB SAUV|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00018341751017|POPULAR (4-$7.99)|WINE|-80.62331|1.4071422133560694|39|1
35.140781|14d5e194aea5985a84c58f642d5c61d7442060bf|5.79|2015-02-28 10:22:00|80.632521683083056|2|7007480240|39|35.153385274882744|0|39|3|-80.654118|1|35.123768|FORMULA RTF|0.0|1|PEDIALYTE GRAPE FLAVOR|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|35.177497916598789|00070074802404|BABY FOOD|G1 GROCERY|-80.62331|80.623314890179671|473|1
35.140781|2c471bbb6c73d4fcfaac2812d0e2e32d815ed28f|3.59|2015-01-24 18:14:00|1.4091206135396188|2|7341016305|39|0.6133223301722653|0|47|1035|-80.62331|163|35.140781|SANDWICH ROLL|0.0|7|ARN SELECT 100% WHEAT HAMS PP|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00073410161456|BUNS/ROLLS|COMMERCIAL BAKERY|-80.62331|1.4071422133560694|39|1
35.140781|445716105d96dabd3f5ed417226f95d3cfd01ce3|7.99|2014-11-09 17:11:00|80.632521683083056|2|20639500000|39|35.153385274882744|0|39|1654|-80.654118|381|35.123768|DESSERT CAKES|0.0|14|CHOCOLATE PATTI CAKE 2 LAYER|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|35.177497916598789|00206395000001|CAKES|BAKERY|-80.62331|80.623314890179671|473|1
35.140781|fc6bd689a390111d4d29681c51dcadbfac959601|12.99|2014-10-08 19:29:00|1.4091206135396188|2|8769201103|39|0.6133223301722653|0|47|458|-80.62331|82|35.140781|CRAFT BEER|0.0|16|SAM ADAMS SEASONAL 12PK|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00087692011033|DOMESTIC BEER|BEER|-80.62331|1.4071422133560694|39|1
35.140781|4570ab44bc10d0ca5d5ccbe4bd7d1ec431f623ad|19.98|2015-02-05 20:34:00|80.632521683083056|2|84715900080|39|35.153385274882744|0|39|9972|-80.654118|888|35.123768|NFS-U/PREM-CAB SAUVIGNON|0.0|13|CONTEMPO CABERNET|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|35.177497916598789|00847159000808|ULTRA PREMIUM ($15-$19.99)|WINE|-80.62331|80.623314890179671|473|2
35.140781|95c6b61a05af353b56cf500fc4cd96406c9c61e0|6.99|2014-10-24 20:00:00|1.4091206135396188|2|1820002992|39|0.6133223301722653|0|47|465|-80.62331|85|35.140781|NON ALCOHOLIC|0.0|16|O'DOULS  AMBER NA 6PK 12OZ BTL|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00018200029929|NON ALCOHOLIC|BEER|-80.62331|1.4071422133560694|39|1
35.140781|1377550565c98d5337d06c64c5e86c494282b9b2|4.29|2014-09-24 13:19:00|1.4091206135396188|2|3450015119|39|0.6133223301722653|0|47|312|-80.62331|51|35.140781|BUTTER|0.0|3|LOL LT BUTTER W CANOLA OIL|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00034500151849|BUTTER & MARGARINE|DAIRY|-80.62331|1.4071422133560694|39|1
35.140781|bb9fb2eb7d9c6252aa95e39a77894ad514fe60aa|9.99|2014-11-16 20:49:00|80.632521683083056|2|89875600105|39|35.153385274882744|0|39|9948|-80.654118|886|35.123768|NFS-PREM-CAB SAUVIGNON|0.0|13|LINE 39 CABERNET SAUVIGNON|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|35.177497916598789|00898756001057|PREMIUM ($8-$10.99)|WINE|-80.62331|80.623314890179671|473|1
35.140781|35115dc894ba7b715e431ef1649f91788f2a46fd|2.69|2014-09-16 18:07:00|1.4091206135396188|2|7203663996|39|0.6133223301722653|0|47|342|-80.62331|57|35.140781|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00072036631299|MILK|DAIRY|-80.62331|1.4071422133560694|39|1
35.140781|a2beb72eb7d44aad17826e9d694769da675d6b45|2.79|2014-09-20 11:29:00|1.4091206135396188|2|2100064353|39|0.6133223301722653|0|47|184|-80.62331|28|35.140781|SALAD DRESSINGS-LIQUID|0.0|1|KRAFT DRS ITALIAN CREAMY|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00021000644261|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.62331|1.4071422133560694|39|1
35.140781|b5cfbf49c99c0399b5d020450f4a4fdffe218358|1.69|2014-12-20 13:02:00|1.4091206135396188|2|4900000044|39|0.6133223301722653|0|47|54|-80.62331|8|35.140781|DIET|0.0|23|CB DIET COKE CONTOUR 20 OZ NR|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00049000000450|CARBONATED BEVERAGES|BEVERAGE|-80.62331|1.4071422133560694|39|1
35.140781|f471806003a5493fea1a339e9401bfab452647e8|1.69|2014-11-12 14:58:00|80.632521683083056|2|4900000044|39|35.153385274882744|0|39|54|-80.654118|8|35.123768|DIET|0.0|23|CB DIET COKE CONTOUR 20 OZ NR|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|35.177497916598789|00049000000450|CARBONATED BEVERAGES|BEVERAGE|-80.62331|80.623314890179671|473|1
35.140781|96559a89bee3a75dd09d69a7de5a1e23d68bbc74|7.99|2014-11-06 18:27:00|1.4091206135396188|2|71280812982|39|0.6133223301722653|0|47|458|-80.62331|82|35.140781|CRAFT BEER|0.0|16|HIGHLAND GAELIC ALE 6PK|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|0.61242566243833529|00712808129820|DOMESTIC BEER|BEER|-80.62331|1.4071422133560694|39|1
35.140781|aa463fc8ed99301020366c52d830673fb2aadcda|3.0|2014-11-02 11:59:00|80.632521683083056|2|7203632021|39|35.153385274882744|0|39|195|-80.654118|30|35.123768|SALAD & COOKING OIL|0.0|1|HT VEGETABLE OIL|8edb490a515b3f5ac535c0386d71709c88f05a50|0.870924999989006|35.177497916598789|00072036320216|SHORTENING/OIL|G1 GROCERY|-80.62331|80.623314890179671|473|1
35.43259|53e10bd6bcaf5423bce3057cdd75ddc3406f95dc|9.99|2015-03-07 09:27:00|80.607132136635443|4|7707117210|202|35.464446622370005|0|9|7185|-80.860108|1600|35.500972|SOFTSIDE COOLERS|0.5|18|HT FOAM COOLER|9085061e409edee3c547b3ce35e831d6f843e4de|2.2012158986689503|35.47365851958088|00077071172103|SEASONAL MERCHANDISE|GM|-80.605588|80.605605637492374|268|1
35.43259|65ca860c8ebdcf929c5d91a170a608f5dece43f0|2.4|2015-01-22 19:59:00|1.4057311447477159|4|3663203732|202|0.6184153580092175|0|52|685|-80.605588|61|35.43259|GREEK|0.0|3|DANNON LNF GREEK CHOC CHERRY|9085061e409edee3c547b3ce35e831d6f843e4de|2.2012158986689503|0.6209993146566879|00036632037503|YOGURT|DAIRY|-80.605588|1.406832906106031|202|2
35.43259|c852e003c1d2f3a55c5d2d3fbec49b272d41bce5|9.99|2015-01-15 20:46:00|1.4057311447477159|4|978055359369|202|0.6184153580092175|0|52|6777|-80.605588|1566|35.43259|PAPER BACK BOOKS|0.0|18|INNOCENCE A NOVEL|9085061e409edee3c547b3ce35e831d6f843e4de|2.2012158986689503|0.6209993146566879|09780553593693|BOOKS|GM|-80.605588|1.406832906106031|202|1
35.43259|e0319c69ab0d562f1ce1dc7c060db170cc0ce6c8|2.19|2014-10-04 21:31:00|1.4057311447477159|4|1200000496|202|0.6184153580092175|0|52|54|-80.605588|8|35.43259|DIET|0.69|23|DIET PEPSI 2 LTR NR|9085061e409edee3c547b3ce35e831d6f843e4de|2.2012158986689503|0.6209993146566879|00012000002311|CARBONATED BEVERAGES|BEVERAGE|-80.605588|1.406832906106031|202|1
35.43259|0da3d0849804a4757136713711293368957307f8|3.29|2015-02-24 14:53:00|1.4057311447477159|4|2840011895|202|0.6184153580092175|0|52|204|-80.605588|31|35.43259|TORTILLA CHIPS|0.0|1|TOSTITOS CANTINA TRADITIONAL|9085061e409edee3c547b3ce35e831d6f843e4de|2.2012158986689503|0.6209993146566879|00028400118958|SNACKS|G1 GROCERY|-80.605588|1.406832906106031|202|1
35.006282|ec611fa8486c3321042814eac4c80fee6526ffed|7.69|2014-10-20 17:46:00|80.562862110758871|4|8087800550|60|35.124799495117799|0|21|3503|-80.64817|1045|35.04711|CONDITIONER-PREMIUM|1.69|17|PANTENE CND DLY MOIS RENEWAL|9295dafccec855564b4746b009ec9a32508d18cb|8.189272709394746|35.054042368968126|00080878171316|HAIR & SCALP CARE|HBC|-80.562829|80.562834660794422|129|1
35.053394|1479f5df44346c8bc2229a3c9e48f40686986c7a|11.99|2015-02-23 21:12:00|80.848351720559364|2|3700088206|11|35.082757871906274|0|25|426|-80.806073|72|35.106477|NFS-PAPER TOWELS|2.0|1|BOUNTY TOWEL 6 RL SAS WHITE|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00037000882022|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.848528|80.848554714125086|4|1
35.053394|1e94877cf6df8eda7c9f704117a71d84fc0a4f23|2.99|2014-10-20 11:58:00|80.848351720559364|2|3700000309|11|35.082757871906274|0|25|4070|-80.806073|1080|35.106477|TOOTHPASTE-BAKING SODA|0.5|17|CREST BAKING SODA& PER-32024|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00037000320241|ORAL HYGIENE|HBC|-80.848528|80.848554714125086|4|1
35.053394|ff14961fc2e945f2b70517a2178d7074be974d01|1.5|2014-10-28 12:54:00|80.848351720559364|2|3663201937|11|35.082757871906274|0|25|685|-80.806073|61|35.106477|GREEK|0.5|3|DANNON INDUL CHOC RSPBRY TRUFL|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00036632019363|YOGURT|DAIRY|-80.848528|80.848554714125086|4|1
35.053394|10d9520ba52f848fa854ea4ac4f3defa76c24099|18.99|2015-01-18 13:03:00|80.848351720559364|2|3700088207|11|35.082757879379905|0|25|426|-80.816172|72|35.059823|NFS-PAPER TOWELS|8.02|1|BOUNTY TOWEL 12 WHITE|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00037000882077|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.848528|80.848535645294604|66|1
35.053394|120b78da40fb67039375e9d9c1d43ea0066ba0e0|8.99|2014-09-29 13:31:00|80.848351720559364|2|3760048620|11|35.082757872007456|0|25|358|-80.78468|100|35.096737|REGULAR BACON|4.0|19|HORMEL BLACK LABEL LOW SALT|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00037600486200|BACON|CASE READY MEATS|-80.848528|80.848554547573357|30|1
35.053394|16db4e884fc0c7ea00ebaff99f2e7ffcd1ff46e3|5.49|2015-03-02 10:02:00|80.848351720559364|2|3700080070|11|35.082757872007456|0|25|417|-80.78468|71|35.096737|NFS-FABRIC SOFTENERS|0.5|1|BOUNCE FRESH LINEN SHEETS 80CT|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00037000800699|LAUNDRY SUPPLIES|G1 GROCERY|-80.848528|80.848554547573357|30|1
35.053394|06e650362534b56cbb7f11478963d356a36a5bba|18.99|2014-12-17 09:56:00|80.848351720559364|2|3700088207|11|35.082757871906274|0|25|426|-80.806073|72|35.106477|NFS-PAPER TOWELS|3.0|1|BOUNTY TOWEL 12 WHITE|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00037000882077|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.848528|80.848554714125086|4|1
35.053394|861bc04272bdd5f4ef3f87fb0216ea9553d28985|3.29|2014-09-26 13:29:00|80.848351720559364|2|5210000444|11|35.082757872007456|0|25|1245|-80.78468|34|35.096737|SINGLE SPICES|0.0|1|E  MC CINNAMON SUGAR|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00052100004440|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.848528|80.848554547573357|30|1
35.053394|e0891e159ac943eb5192aaae17cfc0fb48dab6b6|6.99|2015-02-05 14:54:00|80.848351720559364|2|7703401130|11|35.082757871906274|0|25|141|-80.806073|21|35.106477|TRAIL MIXES AND BLENDS|0.0|1|SECOND NATURE CALIFORNIA MEDLY|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00077034011487|NUTS|G1 GROCERY|-80.848528|80.848554714125086|4|1
35.053394|0217c2d76cb97528165975bd477a879570cc14a6|6.99|2015-02-14 12:26:00|80.848351720559364|2|7703401130|11|35.082757852291103|0|25|141|-80.709466|21|35.124987|TRAIL MIXES AND BLENDS|0.0|1|SECOND NATURE CALIFORNIA MEDLY|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00077034011487|NUTS|G1 GROCERY|-80.848528|80.848577328019871|157|1
35.053394|9be3fae0362cbecbae5d182baf607bbc98f4c1a1|12.98|2014-12-11 12:39:00|80.848351720559364|2|7703401130|11|35.082757871906274|0|25|141|-80.806073|21|35.106477|TRAIL MIXES AND BLENDS|1.5|1|SECOND NATURE CALIFORNIA MEDLY|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00077034011487|NUTS|G1 GROCERY|-80.848528|80.848554714125086|4|2
35.053394|8007575fb7b1666b3a4f75c0654e8ada4175541b|6.49|2014-12-04 13:08:00|80.848351720559364|2|7703401130|11|35.082757879379905|0|25|141|-80.816172|21|35.059823|TRAIL MIXES AND BLENDS|0.0|1|SECOND NATURE CALIFORNIA MEDLY|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00077034011487|NUTS|G1 GROCERY|-80.848528|80.848535645294604|66|1
35.053394|8ae0bd956dcf48422f85a5967df66399e0bef5b4|6.99|2015-03-04 16:22:00|80.848351720559364|2|7703401130|11|35.082757879379905|0|25|141|-80.816172|21|35.059823|TRAIL MIXES AND BLENDS|0.0|1|SECOND NATURE CALIFORNIA MEDLY|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00077034011487|NUTS|G1 GROCERY|-80.848528|80.848535645294604|66|1
35.053394|b0d53f36163f404dcc701858e410c36034e60605|6.49|2014-12-24 17:16:00|80.848351720559364|2|7703401130|11|35.082757871906274|0|25|141|-80.806073|21|35.106477|TRAIL MIXES AND BLENDS|0.7|1|SECOND NATURE CALIFORNIA MEDLY|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00077034011487|NUTS|G1 GROCERY|-80.848528|80.848554714125086|4|1
35.053394|7f8863ba48e15089838d4bfd64f78f4bc4343625|6.99|2015-02-18 16:07:00|80.848351720559364|2|7703401130|11|35.082757852291103|0|25|141|-80.709466|21|35.124987|TRAIL MIXES AND BLENDS|1.5|1|SECOND NATURE CALIFORNIA MEDLY|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00077034011487|NUTS|G1 GROCERY|-80.848528|80.848577328019871|157|1
35.053394|c14c6cbb67ad5c63d3178b09fa6eba39e6719c91|6.49|2014-11-17 19:26:00|80.848351720559364|2|7703401130|11|35.082757852291103|0|25|141|-80.709466|21|35.124987|TRAIL MIXES AND BLENDS|0.0|1|SECOND NATURE CALIFORNIA MEDLY|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00077034011487|NUTS|G1 GROCERY|-80.848528|80.848577328019871|157|1
35.053394|821fa81cce82f86ddca098df90563e5b029a500d|8.58|2014-09-17 14:07:00|80.848351720559364|2|7341001375|11|35.082757874444468|0|25|1027|-80.85753|162|35.116638|GRAIN|2.15|7|ARN HEALTHNUT BRD WP PP|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00073410013656|SLICED BREAD|COMMERCIAL BAKERY|-80.848528|80.848550161395963|204|2
35.053394|2844db25336404c79c9ae612432541a3c29f81e1|6.49|2014-12-29 18:39:00|80.848351720559364|2|7703401130|11|35.082757852291103|0|25|141|-80.709466|21|35.124987|TRAIL MIXES AND BLENDS|0.0|1|SECOND NATURE CALIFORNIA MEDLY|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00077034011487|NUTS|G1 GROCERY|-80.848528|80.848577328019871|157|1
35.053394|a5e126ccb429074a7b811b27cc73b095a6494487|6.99|2015-01-26 17:02:00|80.848351720559364|2|7703401130|11|35.082757852291103|0|25|141|-80.709466|21|35.124987|TRAIL MIXES AND BLENDS|0.0|1|SECOND NATURE CALIFORNIA MEDLY|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00077034011487|NUTS|G1 GROCERY|-80.848528|80.848577328019871|157|1
35.053394|9c0eb9a5afd36ca5dfdcb10581ddb645bba00e3c|3.99|2014-11-20 18:58:00|80.848351720559364|2|7341001375|11|35.082757852291103|0|25|1027|-80.709466|162|35.124987|GRAIN|2.0|7|ARN HEALTHNUT BRD WP PP|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00073410013656|SLICED BREAD|COMMERCIAL BAKERY|-80.848528|80.848577328019871|157|1
35.053394|dff0c76004f1d57ec6c870ace9caee13cbdb41e1|6.49|2015-01-05 14:50:00|80.848351720559364|2|7703401130|11|35.082757871906274|0|25|141|-80.806073|21|35.106477|TRAIL MIXES AND BLENDS|0.0|1|SECOND NATURE CALIFORNIA MEDLY|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00077034011487|NUTS|G1 GROCERY|-80.848528|80.848554714125086|4|1
35.053394|025665199f3fda2407626abe3445244350e1efee|1.69|2014-12-01 12:00:00|80.848351720559364|2||11|35.082757872007456|0|25|524|-80.78468|64|35.096737|FRESH PROD FRESH ONIONS|0.5|4|COO SWEET ONIONS|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00204159000007|FRESH PRODUCE|PRODUCE|-80.848528|80.848554547573357|30|1
35.053394|0879897570cb783be2c8048862cc6d61809f4aa5|1.67|2014-10-07 13:08:00|80.848351720559364|2|76101040154|11|35.082757871906274|0|25|511|-80.806073|64|35.106477|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS 2 CT BAG|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00761010401545|FRESH PRODUCE|PRODUCE|-80.848528|80.848554714125086|4|1
35.053394|7b086ce23073074b184f436dbb1477d942438079|1.79|2014-11-11 22:49:00|80.848351720559364|2|1800000261|11|35.082757852291103|0|25|325|-80.709466|54|35.124987|BISCUITS-REFRIGERATED|0.0|3|GRANDS BUTTERMILK BISCUITS|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00018000001873|DOUGH PRODUCTS|DAIRY|-80.848528|80.848577328019871|157|1
35.053394|e13e575023f57c8b32ddf6e13d5407f7c979ddca|2.89|2014-09-12 15:02:00|80.848351720559364|2|3800040260|11|35.082757871906274|0|25|1269|-80.806073|41|35.106477|BREAKFAST SYRUP CARRIER|0.0|5|EGGO HOMESTYLE WAFFLES|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00038000402609|BREAKFAST FOODS FROZEN|FROZEN|-80.848528|80.848554714125086|4|1
35.053394|1229d349d9f101a09dab061d157698afbe08a1b0|3.99|2014-10-06 10:38:00|80.848351720559364|2|2500005542|11|35.082757872007456|0|25|335|-80.78468|56|35.096737|ORANGE JUICE-REGRIGERATED|0.99|3|SIMPLY ORANGE GROVE MADE|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00025000055447|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.848528|80.848554547573357|30|1
35.053394|2cd9717c7cd9adafcd4eec516e5193b5a0e6e88e|3.79|2014-09-15 17:55:00|80.848351720559364|2|2500005542|11|35.082757871906274|0|25|335|-80.806073|56|35.106477|ORANGE JUICE-REGRIGERATED|0.0|3|SIMPLY ORANGE GROVE MADE|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00025000055447|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.848528|80.848554714125086|4|1
35.053394|180dbb71782d0618fa406dae48eebc1ae14c0fe1|2.99|2014-09-20 20:58:00|80.848351720559364|2|20789700000|11|35.082757871906274|0|25|1677|-80.806073|383|35.106477|INDIVIDUALS (PASTRY CASE)|0.0|14|MEGA RED VELVET CUPCAKE|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00207897000001|PASTRY CASE|BAKERY|-80.848528|80.848554714125086|4|1
35.053394|7e67950ef530127eab9ec0c9dd398c8f32853433|3.69|2015-02-02 12:58:00|80.848351720559364|2|68833992319|11|35.082757871906274|0|25|1611|-80.806073|371|35.106477|PITA'S AND FLAT BREADS|0.0|14|TRADITIONAL WHITE FOLDIT|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00688339924336|BREAD|BAKERY|-80.848528|80.848554714125086|4|1
35.053394|94828b9fb124393d325370bac40fba9178ac6689|2.99|2015-01-10 21:03:00|80.848351720559364|2|3000004760|11|35.082757872007456|0|25|60|-80.78468|9|35.096737|HOT CEREAL|0.0|1|QUAKER INST GRITS ORIGINAL|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00030000047606|CEREAL|G1 GROCERY|-80.848528|80.848554547573357|30|1
35.053394|ca4b9c9650b44fdde2b865204bd7b10384817fcc|3.49|2014-10-13 22:47:00|80.848351720559364|2|3000001190|11|35.082757852291103|0|25|60|-80.709466|9|35.124987|HOT CEREAL|0.99|1|QUAKER OATML RSN DATE WALNT|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00030000012406|CEREAL|G1 GROCERY|-80.848528|80.848577328019871|157|1
35.053394|9835cd2abca6df34ba5ef5cd9b1f53bbe57d1077|3.89|2014-09-11 12:51:00|80.848351720559364|2|5150014110|11|35.082757871906274|0|25|126|-80.806073|19|35.106477|PRESERVES/MARMALADE|0.9|1|SMUCK ORCH FINEST CHERRY PRES|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00051500141137|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.848528|80.848554714125086|4|1
35.053394|cb70e7e434a6c50f1d453dfcd4f0fd43aaf489f2|2.99|2014-10-27 18:26:00|80.848351720559364|2|7073400003|11|35.082757871906274|0|25|230|-80.806073|37|35.106477|HERBAL TEA|0.49|1|CELESTIAL SLEEPYTIME|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00070734000034|TEA|G1 GROCERY|-80.848528|80.848554714125086|4|1
35.053394|a2e3e286208630e6b418698dd2a442310d40a371|4.99|2015-01-24 19:20:00|80.848351720559364|2|6827493471|11|35.082757872007456|0|25|31|-80.78468|4|35.096737|NON CARBONATED WATER|0.0|1|NESTLE PURE LIFE .5L 24PK|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00068274934711|BOTTLED WATER|G1 GROCERY|-80.848528|80.848554547573357|30|1
35.053394|3ba48b8003134177be2d7c23fd1b85227bce40cb|4.99|2015-03-08 21:15:00|80.848351720559364|2|6827493471|11|35.082757872007456|0|25|31|-80.78468|4|35.096737|NON CARBONATED WATER|1.0|1|NESTLE PURE LIFE .5L 24PK|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00068274934711|BOTTLED WATER|G1 GROCERY|-80.848528|80.848554547573357|30|1
35.053394|d9f8c69e646a11550b4debb146b263dedd704e5a|4.99|2014-12-18 12:16:00|80.848351720559364|2|6827493471|11|35.082757852291103|0|25|31|-80.709466|4|35.124987|NON CARBONATED WATER|1.2|1|NESTLE PURE LIFE .5L 24PK|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00068274934711|BOTTLED WATER|G1 GROCERY|-80.848528|80.848577328019871|157|1
35.053394|bbcc0504ff9dee189c02bffd9c729767617d978c|4.99|2015-02-10 22:39:00|80.848351720559364|2|6827493471|11|35.082757872007456|0|25|31|-80.78468|4|35.096737|NON CARBONATED WATER|2.0|1|NESTLE PURE LIFE .5L 24PK|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00068274934711|BOTTLED WATER|G1 GROCERY|-80.848528|80.848554547573357|30|1
35.053394|103edd3ae11698571af59cf4fb224700cca7bf58|14.7|2014-12-20 14:32:00|80.848351720559364|2|4470002268|11|35.082757871906274|0|25|358|-80.806073|100|35.106477|REGULAR BACON|3.68|19|OSCAR MAYER LOW SALT BACON|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00044700019917|BACON|CASE READY MEATS|-80.848528|80.848554714125086|4|2
35.053394|579bb35eaa538020e3d18bb3b1b51b2c48785a55|14.7|2015-01-07 11:52:00|80.848351720559364|2|4470002268|11|35.082757871906274|0|25|358|-80.806073|100|35.106477|REGULAR BACON|3.67|19|OSCAR MAYER LOW SALT BACON|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00044700019917|BACON|CASE READY MEATS|-80.848528|80.848554714125086|4|2
35.053394|f2ac6c1c1d5cfbbdecb4ee0bceba15288680b10c|5.99|2014-11-21 21:13:00|80.848351720559364|2|3700012880|11|35.082757871906274|0|25|389|-80.806073|66|35.106477|NFS-LAUNDRY DETERGENTS|0.0|1|IVORY SNOW GENTLE CARE 25OZ|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00037000128809|DETERGENTS|G1 GROCERY|-80.848528|80.848554714125086|4|1
35.053394|0846fb708ba756b97207d0d9e9a2efbd5080f7c0|0.91|2015-01-21 19:28:00|80.848351720559364|2||11|35.082757852291103|0|25|502|-80.709466|64|35.124987|FRESH BANANAS|0.0|4|BANANAS, YELLOW|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00204011000008|FRESH PRODUCE|PRODUCE|-80.848528|80.848577328019871|157|1
35.053394|6ceff966be0e82350dc0ffcb68ea502ba7bd439d|2.09|2014-10-23 20:53:00|80.848351720559364|2||11|35.082757879379905|0|25|502|-80.816172|64|35.059823|FRESH BANANAS|0.0|4|BANANAS, YELLOW|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00204011000008|FRESH PRODUCE|PRODUCE|-80.848528|80.848535645294604|66|1
35.053394|1c54e2c573ae6d89b9385e0b6cbe97294900c279|1.49|2015-02-25 19:37:00|80.848351720559364|2||11|35.082757871906274|0|25|502|-80.806073|64|35.106477|FRESH BANANAS|0.0|4|BANANAS, YELLOW|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00204011000008|FRESH PRODUCE|PRODUCE|-80.848528|80.848554714125086|4|1
35.053394|65b9475fcffe989713db27283e89608c1de8440f|1.31|2014-12-05 12:56:00|80.848351720559364|2||11|35.082757871906274|0|25|502|-80.806073|64|35.106477|FRESH BANANAS|0.0|4|BANANAS, YELLOW|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00204011000008|FRESH PRODUCE|PRODUCE|-80.848528|80.848554714125086|4|1
35.053394|7b3a6ad744999fe41b27425b9ec522caa3221e39|1.64|2014-11-24 13:17:00|80.848351720559364|2||11|35.082757871906274|0|25|502|-80.806073|64|35.106477|FRESH BANANAS|0.0|4|BANANAS, YELLOW|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00204011000008|FRESH PRODUCE|PRODUCE|-80.848528|80.848554714125086|4|1
35.053394|9c86abe5b0bccd4738cc245d8a329b64651f37b8|1.11|2014-11-15 20:30:00|80.848351720559364|2||11|35.082757871906274|0|25|502|-80.806073|64|35.106477|FRESH BANANAS|0.0|4|BANANAS, YELLOW|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00204011000008|FRESH PRODUCE|PRODUCE|-80.848528|80.848554714125086|4|1
35.053394|45c2448a5481c124898f94d3050494c80b4bc136|1.3|2014-12-10 14:30:00|80.848351720559364|2||11|35.082757871906274|0|25|502|-80.806073|64|35.106477|FRESH BANANAS|0.0|4|BANANAS, YELLOW|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00204011000008|FRESH PRODUCE|PRODUCE|-80.848528|80.848554714125086|4|1
35.053394|def3cf4900599cc1b1bb1739e4acaec622bdd149|1.31|2014-09-30 18:32:00|80.848351720559364|2||11|35.082757872007456|0|25|502|-80.78468|64|35.096737|FRESH BANANAS|0.0|4|BANANAS, YELLOW|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00204011000008|FRESH PRODUCE|PRODUCE|-80.848528|80.848554547573357|30|1
35.053394|093ba377d86b559c224545ec60229575b479c393|3.14|2014-09-25 12:59:00|80.848351720559364|2|7009030410|11|35.082757874444468|0|25|225|-80.85753|35|35.116638|SUGAR-GRANULATED|0.07|1|CRYSTAL FINE GRANULATED SUGAR|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00070090304104|SUGAR/SUBSTITUTES|G1 GROCERY|-80.848528|80.848550161395963|204|2
35.053394|1cd55a8dd91b0411b35f5c9fe426bbda01ee5bca|1.49|2014-12-19 14:15:00|80.848351720559364|2|7203653022|11|35.082757874444468|0|25|1273|-80.85753|50|35.116638|BAG VEG NON STEAM|0.0|5|HT CUT OKRA|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00072036537522|VEGETABLES-FROZEN|FROZEN|-80.848528|80.848550161395963|204|1
35.053394|8539f1539cd20f3aa3445c561aa04c628a55940b|0.99|2014-09-10 14:18:00|80.848351720559364|2|7203653022|11|35.082757874444468|0|25|1273|-80.85753|50|35.116638|BAG VEG NON STEAM|0.0|5|HT CUT OKRA|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00072036537522|VEGETABLES-FROZEN|FROZEN|-80.848528|80.848550161395963|204|1
35.053394|8b4d45d35f04c9d52acd7aeb6b2611aa1c74806d|3.38|2015-02-05 20:06:00|80.848351720559364|2|3660207290|11|35.082757852291103|0|25|4207|-80.709466|1200|35.124987|COUGH DROP-ADULT|0.84|17|RICOLA NATURAL HERB -07917|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00036602079175|COUGH/COLD/SINUS|HBC|-80.848528|80.848577328019871|157|2
35.053394|1fb15bddc0fe8d77f26a04181e89bfe841369c2f|6.49|2015-01-03 10:44:00|80.848351720559364|2|89604000100|11|35.082757871906274|0|25|1866|-80.806073|435|35.106477|PIMENTO|0.0|6|PALMETTO PIMENTO CHEESE|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00896040001004|SALADS|DELI|-80.848528|80.848554714125086|4|1
35.053394|a099da3d85a03a37e9b991b561d414e4c69a466a|3.99|2015-01-13 17:43:00|80.848351720559364|2|85290900329|11|35.082757872007456|0|25|1265|-80.78468|57|35.096737|ALMOND MILK|0.0|3|CALIFIA FRM ALM UNSWT VAN MILK|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00852909003695|MILK|DAIRY|-80.848528|80.848554547573357|30|1
35.053394|35d165b3b060ea598d687fa636ac2fed9fa19e2c|3.99|2015-02-11 19:30:00|80.848351720559364|2|85290900329|11|35.082757872007456|0|25|1265|-80.78468|57|35.096737|ALMOND MILK|0.0|3|CALIFIA FRM ALM UNSWT VAN MILK|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00852909003695|MILK|DAIRY|-80.848528|80.848554547573357|30|1
35.053394|6feb7ed244ca4195cdeef970aedd1acdec650ec5|8.29|2015-02-16 14:16:00|80.848351720559364|2|1258760034|11|35.082757871906274|0|25|443|-80.806073|76|35.106477|NFS-GARBAGE BAGS|0.0|1|GLAD FF D/S TALL KITCHEN|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00012587703557|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.848528|80.848554714125086|4|1
35.053394|ea9efb0a150593ac535e4a5b7796984b296cc20a|3.99|2015-02-07 16:06:00|80.848351720559364|2|1090000015|11|35.082757860980912|0|25|440|-80.825175|76|35.152722|NFS-ALUMINUM FOIL|0.0|1|REYNOLDS FOIL HEAVY DUTY 50 FT|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00010900000215|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.848528|80.848568883274552|160|1
35.053394|68816cfc768c57b4d3ceded29cf49fac55ef407a|9.98|2015-01-28 16:37:00|80.848351720559364|2|7203688187|11|35.082757872007456|0|25|561|-80.78468|64|35.096737|FR PROD ORGANIC PRODUCE|0.0|4|ORG HT BABY SPINACH 11 OZ|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00072036881878|FRESH PRODUCE|PRODUCE|-80.848528|80.848554547573357|30|2
35.053394|5a69e8bde66020825d448b2b64af97388e356291|4.99|2015-02-06 15:24:00|80.848351720559364|2|7203688187|11|35.082757872007456|0|25|561|-80.78468|64|35.096737|FR PROD ORGANIC PRODUCE|0.0|4|ORG HT BABY SPINACH 11 OZ|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00072036881878|FRESH PRODUCE|PRODUCE|-80.848528|80.848554547573357|30|1
35.053394|310b48bf4bfa1ea52a1fb338fa0a631667a5183f|3.55|2014-10-28 16:42:00|80.848351720559364|2|7332100027|11|35.082757872007456|0|25|251|-80.78468|43|35.096737|NON-DAIRY NOVELTIES|1.05|5|LUIGI'S MANGO ITALIAN ICE|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00073321044053|FROZEN NOVELTIES|FROZEN|-80.848528|80.848554547573357|30|1
35.053394|775d0a9a0c34ea7bb870f32fb7d31d3fa303d494|2.95|2015-02-18 19:16:00|80.848351720559364|2|7203663125|11|35.082757871906274|0|25|1262|-80.806073|57|35.106477|HALF N HALF WHIPPING CREAM|0.0|3|HT HEAVY WHIPPING CREAM|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00072036630988|MILK|DAIRY|-80.848528|80.848554714125086|4|1
35.053394|398394c0fd9a1c4a8dc047a01c4859c77c7dfa03|3.85|2014-09-18 18:34:00|80.848351720559364|2|7203663089|11|35.082757871906274|0|25|345|-80.806073|57|35.106477|ORGANIC MILK|0.0|3|HTO ORGANIC CRTN MILK 2%|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00072036630889|MILK|DAIRY|-80.848528|80.848554714125086|4|1
35.053394|11fbf77d905b615fecdb73b8bcd55336e22058b7|4.19|2015-03-06 13:34:00|80.848351720559364|2|7203663089|11|35.082757872007456|0|25|345|-80.78468|57|35.096737|ORGANIC MILK|0.0|3|HTO ORGANIC CRTN MILK 2%|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00072036630889|MILK|DAIRY|-80.848528|80.848554547573357|30|1
35.053394|8ec923b82ef0bf43f52e73a2305faff5d497760d|3.65|2014-11-07 11:31:00|80.848351720559364|2|4610000012|11|35.082757871906274|0|25|318|-80.806073|52|35.106477|SHREDDED/GRATED CHEESE|1.15|3|SARGENTO OTB MILD CHED FINE|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00046100000519|CHEESE|DAIRY|-80.848528|80.848554714125086|4|1
35.053394|66d571b5a1b8b1c38d8d1c74faaf9f29249b6cbf|9.99|2014-10-21 17:28:00|80.848351720559364|2|7203695679|11|35.082757872007456|0|25|1675|-80.78468|383|35.096737|PASTRY CASE PIES|0.0|14|"9"" TOPPED COCONUT CREAM PIE"|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00072036956798|PASTRY CASE|BAKERY|-80.848528|80.848554547573357|30|1
35.053394|ca4f3560212ad9204ceba90025da6073d7b5f252|0.79|2014-11-08 10:47:00|80.848351720559364|2|7203698208|11|35.082757874444468|0|25|257|-80.85753|39|35.116638|TOMATOES|0.0|1|HT TOMATO PASTE 6 BGO|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00072036982087|VEGETABLES-CAN/JAR|G1 GROCERY|-80.848528|80.848550161395963|204|1
35.053394|d3dc38b4a30fb64af3f7345f71a5ea9039a80237|1.0|2014-11-04 15:45:00|80.848351720559364|2||11|35.082757872007456|0|25|502|-80.78468|64|35.096737|FRESH BANANAS|0.0|4|BANANAS, YELLOW|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00204011000008|FRESH PRODUCE|PRODUCE|-80.848528|80.848554547573357|30|1
35.053394|f797659d92ff2828c62fe1f95f44dc50baac3ef9|1.1|2014-11-02 20:02:00|80.848351720559364|2||11|35.082757872007456|0|25|502|-80.78468|64|35.096737|FRESH BANANAS|0.0|4|BANANAS, YELLOW|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00204011000008|FRESH PRODUCE|PRODUCE|-80.848528|80.848554547573357|30|1
35.053394|0b3e074dfc9cd6b116c6992dc945001c75ed1001|5.37|2014-11-25 12:14:00|80.848351720559364|2|7348415501|11|35.082757852291103|0|25|13|-80.709466|2|35.124987|ROLLS/BISCUIT MIXES|0.5|1|HOUSE AUTRY SWT CORN BREAD MIX|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00073484155016|BAKING MIXES|G1 GROCERY|-80.848528|80.848577328019871|157|3
35.053394|0d90625c3bcd4128c297212280aca63b81e6c30a|1.79|2015-01-20 14:37:00|80.848351720559364|2|7348415501|11|35.082757871906274|0|25|13|-80.806073|2|35.106477|ROLLS/BISCUIT MIXES|0.0|1|HOUSE AUTRY SWT CORN BREAD MIX|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00073484155016|BAKING MIXES|G1 GROCERY|-80.848528|80.848554714125086|4|1
35.053394|daf4eec7c2529808e35661036a04d64ff30494cb|3.58|2015-01-01 11:51:00|80.848351720559364|2|7348415501|11|35.082757872007456|0|25|13|-80.78468|2|35.096737|ROLLS/BISCUIT MIXES|1.0|1|HOUSE AUTRY SWT CORN BREAD MIX|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00073484155016|BAKING MIXES|G1 GROCERY|-80.848528|80.848554547573357|30|2
35.053394|b584c7eea4677585c11dfdb91f7fe2d26adc2c75|0.47|2014-11-22 21:53:00|80.848351720559364|2|7248600220|11|35.082757871906274|0|25|11|-80.806073|2|35.106477|MUFFIN MIXES|0.0|1|JIFFY CORN MUFFIN MIX|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00072486002205|BAKING MIXES|G1 GROCERY|-80.848528|80.848554714125086|4|1
35.053394|5e0aebcec92643d3361b424c4756c14c038b0dec|3.97|2014-09-14 12:13:00|80.848351720559364|2|7203658035|11|35.082757874444468|0|25|358|-80.85753|100|35.116638|REGULAR BACON|0.97|19|HT REGULAR SLICED BACON|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00072036580351|BACON|CASE READY MEATS|-80.848528|80.848550161395963|204|1
35.053394|62eecef6df1e6415c6cfc357143eabf7e435ec4c|5.18|2014-11-15 21:12:00|80.848351720559364|2|2100061247|11|35.082757872007456|0|25|316|-80.78468|52|35.096737|CREAM CHEESE|1.18|3|PHILLY 1/3 FAT CREAM CHEESE|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00021000612475|CHEESE|DAIRY|-80.848528|80.848554547573357|30|2
35.053394|996b6cc79fb17020c031d6bca0498369f235e857|3.39|2014-09-21 18:56:00|80.848351720559364|2|1960005480|11|35.082757872007456|0|25|1269|-80.78468|41|35.096737|BREAKFAST SYRUP CARRIER|0.0|5|AUNT JEM BUTTERMILK PANCAKES|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00019600068204|BREAKFAST FOODS FROZEN|FROZEN|-80.848528|80.848554547573357|30|1
35.053394|af4ef4d5ab6a15e912b9f349967312a254b43cb7|0.69|2015-02-13 16:29:00|80.848351720559364|2||11|35.082757872007456|0|25|509|-80.78468|64|35.096737|FRESH CITRUS-REMAINING|0.0|4|LEMONS, LARGE|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00204053000004|FRESH PRODUCE|PRODUCE|-80.848528|80.848554547573357|30|1
35.053394|47676c961282022f9a132e7b6a3b1b8fab65b8ec|2.67|2014-09-11 14:52:00|80.848351720559364|2|7203670830|11|35.082757874444468|0|25|31|-80.85753|4|35.116638|NON CARBONATED WATER|0.0|1|(U)HT PURIFIED WATER .5L 32 PK|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00072036708304|BOTTLED WATER|G1 GROCERY|-80.848528|80.848550161395963|204|1
35.053394|6ce7a14bd6e6f6ecdd9b2d9094e5f2e9370fefe5|4.89|2014-09-12 21:32:00|80.848351720559364|2|4154861004|11|35.082757852291103|0|25|251|-80.709466|43|35.124987|NON-DAIRY NOVELTIES|0.0|5|EDY'S CREAMY COCONUT BARS|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00041548047638|FROZEN NOVELTIES|FROZEN|-80.848528|80.848577328019871|157|1
35.053394|7ac7f4d84f16115761e8daa4ca1e4b38a0f06972|3.99|2014-09-25 13:48:00|80.848351720559364|2|9418456076|11|35.082757879379905|0|25|583|-80.816172|136|35.059823|NUTS|0.0|4|TROPICAL DRIED CRANBERRIES|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00094184560764|OTHER MERCHANDISE|PRODUCE|-80.848528|80.848535645294604|66|1
35.053394|13c37ef2d38d0a27797534ad7e82d34247cc2aec|6.99|2014-11-20 13:05:00|80.848351720559364|2|3700013885|11|35.082757874444468|0|25|389|-80.85753|66|35.116638|NFS-LAUNDRY DETERGENTS|0.0|1|TIDE FREE & GENTLE 50OZ|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00037000138853|DETERGENTS|G1 GROCERY|-80.848528|80.848550161395963|204|1
35.053394|ffa2cd5b574bbd60a358c402c8655893819605a7|1.45|2014-10-28 16:45:00|80.848351720559364|2|7056097811|11|35.082757874444468|0|25|1272|-80.85753|50|35.116638|BAG VEG STEAM|0.0|5|PCTSWT STEAM BBY BRUSSELS|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00070560979511|VEGETABLES-FROZEN|FROZEN|-80.848528|80.848550161395963|204|1
35.053394|d36558911295158e29d70c1213294634fcdc8f8d|2.16|2014-12-23 17:57:00|80.848351720559364|2||11|35.082757871906274|0|25|561|-80.806073|64|35.106477|FR PROD ORGANIC PRODUCE|0.0|4|ORG BANANAS|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00294011000009|FRESH PRODUCE|PRODUCE|-80.848528|80.848554714125086|4|1
35.053394|5b36f5ce984e39948c3091762b9a3ddcc9eaef90|2.5|2015-01-15 17:45:00|80.848351720559364|2|7203698557|11|35.082757872007456|0|25|424|-80.78468|72|35.096737|NFS-FACIAL TISSUE|0.5|1|HT FACIAL TISSUE LOTION|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00072036985583|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.848528|80.848554547573357|30|2
35.053394|c6e6b1e2c6ec15cf4e070f6768018797e4e8d3dc|4.29|2015-02-18 16:03:00|80.848351720559364|2|7225000862|11|35.082757852291103|0|25|1038|-80.709466|164|35.124987|SWIRL/TOASTING|1.3|7|NATOWN CINNRAISIN BREAD|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00072250008624|BREAKFAST|COMMERCIAL BAKERY|-80.848528|80.848577328019871|157|1
35.053394|e4aff38668968497f471ed27b7fe99563568018c|6.98|2015-01-17 11:23:00|80.848351720559364|2|7203663995|11|35.082757874444468|0|25|342|-80.85753|57|35.116638|FRESH MILK|1.92|3|HARRIS TEETER 2% MILK|93ccf40dcbd22058bcfe4663b6f98bfa19c22aa1|2.0289731999909626|35.082633588753836|00072036639981|MILK|DAIRY|-80.848528|80.848550161395963|204|2
35.17335|c39f0b7c4f47f96b213f414cb59e40501b7a0c50|2.0|2014-10-02 09:35:00|1.4094857484078087|2|7203698753|174|0.6138907664563474|0|26|1272|-80.70901|50|35.17335|BAG VEG STEAM|0.0|5|HT RDY QUK YELLOW CORN|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00072036704191|VEGETABLES-FROZEN|FROZEN|-80.70901|1.4086379605250285|174|1
35.17335|5687cb547e5d01b77bf59b20816c692deb5cc90a|2.0|2014-10-16 10:18:00|1.4094857484078087|2|7203698753|174|0.6138907664563474|0|26|1272|-80.70901|50|35.17335|BAG VEG STEAM|0.0|5|HT RDY QUK YELLOW CORN|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00072036704191|VEGETABLES-FROZEN|FROZEN|-80.70901|1.4086379605250285|174|1
35.17335|31427ea63f3c6f144390f2dcde864fcae3db5eef|2.45|2014-10-30 10:07:00|1.4094857484078087|2|7040400100|174|0.6138907664563474|0|26|82|-80.70901|11|35.17335|VINEGAR|0.45|1|POMPEIAN VINEGAR RED WINE.|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00070404001002|CONDIMENTS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|18b43ddc1c603398fb40129e097d0941df5ddf4b|1.29|2015-02-12 10:24:00|1.4094857484078087|2|4920005675|174|0.6138907664563474|0|26|224|-80.70901|35|35.17335|SUGAR-BROWN|0.3|1|DOMINO DARK BROWN SUGAR-BX|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00049200056004|SUGAR/SUBSTITUTES|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|f92f778ecb36aef1fad7eef1e4d9c81cf1a5821f|1.29|2014-11-20 10:20:00|1.4094857484078087|2|4920005675|174|0.6138907664563474|0|26|224|-80.70901|35|35.17335|SUGAR-BROWN|0.3|1|DOMINO DARK BROWN SUGAR-BX|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00049200056004|SUGAR/SUBSTITUTES|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|68bc2c178a759b1c81916e6858429c94f0cfa809|3.99|2015-02-19 10:04:00|1.4094857484078087|2|5150000686|174|0.6138907664563474|0|26|123|-80.70901|19|35.17335|JELLY/JAMS|1.49|1|SMUCKER SEEDLES BLACKBERRY JAM|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00051500006849|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|3442471caab349bff3811afd7994c809ab50c56c|3.99|2014-10-23 13:22:00|1.4094857484078087|2|3425600064|174|0.6138907664563474|0|26|577|-80.70901|136|35.17335|OTHER MERCH FR MSC JUICE|0.49|4|HT APPLE CIDER, 64 OZ|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00072036880888|OTHER MERCHANDISE|PRODUCE|-80.70901|1.4086379605250285|174|1
35.17335|3ea7e5a7449ae614750c3257d6dc33e40cf2e383|7.98|2014-09-17 13:43:00|1.4094857484078087|2|3425600064|174|0.6138907664563474|0|26|577|-80.70901|136|35.17335|OTHER MERCH FR MSC JUICE|0.0|4|HT APPLE CIDER, 64 OZ|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00072036880888|OTHER MERCHANDISE|PRODUCE|-80.70901|1.4086379605250285|174|2
35.17335|c169791780ae991efb5a4acd1bc07c3ed1ba5a62|3.99|2015-01-15 10:17:00|1.4094857484078087|2|7203688078|174|0.6138907664563474|0|26|523|-80.70901|64|35.17335|FRESH POTATOES|0.0|4|HT RED POTATO 3LB BAG|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00072036880789|FRESH PRODUCE|PRODUCE|-80.70901|1.4086379605250285|174|1
35.17335|c20b09caab7a421013119c3b9dbcf363647f369b|1.77|2015-02-05 09:50:00|1.4094857484078087|2|7203657031|174|0.6138907664563474|0|26|322|-80.70901|53|35.17335|SOUR CREAM|0.0|3|HT SOUR CREAM|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00072036570314|CULTURES|DAIRY|-80.70901|1.4086379605250285|174|1
35.17335|c9da6a4412cbf1ccf227a398e72477a9be4aa408|2.79|2014-09-11 10:22:00|1.4094857484078087|2|1740011805|174|0.6138907664563474|0|26|239|-80.70901|38|35.17335|RICE-PACKAGED & BULK|0.0|1|MINUTE RICE INSTANT BROWN 14|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00017400118457|RICE GRAINS AND BEANS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|12240d79ad9281fa22fa9c8b751f8cd2eb7a0040|2.39|2014-12-18 10:14:00|1.4094857484078087|2|1340934115|174|0.6138907664563474|0|26|68|-80.70901|11|35.17335|BARBECUE SAUCES|0.51|1|SWEET BABY RAY BBQ SC SWT HOT|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00013409351000|CONDIMENTS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|9d1e62c9c58ac429edc721540e9042c04244aa6f|5.99|2014-11-28 15:50:00|1.4094857484078087|2|3760018888|174|0.6138907664563474|0|26|175|-80.70901|27|35.17335|CANNED MEATS|0.0|1|HORMEL CORNED BEEF|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00037600188883|PREPARED FOODS-RTS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|686b41e74eebbc85826befeb68bb60b20e1cd05e|1.67|2015-01-08 10:17:00|1.4094857484078087|2|7110000407|174|0.6138907664563474|0|26|183|-80.70901|28|35.17335|SALAD DRESSINGS-DRY|0.0|1|HVR DRS MIX RANCH ORIG 1OZ|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00071100004434|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|51dce5608221a12dd494f5a0490c536a28739970|1.27|2014-11-20 16:35:00|1.4094857484078087|2|7203628032|174|0.6138907664563474|0|26|163|-80.70901|25|35.17335|RELISHES|0.0|1|HT RELISH SWEET 16|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00072036280329|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|c839fa2425ae56b2bdf4800d928d515cb3c1b0ff|13.58|2015-01-22 09:35:00|1.4094857484078087|2|1200080994|174|0.6138907664563474|0|26|55|-80.70901|8|35.17335|REGULAR|3.39|23|CF PEPSI FRIDGEMATE|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00012000810022|CARBONATED BEVERAGES|BEVERAGE|-80.70901|1.4086379605250285|174|2
35.17335|c36353cb293a20dca7210c797105afa72414af30|2.99|2014-11-13 10:16:00|1.4094857484078087|2|1410009435|174|0.6138907664563474|0|26|28|-80.70901|26|35.17335|STUFFING PRODUCTS|0.3|1|PP2.99 PEP FARM HERB STUFFING|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00014100094357|PREPARED FOODS-DRY MIXES|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|52259fdd8ae120de694f2616af921ce1a0b6b3e6|3.35|2014-12-04 10:23:00|1.4094857484078087|2|1600042040|174|0.6138907664563474|0|26|13|-80.70901|2|35.17335|ROLLS/BISCUIT MIXES|0.0|1|BC BISQUICK|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00016000420403|BAKING MIXES|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|119d9fac1785968e562bd0b3574a44e2abef7b53|2.99|2014-11-06 10:50:00|1.4094857484078087|2|1410009435|174|0.6138907664563474|0|26|28|-80.70901|26|35.17335|STUFFING PRODUCTS|0.3|1|PP2.99 PEP FARM HERB STUFFING|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00014100094357|PREPARED FOODS-DRY MIXES|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|c2dc502b6f5031f48024d562650c77186c2f06d0|6.99|2014-10-24 09:25:00|1.4094857484078087|2|4100000873|174|0.6138907664563474|0|26|231|-80.70901|37|35.17335|INSTANT TEA|0.0|1|LIPTON DT ICE TEA MIX LMN FLVR|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00041000008733|TEA|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|b1d9ab0ab2a0c38406f091a4ff63e6b722dfe408|6.99|2015-01-29 10:04:00|1.4094857484078087|2|4100000873|174|0.6138907664563474|0|26|231|-80.70901|37|35.17335|INSTANT TEA|0.0|1|LIPTON DT ICE TEA MIX LMN FLVR|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00041000008733|TEA|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|2006fd18e05e6113e8729c345aada4d9b8315d52|6.99|2014-12-11 09:52:00|1.4094857484078087|2|4100000873|174|0.6138907664563474|0|26|231|-80.70901|37|35.17335|INSTANT TEA|0.0|1|LIPTON DT ICE TEA MIX LMN FLVR|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00041000008733|TEA|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|2c9bc21ff2070c54e0b4bdd53b5f6aa18371113d|6.99|2014-09-25 10:17:00|1.4094857484078087|2|4100000873|174|0.6138907664563474|0|26|231|-80.70901|37|35.17335|INSTANT TEA|0.0|1|LIPTON DT ICE TEA MIX LMN FLVR|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00041000008733|TEA|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|2a261685cd6300c3e0a20bcc016b4db49275e2ed|2.99|2014-12-31 10:03:00|1.4094857484078087|2|5209222318|174|0.6138907664563474|0|26|5826|-80.70901|1536|35.17335|FOILWARE BAKING|0.0|18|HANDI-FOIL 5LB LOAF PAN 2CT|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00052092223188|FOILWARE|GM|-80.70901|1.4086379605250285|174|1
35.17335|f6baa25734c79c877d98d2e2e57397be8586cdd6|5.49|2014-10-09 10:08:00|1.4094857484078087|2|7092200496|174|0.6138907664563474|0|26|5544|-80.70901|1508|35.17335|LDRY/IRON/VAC CLOSET STR|0.0|18|ENOZ MOTH BAR LAVENDER|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00070922004967|LAUNDRY/IRONING/VACUUM|GM|-80.70901|1.4086379605250285|174|1
35.17335|c5ae153737d583b02b1a5e03a5eae400cd08ab73|2.57|2015-03-05 09:57:00|1.4094857484078087|2|7203655996|174|0.6138907664563474|0|26|316|-80.70901|52|35.17335|CREAM CHEESE|0.0|3|HT LIGHT SOFT CREAM CHEESE|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00072036559975|CHEESE|DAIRY|-80.70901|1.4086379605250285|174|1
35.17335|d33ad12116752df134840aaf49ef936ad5a8c7ae|3.99|2015-02-25 11:34:00|1.4094857484078087|2|4300000037|174|0.6138907664563474|0|26|228|-80.70901|36|35.17335|TABLE SYRUP|2.0|1|LOG CABIN SYRUP|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00043000000373|TABLE SYRUPS|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|c994b1f56e67d253690aada092163bc1a7b51444|2.59|2014-11-08 10:49:00|1.4094857484078087|2|7203663996|174|0.6138907664563474|0|26|342|-80.70901|57|35.17335|FRESH MILK|0.0|3|HARRIS TEETER 2%   MILK|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00072036639998|MILK|DAIRY|-80.70901|1.4086379605250285|174|1
35.17335|659548f3722eec750ff50a3af41b56800f3f617a|2.19|2014-09-19 17:03:00|1.4094857484078087|2|76857300210|174|0.6138907664563474|0|26|544|-80.70901|64|35.17335|FRESH PRODUCE FRSH HERBS|0.2|4|PKG FRESH THYME|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00768573001601|FRESH PRODUCE|PRODUCE|-80.70901|1.4086379605250285|174|1
35.17335|45a3e3b3a995227154c389cc53a007fced7efec0|1.67|2015-02-07 17:03:00|1.4094857484078087|2|7203614064|174|0.6138907664563474|0|26|110|-80.70901|16|35.17335|FRUIT-CORE|0.33|1|HT PEAR LITE SLICES JC 15|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00072036140647|FRUIT-CAN/JAR|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|6ce3820203d7da71b69367db4a6fc20d244a7c8b|19.84|2014-12-22 10:44:00|1.4094857484078087|2|23520300000|174|0.6138907664563474|0|26|646|-80.70901|202|35.17335|COUNTRY HAMS|0.0|2|OLD WAYNESBORO CENTER SLICES|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00235203000001|SMOKED HAMS|MEAT|-80.70901|1.4086379605250285|174|3
35.17335|cb6c87b55f218d89afaf08c2c364cc2787bf4eb5|11.97|2014-10-28 09:44:00|80.709059419360486|2|7203698238|174|35.211915308165963|0|31|402|-80.810056|76|35.219587|NFS-DISPOSABLE CONTAINER|1.47|1|YH SOUP/SALAD CONTAINER|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|35.187384292804154|00072036982384|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.70901|80.709011080270145|401|3
35.17335|4763cac8a64b5ec5c9eb989d5be90cc2d2b72062|2.19|2014-09-18 15:20:00|1.4094857484078087|2|64420931131|174|0.6138907664563474|0|26|8|-80.70901|2|35.17335|BROWNIE MIXES|0.0|1|D HINES DARK CHOC FUDGE BRWNIE|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00644209420957|BAKING MIXES|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|5f3f27808e3425cb2769b9b4d1fdac919b70efdd|7.3|2015-03-09 14:10:00|1.4094857484078087|2|3010003012|174|0.6138907664563474|0|26|91|-80.70901|13|35.17335|SPRAYED BUTTER CRACKERS|2.3|1|KEELBER CLUB ORIGINAL|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00030100100577|CRACKERS|G1 GROCERY|-80.70901|1.4086379605250285|174|2
35.17335|64226ec4a0bf8e9848bff40355e6197cba0d977b|2.45|2014-11-18 12:19:00|1.4094857484078087|2|5100013279|174|0.6138907664563474|0|26|214|-80.70901|33|35.17335|BROTH|0.45|1|SWANSON BROTH LOW SOD CHICKEN|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00051000132796|SOUP|G1 GROCERY|-80.70901|1.4086379605250285|174|1
35.17335|a0b4b2b4d950d68d0af30fa10972139516080013|8.98|2014-12-07 15:39:00|1.4094857484078087|2|7203695755|174|0.6138907664563474|0|26|1647|-80.70901|379|35.17335|PACKAGED MUFFINS|0.0|14|12CT MINI ASSORTED MUFFINS|943ba52037ce2811260d80d0feddae09a98bca6a|2.6647696630818323|0.61471665291522548|00072036957573|MUFFINS|BAKERY|-80.70901|1.4086379605250285|174|2
35.603432|2406c138b82c7d833d0e654b870767bf869b553d|3.99|2014-12-18 22:19:00|1.4102725052409182|2|84921900730|274|0.6213971134099097|0|1|7350|-80.895009|1600|35.603432|CHRISTMAS GIFT BOX IMP|1.5|18|HDAY G/CARD HLDR 3 PK|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00849219007307|SEASONAL MERCHANDISE|GM|-80.895009|1.4118842554804456|274|1
35.603432|a01e32a57f19a45af00b87f25ca261b90086ed28|5.99|2014-11-17 16:41:00|1.4102725052409182|2|7430500132|274|0.6213971134099097|0|1|82|-80.895009|11|35.603432|VINEGAR|0.0|1|BRAGG ORG VINEGAR APPLE CIDER|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00074305001321|CONDIMENTS|G1 GROCERY|-80.895009|1.4118842554804456|274|1
35.603432|93912ece7b8dad6d6c7899411005bbd8f34ad022|6.49|2014-12-04 21:12:00|1.4102725052409182|2|7800001180|274|0.6213971134099097|0|1|55|-80.895009|8|35.603432|REGULAR|0.0|23|CRUSH ORANGE 12PK|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00078000013054|CARBONATED BEVERAGES|BEVERAGE|-80.895009|1.4118842554804456|274|1
35.603432|9625b9a72b18cf4920cb4941092b42972de6ae43|3.77|2015-02-14 09:00:00|1.4102725052409182|2|7203603040|274|0.6213971134099097|0|1|217|-80.895009|34|35.603432|EXTRACTS FOOD COLORING|0.0|1|HT VANILLA EXTRACT|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00072036030405|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.895009|1.4118842554804456|274|1
35.603432|77c3b1fb20cf0f0b2d7c93bbf40f79553ed487ca|1.79|2014-09-18 17:33:00|1.4102725052409182|2|8079380770|274|0.6213971134099097|0|1|99|-80.895009|32|35.603432|LIQUID TEA|0.68|1|D FUZE SLENDER TROPICAL PUNCH|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00080793807765|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.895009|1.4118842554804456|274|1
35.603432|08b539dfb888d63fa00cc90c576db37f8cbcc566|5.99|2014-12-22 17:44:00|1.4102725052409182|2|7756725423|274|0.6213971134099097|0|1|252|-80.895009|45|35.603432|PREMIUM ICE CREAM|3.0|5|BREYERS STRAWBERRY ICE CREAM|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00077567254344|ICE CREAM|FROZEN|-80.895009|1.4118842554804456|274|1
35.603432|4bee73f98a643d6dae84b1b9e50f842dd145ad82|1.88|2015-01-01 15:42:00|1.4102725052409182|2|7248600220|274|0.6213971134099097|0|1|11|-80.895009|2|35.603432|MUFFIN MIXES|0.12|1|JIFFY CORN MUFFIN MIX|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00072486002205|BAKING MIXES|G1 GROCERY|-80.895009|1.4118842554804456|274|4
35.603432|ac178e0b6e6f7d6577d60b77e6a5656e33036f8d|1.99|2014-10-18 17:53:00|1.4102725052409182|2|7294075600|274|0.6213971134099097|0|1|257|-80.895009|39|35.603432|TOMATOES|0.49|1|TUTTOROSSO TOMATO CRUSH BASIL|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00072940756002|VEGETABLES-CAN/JAR|G1 GROCERY|-80.895009|1.4118842554804456|274|1
35.603432|f847e9fbf2deb7d8e256bac9d4c0ff9baa4c1ab7|8.38|2015-02-04 15:49:00|1.4102725052409182|2|76026300010|274|0.6213971134099097|0|1|213|-80.895009|33|35.603432|SOUP MIXES|0.5|1|BEARCREEK SOUP MIX CRMY POTATO|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00760263000161|SOUP|G1 GROCERY|-80.895009|1.4118842554804456|274|2
35.603432|99be7bd376cdf40cf2c7adfe2baced7d2d79465e|1.99|2014-09-27 09:39:00|1.4102725052409182|2|7203648011|274|0.6213971134099097|0|1|274|-80.895009|44|35.603432|ICE|0.0|5|HT BAGGED ICE 10LB (456)|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00000000004560|ICE|FROZEN|-80.895009|1.4118842554804456|274|1
35.603432|89a2b1340ceefefca911f659f5bfec9efc38146d|2.39|2014-10-30 14:56:00|1.4102725052409182|2|1410008550|274|0.6213971134099097|0|1|89|-80.895009|12|35.603432|GRAHAM CRACKERS|0.2|1|PP GF SWEET GRAHAM VANILLA CUP|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00014100096061|COOKIES|G1 GROCERY|-80.895009|1.4118842554804456|274|1
35.603432|dabf4bf23667729abc9030a0214f00706afbb934|6.67|2015-01-01 19:41:00|1.4102725052409182|2|7203642992|274|0.6213971134099097|0|1|236|-80.895009|38|35.603432|DRY BEANS|0.34|1|HT PEAS DRY GREEN SPLIT|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00072036420671|RICE GRAINS AND BEANS|G1 GROCERY|-80.895009|1.4118842554804456|274|5
35.603432|8e2bcf8924eb46af2ab88495f9f70c47f67b28e3|2.99|2014-12-12 07:02:00|1.4102725052409182|2|3080000189|274|0.6213971134099097|0|1|52|-80.895009|7|35.603432|PKG NON CHOC|0.0|1|DUM DUM POPS SPANGLER LAY DOWN|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00030800001891|CANDY|G1 GROCERY|-80.895009|1.4118842554804456|274|1
35.603432|d55c8db7a1def77a224853da826c082b1b9de44f|5.98|2015-01-09 07:03:00|1.4102725052409182|2|3080000189|274|0.6213971134099097|0|1|52|-80.895009|7|35.603432|PKG NON CHOC|0.0|1|DUM DUM POPS SPANGLER LAY DOWN|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00030800001891|CANDY|G1 GROCERY|-80.895009|1.4118842554804456|274|2
35.603432|496733c13e83a6316fa95ac254a57435a56abdfc|2.99|2014-10-02 06:54:00|1.4102725052409182|2|3080000189|274|0.6213971134099097|0|1|52|-80.895009|7|35.603432|PKG NON CHOC|0.0|1|DUM DUM POPS SPANGLER LAY DOWN|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00030800001891|CANDY|G1 GROCERY|-80.895009|1.4118842554804456|274|1
35.603432|aeac16206bc17ffc8777c7b8a04b3271492644a3|5.98|2015-01-22 14:41:00|1.4102725052409182|2|3080000189|274|0.6213971134099097|0|1|52|-80.895009|7|35.603432|PKG NON CHOC|0.98|1|DUM DUM POPS SPANGLER LAY DOWN|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00030800001891|CANDY|G1 GROCERY|-80.895009|1.4118842554804456|274|2
35.603432|833ddfb582738236c19dcc33353f09229737c1ac|3.11|2014-12-10 21:21:00|1.4102725052409182|2||274|0.6213971134099097|0|1|524|-80.895009|64|35.603432|FRESH PROD FRESH ONIONS|0.0|4|COO PEELED RED ONIONS|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00204667000001|FRESH PRODUCE|PRODUCE|-80.895009|1.4118842554804456|274|1
35.603432|9cf6bb6be58178e16285f5943e6299ab1695af92|1.77|2014-10-29 18:08:00|1.4102725052409182|2|7203657031|274|0.6213971134099097|0|1|322|-80.895009|53|35.603432|SOUR CREAM|0.0|3|HT LIGHT SOUR CREAM|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00072036590343|CULTURES|DAIRY|-80.895009|1.4118842554804456|274|1
35.603432|77aadfe6b0591b986cb29b781e7fd4d3fd0aaed0|3.75|2014-11-13 17:33:00|1.4102725052409182|2|1600048796|274|0.6213971134099097|0|1|74|-80.895009|9|35.603432|RTE CEREAL ALL FAMILY|0.0|1|GM RICE CHEX|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00016000487949|CEREAL|G1 GROCERY|-80.895009|1.4118842554804456|274|1
35.603432|69c159b21241f5a3ede1329b66684c4e6029294b|8.97|2014-09-27 07:39:00|1.4102725052409182|2|1600018910|274|0.6213971134099097|0|1|1200|-80.895009|6|35.603432|FRUIT SNACKS|0.99|1|FRUIT ROLL-UPS FLAVOR MIXERS|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00016000454729|BREAKFAST FOODS|G1 GROCERY|-80.895009|1.4118842554804456|274|3
35.603432|928bc80903a18e2c71b2f673689f9a2e6d259736|3.0|2014-12-24 07:01:00|1.4102725052409182|2|7203632016|274|0.6213971134099097|0|1|195|-80.895009|30|35.603432|SALAD & COOKING OIL|0.5|1|HT CANOLA OIL|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00072036320162|SHORTENING/OIL|G1 GROCERY|-80.895009|1.4118842554804456|274|1
35.603432|3947b46e2e8ac5212d0e7f5e4f13dd90fd08f46e|5.78|2014-12-22 06:52:00|1.4102725052409182|2|7203663102|274|0.6213971134099097|0|1|339|-80.895009|57|35.603432|EGGNOGS/DRINKS|0.89|3|I/O HARRIS TEETER EGG NOG|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00072036631022|MILK|DAIRY|-80.895009|1.4118842554804456|274|2
35.603432|fcff95893c607b58235ea7d1e9a35b17086e322d|2.39|2015-02-01 14:38:00|1.4102725052409182|2|7357013000|274|0.6213971134099097|0|1|1267|-80.895009|53|35.603432|DIPS AND SPREADS|0.89|3|HELUVA GOOD FRENCH ONION DIP|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00073570130002|CULTURES|DAIRY|-80.895009|1.4118842554804456|274|1
35.603432|0cda9e8bb25161f8c25124852f7a250e710faf7f|4.78|2015-02-16 14:14:00|1.4102725052409182|2|7357013000|274|0.6213971134099097|0|1|1267|-80.895009|53|35.603432|DIPS AND SPREADS|1.2|3|HELUVA GOOD FRENCH ONION DIP|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00073570130002|CULTURES|DAIRY|-80.895009|1.4118842554804456|274|2
35.603432|8a472f4cb7b043d90cefc826c355df9c207f5bbc|5.85|2014-12-21 19:59:00|1.4102725052409182|2|64420941000|274|0.6213971134099097|0|1|10|-80.895009|2|35.603432|LAYER CAKE MIX|2.0999999999999996|1|D HINES YELLOW CAKE MIX|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00644209410200|BAKING MIXES|G1 GROCERY|-80.895009|1.4118842554804456|274|3
35.603432|901d0c0bde7ec347271c83fc62c9d2625ed87bbf|15.599999999999998|2014-12-16 18:32:00|1.4102725052409182|2|64420941000|274|0.6213971134099097|0|1|10|-80.895009|2|35.603432|LAYER CAKE MIX|0.7|1|D HINES YELLOW CAKE MIX|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00644209410200|BAKING MIXES|G1 GROCERY|-80.895009|1.4118842554804456|274|8
35.603432|53833be59e22d0f6ff740816c79c8712735d4a0c|4.29|2014-09-13 18:39:00|1.4102725052409182|2|70897111899|274|0.6213971134099097|0|1|1703|-80.895009|387|35.603432|SEASONAL COOKIES|0.8|14|HARVEST ORANGE FRSTD SGR COOK|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00708971118990|COOKIES|BAKERY|-80.895009|1.4118842554804456|274|1
35.603432|97d0b77d1eab9de9bd4b92ef581db8a6e4dc69a1|4.69|2014-12-23 20:26:00|80.891462859624312|2|5210007064|274|35.624236450782313|0|45|217|-80.875654|34|35.585842|EXTRACTS FOOD COLORING|1.41|1|MC BUTTER FLAVORING|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|35.636605227883024|00052100070711|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.895009|80.895011405058398|99|1
35.603432|a13bf981764dbdaa2b40ee35d03533250c0e352f|10.649999999999999|2015-02-25 16:43:00|1.4102725052409182|2|3800039125|274|0.6213971134099097|0|1|74|-80.895009|9|35.603432|RTE CEREAL ALL FAMILY|1.05|1|KELLOGG RICE KRISPIES 9|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00038000318443|CEREAL|G1 GROCERY|-80.895009|1.4118842554804456|274|3
35.603432|6a2df3b0b5a237f1843e31a43cdff24c9c34251b|8.99|2015-01-31 18:33:00|1.4102725052409182|2|7203695532|274|0.6213971134099097|0|1|1659|-80.895009|381|35.603432|VARIETY SINGLE LAYER|2.0|14|SGL LAYER RED VELVET CAKE|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00072036955326|CAKES|BAKERY|-80.895009|1.4118842554804456|274|1
35.603432|6ba3a70d96df570bd2f9da4227512f83d10a83b7|2.99|2015-02-13 19:32:00|1.4102725052409182|2|1800000338|274|0.6213971134099097|0|1|327|-80.895009|54|35.603432|DINNER ROLLS-REFRIGERATED|0.0|3|PILLS CRUSTY FRENCH LOAF BREAD|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00018000004683|DOUGH PRODUCTS|DAIRY|-80.895009|1.4118842554804456|274|1
35.603432|79b37b074ee538cc772a61351eeab7ee2ae62225|3.39|2014-09-18 21:33:00|1.4102725052409182|2|5100012573|274|0.6213971134099097|0|1|137|-80.895009|20|35.603432|TOMATO & VEGETABLE JUICE|0.89|1|V8 SPLASH BERRY BLEND|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00051000127112|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.895009|1.4118842554804456|274|1
35.603432|7c4e95be0c39b4644c067f4e20309449b7d5691d|3.99|2014-10-05 11:38:00|1.4102725052409182|2|4000015140|274|0.6213971134099097|0|1|46|-80.895009|7|35.603432|PKG CHOC|0.49|1|TWIX FUNSIZE|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00040000151784|CANDY|G1 GROCERY|-80.895009|1.4118842554804456|274|1
35.603432|960e6412ff61177624a7b3635df967201f5db322|2.97|2014-10-08 06:58:00|80.891462859624312|2|7203675058|274|35.624236450782313|0|45|3917|-80.875654|1075|35.585842|DISPOSABLE RAZOE-MEN|0.0|17|HT TRIPLE BLADE DISPOSABLE MEN|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|35.636605227883024|00072036750587|SHAVING NEEDS/MEN HAIR|HBC|-80.895009|80.895011405058398|99|1
35.603432|7988f8447ce1f25d443f331e534dc1820c825061|5.77|2014-09-24 16:18:00|1.4102725052409182|2|7203698516|274|0.6213971134099097|0|1|426|-80.895009|72|35.603432|NFS-PAPER TOWELS|0.8|1|YH TOWEL 8RL WHITE|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00072036985156|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.895009|1.4118842554804456|274|1
35.603432|d52ceea8ccc1774c76d3a705d1bc79745e6c23cc|9.98|2015-01-14 16:41:00|1.4102725052409182|2|6827493471|274|0.6213971134099097|0|1|31|-80.895009|4|35.603432|NON CARBONATED WATER|2.0|1|NESTLE PURE LIFE .5L 24PK|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00068274934711|BOTTLED WATER|G1 GROCERY|-80.895009|1.4118842554804456|274|2
35.603432|4f7078f6da4e0a14bd8a9f2aaa47804739d758fd|3.98|2014-12-13 07:17:00|1.4102725052409182|2|4900004574|274|0.6213971134099097|0|1|171|-80.895009|20|35.603432|ISOTONIC DRINKS|2.6|1|POWERADE LEMON LIME|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00049000045734|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.895009|1.4118842554804456|274|2
35.603432|2d44da157f4e99531886e866e75d8a354f436699|4.49|2014-12-29 09:09:00|1.4102725052409182|2|4000031532|274|0.6213971134099097|0|1|727|-80.895009|7|35.603432|SEASONAL CANDY-SINGLE FAC|2.25|1|I/O(C14)M&M PLAIN CHRISTMAS|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00040000315322|CANDY|G1 GROCERY|-80.895009|1.4118842554804456|274|1
35.603432|5d5a58bcc9103d4460128e29227e342b87ca383c|4.99|2015-02-09 19:34:00|1.4102725052409182|2|4900002468|274|0.6213971134099097|0|1|54|-80.895009|8|35.603432|DIET|0.0|23|DIET COKE .5 LITER/6 PK.|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00049000024692|CARBONATED BEVERAGES|BEVERAGE|-80.895009|1.4118842554804456|274|1
35.603432|ad078d980ae394246dd9b2ed897123ea8c86e062|3.99|2014-11-03 15:07:00|1.4102725052409182|2|3400038826|274|0.6213971134099097|0|1|727|-80.895009|7|35.603432|SEASONAL CANDY-SINGLE FAC|2.0|1|I/O(H15)FH ROLO MINIATURES BAG|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00034000388264|CANDY|G1 GROCERY|-80.895009|1.4118842554804456|274|1
35.603432|0776b6f858cfca5e5cfb4c6c8c7e3f2ead20282f|6.39|2014-10-05 17:14:00|1.4102725052409182|2|3040077377|274|0.6213971134099097|0|1|427|-80.895009|72|35.603432|NFS-TOILET TISSUE|0.0|1|ANGEL SOFT SOFT/STRONG 12DR|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00030400773778|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.895009|1.4118842554804456|274|1
35.603432|c790ae37ce7a3c6989ab1d976152e11a1b83b050|7.58|2014-12-31 15:42:00|1.4102725052409182|2|2500005542|274|0.6213971134099097|0|1|335|-80.895009|56|35.603432|ORANGE JUICE-REGRIGERATED|1.58|3|SIMPLY ORANGE GROVE MADE|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00025000055447|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.895009|1.4118842554804456|274|2
35.603432|359fd2a7cd8626fb61f914e0512431c040cdb23a|1.79|2015-01-02 08:05:00|1.4102725052409182|2|1200000157|274|0.6213971134099097|0|1|31|-80.895009|4|35.603432|NON CARBONATED WATER|0.79|1|AQUAFINA WATER  1 LITER|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00012000001574|BOTTLED WATER|G1 GROCERY|-80.895009|1.4118842554804456|274|1
35.603432|c3535a30a5e5429084260e5e8ddc73888f92e42a|7.78|2015-01-04 14:26:00|1.4102725052409182|2|4900002468|274|0.6213971134099097|0|1|54|-80.895009|8|35.603432|DIET|0.0|23|DT SUNDROP .5 LITER 6PK|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00078000231427|CARBONATED BEVERAGES|BEVERAGE|-80.895009|1.4118842554804456|274|2
35.603432|81944c618a7f0add53191c683c8f76cd9988b9b3|2.99|2015-02-25 20:27:00|1.4102725052409182|2|9418456066|274|0.6213971134099097|0|1|583|-80.895009|136|35.603432|NUTS|0.0|4|TROPICAL SUNFLOWER SEEDS R/S|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00094184560665|OTHER MERCHANDISE|PRODUCE|-80.895009|1.4118842554804456|274|1
35.603432|6417f7ed3f9a20372790028be3a97e1443029f40|3.55|2014-11-29 16:07:00|1.4102725052409182|2|7433610102|274|0.6213971134099097|0|1|342|-80.895009|57|35.603432|FRESH MILK|1.08|3|HIGHLAND CREST SKIM MILK|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00074336101083|MILK|DAIRY|-80.895009|1.4118842554804456|274|1
35.603432|b8d5f40c613c2cd5c3be4db995c3c5305923d7c4|4.49|2014-10-13 18:45:00|1.4102725052409182|2|71575620002|274|0.6213971134099097|0|1|504|-80.895009|64|35.603432|FRESH BERRIES|0.5|4|STRAWBERRIES 1LB CLAM|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00812049005102|FRESH PRODUCE|PRODUCE|-80.895009|1.4118842554804456|274|1
35.603432|afa19876fdfe1c56e1a1bfe306582e927ee13651|3.49|2015-01-19 18:36:00|1.4102725052409182|2|7092500046|274|0.6213971134099097|0|1|54|-80.895009|8|35.603432|DIET|0.0|23|DIET CHEERWINE .5 LTR 6 PK|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00070925000461|CARBONATED BEVERAGES|BEVERAGE|-80.895009|1.4118842554804456|274|1
35.603432|6028d2fe0aafb5673aaab29cad09b9553d7b57f5|6.99|2015-01-01 18:35:00|1.4102725052409182|2|7203670333|274|0.6213971134099097|0|1|443|-80.895009|76|35.603432|NFS-GARBAGE BAGS|1.02|1|YH TALL KITCHN BAGS VANILLA 13|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00072036707024|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.895009|1.4118842554804456|274|1
35.603432|27c1b448514ff363d9da7012a4bedc372a411a8e|1.59|2014-11-23 08:53:00|1.4102725052409182|2|7203698008|274|0.6213971134099097|0|1|442|-80.895009|76|35.603432|NFS-COOKING-STORAGE BAGS|0.0|1|YOUR HOME LUNCH BAGS 50 CT|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00072036980083|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.895009|1.4118842554804456|274|1
35.603432|551e626e577ae4ff12cb7250004b9d6250239ca0|3.88|2014-12-17 06:13:00|80.891462859624312|2|4300020431|274|35.624236450782313|0|45|94|-80.875654|14|35.585842|PUDDING MIXES|0.22|1|JELLO INST PUDDING VANILLA|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|35.636605227883024|00043000204337|DESSERTS/GELS/SYRUPS|G1 GROCERY|-80.895009|80.895011405058398|99|4
35.603432|b8f5c42a75eac82161280d21ab1aca76bd4aa48e|8.97|2015-01-22 17:39:00|1.4102725052409182|2|7203659051|274|0.6213971134099097|0|1|318|-80.895009|52|35.603432|SHREDDED/GRATED CHEESE|0.0|3|(U)HT FANCY SHRED MEXICAN CHS|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00072036590503|CHEESE|DAIRY|-80.895009|1.4118842554804456|274|1
35.603432|fb44d476b6d9c13b4484f498e1be93fd4865f9cd|0.99|2014-09-18 14:48:00|1.4102725052409182|2|3400000031|274|0.6213971134099097|0|1|47|-80.895009|7|35.603432|REGISTER BARS|0.5|1|HERSHEY MILK CHOC BAR|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00034000002405|CANDY|G1 GROCERY|-80.895009|1.4118842554804456|274|1
35.603432|49a204f0592a20be898342138c9d1c46af07f4d4|5.0|2015-02-14 20:06:00|1.4102725052409182|2||274|0.6213971134099097|0|1|1645|-80.895009|379|35.603432|BULK (MUFFINS)|0.0|14|BULK MUFFINS|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00072036959591|MUFFINS|BAKERY|-80.895009|1.4118842554804456|274|4
35.603432|f3fbc27696fc58ac0148d97c966074fb6d9e0e9d|6.5|2014-12-30 10:06:00|1.4102725052409182|2|3700007100|274|0.6213971134099097|0|1|393|-80.895009|68|35.603432|NFS-AIR FRESHENERS|0.25|1|I/O FEBREZE AE VANILLA LATTE|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00037000866961|FRESHENERS/DEODORIZERS|G1 GROCERY|-80.895009|1.4118842554804456|274|2
35.603432|89a597ff186e2972b94e65cc24c082989e832d60|6.98|2014-12-31 15:43:00|1.4102725052409182|2|7203663995|274|0.6213971134099097|0|1|342|-80.895009|57|35.603432|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00072036631282|MILK|DAIRY|-80.895009|1.4118842554804456|274|2
35.603432|50984b138f8d3593ed48245cb7b0eb90382fea88|13.98|2015-02-16 17:22:00|1.4102725052409182|2|71921820201|274|0.6213971134099097|0|1|6204|-80.895009|1548|35.603432|HIGH END|0.0|18|PURAFILTER GOLD 20/20/1|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00719218202013|FURNACE FILTERS|GM|-80.895009|1.4118842554804456|274|2
35.603432|f763dcb8028ecbada1cefaaa284db3563761f604|6.99|2015-01-12 14:47:00|1.4102725052409182|2|4900002890|274|0.6213971134099097|0|1|54|-80.895009|8|35.603432|DIET|2.0|23|FRESCA 12OZ 12PK FRIDGEPACK CN|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00049000031058|CARBONATED BEVERAGES|BEVERAGE|-80.895009|1.4118842554804456|274|1
35.603432|d153384de3ff072ea6a48132395f46066233d682|3.38|2014-09-19 18:30:00|1.4102725052409182|2|4900000044|274|0.6213971134099097|0|1|54|-80.895009|8|35.603432|DIET|0.0|23|CB DIET COKE CONTOUR 20 OZ NR|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00049000000450|CARBONATED BEVERAGES|BEVERAGE|-80.895009|1.4118842554804456|274|2
35.603432|46121f090b0cc22787ac8151f46913d6f57421c4|5.45|2014-09-25 16:08:00|1.4102725052409182|2|7203697668|274|0.6213971134099097|0|1|317|-80.895009|52|35.603432|CHUNK AND BAR CHEESE|1.95|3|HT NY SHARP CHEDDAR CHEESE|9926159a4d1f7d29adb4c13db62798e9b22d38e8|1.4375373144565273|0.61833652052202714|00072036979551|CHEESE|DAIRY|-80.895009|1.4118842554804456|274|1
35.444615|b0d0fde42bece58fb0786d4c5177c30ae0e20369|0.67|2014-11-15 11:05:00|1.4102725052409182|2|7203641111|340|0.6186252338517699|0|1|242|-80.861571|39|35.444615|CANNED BEANS|0.0|1|HT BEANS PINTO|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00072036411112|VEGETABLES-CAN/JAR|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.444615|dd84464d2fecb3da13b49020f2fff12b98bf504d|2.89|2014-12-07 12:33:00|1.4102725052409182|2|7203655029|340|0.6186252338517699|0|1|331|-80.861571|52|35.444615|NATURAL SLICED|0.39|3|HT PROVOLONE SLICES|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00072036550170|CHEESE|DAIRY|-80.861571|1.4113006522851637|340|1
35.444615|e66cd34eb2b4f317ad8b4207bf1bbb49246facc1|2.35|2014-10-05 13:16:00|1.4102725052409182|2|4112907700|340|0.6186252338517699|0|1|1219|-80.861571|275|35.444615|PASTA SC CORE|0.0|1|CLASSICO SC SPICY TOMATO PESTO|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00041129077757|PASTA SAUCES|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.444615|33b0e0a3a027517af755c7b53000fc1255677366|3.49|2014-10-19 13:26:00|1.4102725052409182|2|7203676172|340|0.6186252338517699|0|1|92|-80.861571|13|35.444615|REMAINING CRACKERS|1.49|1|HTT WHEAT SNACK CRACKER|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00072036761712|CRACKERS|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.444615|7e0ca0be5d264ce5b0e9f2a98bd824701129d89e|3.99|2014-10-14 17:07:00|1.4102725052409182|2|7203688076|340|0.6186252338517699|0|1|523|-80.861571|64|35.444615|FRESH POTATOES|0.5|4|HT RUSSET POTATO 5LB BAG|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00072036880765|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|746b19b2fba990811427187fbe679f6ae023e2f6|1.69|2014-10-18 18:40:00|1.4102725052409182|2|7203688003|340|0.6186252338517699|0|1|527|-80.861571|64|35.444615|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00072036880031|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|afdec51a58dc46c730e6a5e2c13cfa9bf1564346|1.69|2014-11-22 13:23:00|1.4102725052409182|2|7203688003|340|0.6186252338517699|0|1|527|-80.861571|64|35.444615|FRESH CARROTS|0.0|4|HT BABY CARROTS 1LB BAG|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00072036880031|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|b8d33f9f63c0a39aabf09f3fefc653bb7e4ba512|1.69|2014-11-01 12:03:00|1.4102725052409182|2|7203688003|340|0.6186252338517699|0|1|527|-80.861571|64|35.444615|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00072036880031|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|bc80859982ff94048c8f177fac5dcbfb59416200|3.38|2014-12-13 15:32:00|1.4102725052409182|2|7203688003|340|0.6186252338517699|0|1|527|-80.861571|64|35.444615|FRESH CARROTS|0.0|4|HT BABY CARROTS 1LB BAG|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00072036880031|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|2
35.444615|28022c816ff7cfb00a60d2e4e051bf0dbef54b16|4.0|2014-11-15 17:34:00|1.4102725052409182|2|84115200793|340|0.6186252338517699|0|1|1165|-80.861571|87|35.444615|NFS-FRESH CONSUMER BUNCH|0.0|9|BUNCH -3/$12 NOVELTY DISBUDS|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00841152007932|FLORAL|FLORAL|-80.861571|1.4113006522851637|340|1
35.444615|65fc9aa57f887ad67dade1ec4dd2700a5b5aa047|2.4|2015-03-03 17:49:00|80.86161257435397|2|81829001314|340|35.455082584258413|0|36|685|-80.860108|61|35.500972|GREEK|0.0|3|CHOBANI 100 PEACH|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|35.472272108304431|00818290013156|YOGURT|DAIRY|-80.861571|80.861578596363103|268|2
35.444615|eadfd6da1f25ca618fdbc1deacb8f2600ff46711|11.99|2015-03-05 19:23:00|1.4102725052409182|2|8254400801|340|0.6186252338517699|0|1|9948|-80.861571|886|35.444615|NFS-PREM-CAB SAUVIGNON|0.0|13|3 GIRLS CABERNET|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00082544008018|PREMIUM ($8-$10.99)|WINE|-80.861571|1.4113006522851637|340|1
35.444615|4da0e3b69c7c96895206788e3a585d3c6ab14376|0.87|2014-11-26 18:08:00|1.4102725052409182|2||340|0.6186252338517699|0|1|524|-80.861571|64|35.444615|FRESH PROD FRESH ONIONS|0.0|4|COO YELLOW ONIONS, LRG|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00204665000003|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|427aeaaba02e1b99b4e89cd5d37e375e281ae229|0.31|2015-01-11 15:31:00|1.4102725052409182|2||340|0.6186252338517699|0|1|524|-80.861571|64|35.444615|FRESH PROD FRESH ONIONS|0.0|4|COO YELLOW ONIONS, LRG|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00204665000003|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|46629537307ffea4647f8abbfd002b03e2cf29a8|2.38|2014-10-11 16:02:00|1.4102725052409182|2||340|0.6186252338517699|0|1|529|-80.861571|64|35.444615|FRESH ASPARAGUS|0.27|4|GREEN  ASPARAGUS|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00204080000008|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|390bc2aa1f42dbfbc25fb1f3b155ab15ca1e7bec|4.15|2015-01-31 17:51:00|1.4102725052409182|2||340|0.6186252338517699|0|1|529|-80.861571|64|35.444615|FRESH ASPARAGUS|2.08|4|GREEN  ASPARAGUS|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00204080000008|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|33a207ccf03b63f143e7caabc196301a20ef311e|0.95|2014-10-21 13:19:00|80.86161257435397|2|61300871771|340|35.455082584258413|0|36|99|-80.860108|32|35.500972|LIQUID TEA|0.0|1|ARIZONA DIET PEACH TEA|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|35.472272108304431|00613008719548|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.861571|80.861578596363103|268|1
35.444615|c76b1e70e5c797222588a311aa9c7a35bf0098c1|0.29|2014-09-14 14:10:00|1.4102725052409182|2||340|0.6186252338517699|0|1|502|-80.861571|64|35.444615|FRESH BANANAS|0.0|4|BANANAS, YELLOW|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|e9210c5cd495ac8f729d59cc4ac14294882b9d8b|2.69|2014-09-24 19:18:00|1.4102725052409182|2|7203663996|340|0.6186252338517699|0|1|342|-80.861571|57|35.444615|FRESH MILK|0.0|3|HARRIS TEETER 2%   MILK|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00072036639998|MILK|DAIRY|-80.861571|1.4113006522851637|340|1
35.444615|ffc39f497e3284ad563ba6094a188a3e03dde6a1|39.96|2014-12-15 17:31:00|1.4102725052409182|2|7203661033|340|0.6186252338517699|0|1|666|-80.861571|145|35.444615|PACKAGED COOKED|8.0|12|HT COOKED SHRIMP RING 10OZ|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00072036610331|SHRIMP|SEAFOOD|-80.861571|1.4113006522851637|340|4
35.444615|3daa0a8bd1bf68f1d87af804eda3422033af1d6f|4.99|2014-09-28 15:53:00|1.4102725052409182|2|2840008313|340|0.6186252338517699|0|1|204|-80.861571|31|35.444615|TORTILLA CHIPS|1.0|1|TOSTITOS RSTC FAMILY SIZE|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00028400083133|SNACKS|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.444615|a01abf7bd140f6f2a35e78cf97df3032e33c6ee5|11.98|2014-10-04 12:52:00|1.4102725052409182|2|827411111|340|0.6186252338517699|0|1|55|-80.861571|8|35.444615|REGULAR|0.0|23|REEDS EXTRA GINGER BREW|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00008274444445|CARBONATED BEVERAGES|BEVERAGE|-80.861571|1.4113006522851637|340|2
35.444615|864a4ffb3d80e56d94355e8bb7c1e68b685c5b4e|6.98|2014-11-09 12:57:00|1.4102725052409182|2|75733955555|340|0.6186252338517699|0|1|68|-80.861571|11|35.444615|BARBECUE SAUCES|1.02|1|STICKY FNGR BBQ SC MEMPHIS.|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00757339222220|CONDIMENTS|G1 GROCERY|-80.861571|1.4113006522851637|340|2
35.444615|53edeb74517ce0aa3962590becbb4152d0882d52|12.99|2014-10-01 19:42:00|1.4102725052409182|2|8769229103|340|0.6186252338517699|0|1|458|-80.861571|82|35.444615|CRAFT BEER|0.0|16|SAM ADAMS VARIETY 12PK|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00087692291039|DOMESTIC BEER|BEER|-80.861571|1.4113006522851637|340|1
35.444615|5d7bf7a56bbe3d61dfa16ba874050d0ee8240b26|3.38|2014-09-13 13:37:00|1.4102725052409182|2|7680828008|340|0.6186252338517699|0|1|149|-80.861571|23|35.444615|WHSE PASTA CORE|1.38|1|BARILLA PASTA VEGGIE SPAGHETTI|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00076808004120|PASTA|G1 GROCERY|-80.861571|1.4113006522851637|340|2
35.444615|9b629fafc8f8c5e076d95eb832dde98a07179566|9.99|2014-11-12 18:21:00|1.4102725052409182|2|67058000417|340|0.6186252338517699|0|1|9948|-80.861571|886|35.444615|NFS-PREM-CAB SAUVIGNON|0.0|13|MCMANIS CABERNET|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00670580004172|PREMIUM ($8-$10.99)|WINE|-80.861571|1.4113006522851637|340|1
35.444615|4f37478cd02d724516b3975d97e7573ddf723c92|9.99|2015-01-28 18:18:00|1.4102725052409182|2|8500001819|340|0.6186252338517699|0|1|9955|-80.861571|886|35.444615|NFS-PREM-MALBEC|0.0|13|ALAMOS MENDOZA MALBEC|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00085000018194|PREMIUM ($8-$10.99)|WINE|-80.861571|1.4113006522851637|340|1
35.444615|d2eb9713532c24aea2e33a930baf77bbe7c561c9|2.0|2014-11-24 11:03:00|1.4102725052409182|2|4300000953|340|0.6186252338517699|0|1|272|-80.861571|307|35.444615|TOPPINGS FROZEN|1.01|5|COOL WHIP WHIPPED TOPPING|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00043000009536|DESSERTS FROZEN|FROZEN|-80.861571|1.4113006522851637|340|1
35.444615|f7337612ea89441cf5724eef5d3cfdafd602039a|4.0|2015-01-09 21:47:00|1.4102725052409182|2|66440100025|340|0.6186252338517699|0|1|1165|-80.861571|87|35.444615|NFS-FRESH CONSUMER BUNCH|0.0|9|BUNCH - 3 ST STOCK ASST   JOLO|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00664401000252|FLORAL|FLORAL|-80.861571|1.4113006522851637|340|1
35.444615|7fc81b1344efc261646662535fdcb2f531cc0ccd|3.49|2014-10-02 17:56:00|1.4102725052409182|2|88491212971|340|0.6186252338517699|0|1|81|-80.861571|9|35.444615|RTE CEREAL KIDS|0.0|1|POST PEBBLES FRUITY|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00884912129710|CEREAL|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.444615|4e501ba3823a72fc0cca02c64dac718288ddd7d6|10.88|2014-10-08 19:01:00|1.4102725052409182|2|20596200000|340|0.6186252338517699|0|1|1821|-80.861571|410|35.444615|BH TURKEY|0.0|6|BOARS HEAD MAPLE HONEY TURKEY|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00205962000000|BH MEAT|DELI|-80.861571|1.4113006522851637|340|1
35.444615|9a71693052877aa6a24046b73abcd8d53be3f007|11.87|2014-10-28 19:03:00|1.4102725052409182|2|20596200000|340|0.6186252338517699|0|1|1821|-80.861571|410|35.444615|BH TURKEY|2.16|6|BOARS HEAD MAPLE HONEY TURKEY|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00205962000000|BH MEAT|DELI|-80.861571|1.4113006522851637|340|1
35.444615|76c963de1581d30ec2b0df950d580c288a99dd8c|5.49|2015-02-04 21:18:00|1.4102725052409182|2|4175700109|340|0.6186252338517699|0|1|2018|-80.861571|505|35.444615|PRESSED CHEESE|0.0|6|MINI WHITE CHEDDAR|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00041757018368|SPECIALTY CHEESE|DELI|-80.861571|1.4113006522851637|340|1
35.444615|14df86f7fc469b8b5985fb8e9685b24d906e5118|3.99|2015-01-05 20:42:00|1.4102725052409182|2|7203670998|340|0.6186252338517699|0|1|31|-80.861571|4|35.444615|NON CARBONATED WATER|0.0|1|HT PURIFIED WATER 8 OZ 24PK|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00072036709981|BOTTLED WATER|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.444615|df1efd6cb6442a951d36e4747cc343eb4bdc65b6|3.49|2014-11-24 18:10:00|1.4102725052409182|2|9235243007|340|0.6186252338517699|0|1|6471|-80.861571|1558|35.444615|PLASTIC UTENSILS|0.0|18|SENS ASST CUTLERY WASABI GREEN|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00092352430222|PARTY NAPKINS/PLATES|GM|-80.861571|1.4113006522851637|340|1
35.444615|3fd93970ec33b137ca89cfe6b9f4ae4f662f3078|4.38|2014-12-20 18:23:00|1.4102725052409182|2|4900005010|340|0.6186252338517699|0|1|55|-80.861571|8|35.444615|REGULAR|1.88|23|SCHWEPPES GINGERALE 2LTR|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00078000206463|CARBONATED BEVERAGES|BEVERAGE|-80.861571|1.4113006522851637|340|2
35.444615|4bd857fd337427cdbe1066acb1ff71fa3221f243|3.49|2014-11-24 11:04:00|1.4102725052409182|2|7797508005|340|0.6186252338517699|0|1|202|-80.861571|31|35.444615|PRETZELS|0.3|1|SOH SNAPS 20% BONUS PK|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00077975091395|SNACKS|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.444615|c6d6a89b07e1675983d210c509d6b1f86a1c8b7c|3.99|2014-12-03 13:47:00|80.86161257435397|2|7203697777|340|35.455082584258413|0|36|31|-80.860108|4|35.500972|NON CARBONATED WATER|1.49|1|(U) HT PURIFIED WATER 24 PK|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|35.472272108304431|00072036977779|BOTTLED WATER|G1 GROCERY|-80.861571|80.861578596363103|268|1
35.444615|85a3f2d15589dde9ba415e2c8ffbc498f1ed7a19|3.15|2014-11-24 11:08:00|1.4102725052409182|2|7225003706|340|0.6186252338517699|0|1|1026|-80.861571|162|35.444615|WHEAT|0.0|7|NATOWN HONEYWHEAT BRD|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00072250037068|SLICED BREAD|COMMERCIAL BAKERY|-80.861571|1.4113006522851637|340|1
35.444615|1422db2aafdfd0117647828e57bf8a8bc25d6a1f|1.99|2014-11-10 17:26:00|1.4102725052409182|2|1360002005|340|0.6186252338517699|0|1|221|-80.861571|34|35.444615|SALT SALT SUBSTITUTES|0.6|1|DIAMOND CRYSTAL FINE SEA SALT|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00013600020064|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.444615|7af5bdf22d645448de101c40b9a4b9829669848e|11.99|2014-11-03 11:51:00|1.4102725052409182|2|20595400000|340|0.6186252338517699|0|1|1823|-80.861571|410|35.444615|BH HAM|2.0|6|BOARS HEAD TRIO|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00205954000001|BH MEAT|DELI|-80.861571|1.4113006522851637|340|1
35.444615|8e268bc4c2e1170c9dc796d45014eb5ea0f13f11|2.99|2014-09-30 11:35:00|1.4102725052409182|2|7203698526|340|0.6186252338517699|0|1|201|-80.861571|31|35.444615|POTATO CHIPS|0.49|1|HT TRADER KETTLE CHIP SALT VIN|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00072036985286|SNACKS|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.444615|e58d0f57650ee072ee09d3799ef38056daf8642a|4.29|2014-10-01 19:45:00|1.4102725052409182|2|7203670353|340|0.6186252338517699|0|1|442|-80.861571|76|35.444615|NFS-COOKING-STORAGE BAGS|0.0|1|YH RESEAL DBL ZIP STORAGE GAL|99bd7a3f2d7304bdb975556c796c3588012430b7|0.7232849203347611|0.61833652052202714|00072036703545|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.667941|d31a6e6d74609691382828d9be48cfee06428c82|2.99|2015-02-11 21:45:00|1.4057311447477159|4|8186422116|178|0.6225230078570788|0|52|583|-80.497332|136|35.667941|NUTS|0.99|4|SALTED PEANUTS IN-SHELL|99f04c72734d00aa457d1a2e5f25c20c74aa380b|6.448336988341629|0.6209993146566879|00081864221169|OTHER MERCHANDISE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|02ca80f3b916a2b030830622a852c9d35994e0ff|2.99|2015-02-16 16:44:00|1.4057311447477159|4|8186422116|178|0.6225230078570788|0|52|583|-80.497332|136|35.667941|NUTS|0.99|4|SALTED PEANUTS IN-SHELL|99f04c72734d00aa457d1a2e5f25c20c74aa380b|6.448336988341629|0.6209993146566879|00081864221169|OTHER MERCHANDISE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|7417e5458de355697122ecf9fe27e7d4535f9394|5.78|2014-12-04 20:24:00|1.4057311447477159|4|7203663102|178|0.6225230078570788|0|52|339|-80.497332|57|35.667941|EGGNOGS/DRINKS|1.78|3|I/O HARRIS TEETER EGG NOG|99f04c72734d00aa457d1a2e5f25c20c74aa380b|6.448336988341629|0.6209993146566879|00072036631022|MILK|DAIRY|-80.497332|1.4049434824709919|178|2
35.667941|1b83ee38c80d90b58c2c2a3ddb340423aeb21256|2.89|2014-11-20 20:28:00|1.4057311447477159|4|7203663102|178|0.6225230078570788|0|52|339|-80.497332|57|35.667941|EGGNOGS/DRINKS|0.39|3|I/O HARRIS TEETER EGG NOG|99f04c72734d00aa457d1a2e5f25c20c74aa380b|6.448336988341629|0.6209993146566879|00072036631022|MILK|DAIRY|-80.497332|1.4049434824709919|178|1
35.667941|415e401cd71a53b63c0b4f2505b20731de95c5d9|5.78|2014-11-23 20:37:00|1.4057311447477159|4|7203663102|178|0.6225230078570788|0|52|339|-80.497332|57|35.667941|EGGNOGS/DRINKS|0.78|3|I/O HARRIS TEETER EGG NOG|99f04c72734d00aa457d1a2e5f25c20c74aa380b|6.448336988341629|0.6209993146566879|00072036631022|MILK|DAIRY|-80.497332|1.4049434824709919|178|2
35.667941|85de9a56add60d974465b3d4792ddaef3852e1a9|5.98|2015-01-19 19:15:00|1.4057311447477159|4|8186420216|178|0.6225230078570788|0|52|583|-80.497332|136|35.667941|NUTS|1.98|4|ROASTED PEANUTS IN-SHELL|99f04c72734d00aa457d1a2e5f25c20c74aa380b|6.448336988341629|0.6209993146566879|00081864222166|OTHER MERCHANDISE|PRODUCE|-80.497332|1.4049434824709919|178|2
35.667941|515cad73e93315194846545ec8d2174875dd66ac|0.97|2014-11-25 19:02:00|1.4057311447477159|4||178|0.6225230078570788|0|52|535|-80.497332|64|35.667941|FRESH GREENS|0.0|4|COO TURNIP GREENS, BULK|99f04c72734d00aa457d1a2e5f25c20c74aa380b|6.448336988341629|0.6209993146566879|00204619000004|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|77c9b9b0cb2bc3f80630144588e107616d1d9e29|1.33|2014-11-17 20:53:00|1.4057311447477159|4||178|0.6225230078570788|0|52|535|-80.497332|64|35.667941|FRESH GREENS|0.0|4|COO TURNIP GREENS, BULK|99f04c72734d00aa457d1a2e5f25c20c74aa380b|6.448336988341629|0.6209993146566879|00204619000004|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|d5d0ae1a99b4482f1aa5983b9386f982f80af598|1.06|2014-09-11 22:31:00|1.4057311447477159|4||178|0.6225230078570788|0|52|535|-80.497332|64|35.667941|FRESH GREENS|0.0|4|COO TURNIP GREENS, BULK|99f04c72734d00aa457d1a2e5f25c20c74aa380b|6.448336988341629|0.6209993146566879|00204619000004|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|d352613a885d01bf72bd5730c52c2655c8fc341e|3.84|2015-01-28 16:33:00|1.4057311447477159|4||178|0.6225230078570788|0|52|558|-80.497332|64|35.667941|SPECIALTY-VEGETABLES|0.0|4|COO HORSERADISH ROOT|99f04c72734d00aa457d1a2e5f25c20c74aa380b|6.448336988341629|0.6209993146566879|00204625000005|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|ea9c791140792d9b7cda2791f89628734baa3989|18.46|2015-01-31 15:17:00|1.4057311447477159|4||178|0.6225230078570788|0|52|503|-80.497332|64|35.667941|FRESH GRAPES|2.64|4|RED GRAPES,SEEDLESS 12/16|99f04c72734d00aa457d1a2e5f25c20c74aa380b|6.448336988341629|0.6209993146566879|00204023000003|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|c4d418dc72e874f841594326c6bd3d3c0656867d|4.99|2014-09-23 18:53:00|1.4057311447477159|4|7203697885|178|0.6225230078570788|0|52|200|-80.497332|31|35.667941|MICROWAVE POPCORN|0.0|1|HTN ORGANIC POPCORN YELLOW|99f04c72734d00aa457d1a2e5f25c20c74aa380b|6.448336988341629|0.6209993146566879|00072036978851|SNACKS|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|c3439ed8649c21b8ba0795e9e34dcd8b8d6c9d9b|3.49|2014-11-22 19:00:00|1.4057311447477159|4|85225100001|178|0.6225230078570788|0|52|339|-80.497332|57|35.667941|EGGNOGS/DRINKS|0.5|3|I/O SUTHRN COMF EGG NOG|99f04c72734d00aa457d1a2e5f25c20c74aa380b|6.448336988341629|0.6209993146566879|00852251000014|MILK|DAIRY|-80.497332|1.4049434824709919|178|1
35.667941|96256af271d7d572775beda51d27a447581dc090|3.34|2015-02-20 19:43:00|1.4057311447477159|4||178|0.6225230078570788|0|52|523|-80.497332|64|35.667941|FRESH POTATOES|0.68|4|COO SWEET POTATOES, BULK|99f04c72734d00aa457d1a2e5f25c20c74aa380b|6.448336988341629|0.6209993146566879|00204091000004|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|fc19da9e8fa7f3bf871075fe9f6463904aaacad8|1.59|2014-12-14 19:35:00|1.4057311447477159|4|6661300009|178|0.6225230078570788|0|52|191|-80.497332|29|35.667941|REMAINING SEAFOOD-CANNED|0.34|1|BRUNSWICK SARDINES IN WATER|99f04c72734d00aa457d1a2e5f25c20c74aa380b|6.448336988341629|0.6209993146566879|00066613000097|SEAFOOD-CANNED|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|5cc65bc763441680d7813af1b5363a2e371da1b8|0.99|2015-02-08 18:26:00|1.4057311447477159|4||178|0.6225230078570788|0|52|535|-80.497332|64|35.667941|FRESH GREENS|0.0|4|COLLARD GREENS, BUN (RPC)|99f04c72734d00aa457d1a2e5f25c20c74aa380b|6.448336988341629|0.6209993146566879|00204614000009|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|0b23b35d968275d69769a4f4d8b04ef1af5da5e1|1.99|2014-12-31 18:06:00|1.4057311447477159|4||178|0.6225230078570788|0|52|535|-80.497332|64|35.667941|FRESH GREENS|1.0|4|COLLARD GREENS, BUN (RPC)|99f04c72734d00aa457d1a2e5f25c20c74aa380b|6.448336988341629|0.6209993146566879|00204614000009|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|835f7618bad5ff0d3d107d69b3819c25c12cb6a0|7.98|2015-03-08 18:25:00|1.4057311447477159|4|7203663061|178|0.6225230078570788|0|52|364|-80.497332|55|35.667941|ORGANIC AND CF EGGS|0.0|3|HTO ORGANIC GRD A LARGE EGG BR|99f04c72734d00aa457d1a2e5f25c20c74aa380b|6.448336988341629|0.6209993146566879|00072036630612|EGGS FRESH|DAIRY|-80.497332|1.4049434824709919|178|2
35.667941|734967ed4a911d0cf9e6e522cd26ab24cf14c7c2|7.98|2014-09-19 18:53:00|1.4057311447477159|4|7203663061|178|0.6225230078570788|0|52|364|-80.497332|55|35.667941|ORGANIC AND CF EGGS|0.0|3|HTO ORGANIC GRD A LARGE EGG BR|99f04c72734d00aa457d1a2e5f25c20c74aa380b|6.448336988341629|0.6209993146566879|00072036630612|EGGS FRESH|DAIRY|-80.497332|1.4049434824709919|178|2
35.667941|6e2e476d33363cb00e63fe355f836612d7bc0128|3.99|2015-02-27 14:10:00|1.4057311447477159|4|7203663061|178|0.6225230078570788|0|52|364|-80.497332|55|35.667941|ORGANIC AND CF EGGS|0.0|3|HTO ORGANIC GRD A LARGE EGG BR|99f04c72734d00aa457d1a2e5f25c20c74aa380b|6.448336988341629|0.6209993146566879|00072036630612|EGGS FRESH|DAIRY|-80.497332|1.4049434824709919|178|1
35.372142|ad056a6f84b66e765554c5c6a0acd067018ddd6a|14.99|2014-11-08 20:51:00|80.779636304526477|3|8992488007|122|35.396821757261272|0|17|455|-80.784334|82|35.384824|DOMESTIC PREMIUM 12PK&>|0.0|16|YUENGLING LAGER 24PK CANS|9a5f1aa555e720c95d43951b8c344ec1127592ac|1.705311640594015|35.392509581117899|00089924880073|DOMESTIC BEER|BEER|-80.782849|80.782852783551135|476|1
35.372142|8a663b4062591e8a98759d997bf45b1261c1ea8f|14.99|2015-01-12 17:25:00|80.779636304526477|3|8992488007|122|35.396821752305151|0|17|455|-80.746334|82|35.41832|DOMESTIC PREMIUM 12PK&>|0.0|16|YUENGLING LAGER 24PK CANS|9a5f1aa555e720c95d43951b8c344ec1127592ac|1.705311640594015|35.392509581117899|00089924880073|DOMESTIC BEER|BEER|-80.782849|80.782868553894019|190|1
35.372142|2e534c6a3fb3f409c170df125e1bc3b72404d814|15.99|2014-09-28 18:22:00|1.4102725052409182|3|8992488007|122|0.617360341382972|0|1|455|-80.782849|82|35.372142|DOMESTIC PREMIUM 12PK&>|0.0|16|YUENGLING LAGER 24PK CANS|9a5f1aa555e720c95d43951b8c344ec1127592ac|1.705311640594015|0.61833652052202714|00089924880073|DOMESTIC BEER|BEER|-80.782849|1.4099266941914086|122|1
35.372142|f1163d4f33fb940cdbeb9740a49e053d030b5a3f|9.13|2014-11-24 20:53:00|80.779636304526477|3||122|35.396821757261272|0|17|1405|-80.784334|21|35.384824|BULK NUTS|0.0|1|CAPITOL MIX II NATURAL #340|9a5f1aa555e720c95d43951b8c344ec1127592ac|1.705311640594015|35.392509581117899|00094184100519|NUTS|G1 GROCERY|-80.782849|80.782852783551135|476|1
35.372142|8ccd8ead21c5ca6880aa5ca8ac52f4d574702241|6.39|2014-12-26 13:38:00|80.779636304526477|3|1030033602|122|35.396821757261272|0|17|1148|-80.784334|21|35.384824|ALMONDS|2.4|1|EMERALD DRY ROASTED ALMONDS|9a5f1aa555e720c95d43951b8c344ec1127592ac|1.705311640594015|35.392509581117899|00010300336020|NUTS|G1 GROCERY|-80.782849|80.782852783551135|476|1
35.372142|732e0caeb401bd7bfeb8915453ebf9445dd2899a|8.99|2014-10-10 21:58:00|80.779636304526477|3|85877000244|122|35.396821757261272|0|17|458|-80.784334|82|35.384824|CRAFT BEER|0.0|16|OMB COPPER 12OZ 6PACK|9a5f1aa555e720c95d43951b8c344ec1127592ac|1.705311640594015|35.392509581117899|00858770002447|DOMESTIC BEER|BEER|-80.782849|80.782852783551135|476|1
35.372142|01055557dcc711d2db18d9a9e88858de08827e10|8.99|2015-02-25 18:27:00|1.4102725052409182|3|7289482424|122|0.617360341382972|0|1|5504|-80.782849|1504|35.372142|TOWELS|0.0|18|3PK KITCHEN TOWEL MOCHA|9a5f1aa555e720c95d43951b8c344ec1127592ac|1.705311640594015|0.61833652052202714|00072894824611|DOMESTICS|GM|-80.782849|1.4099266941914086|122|1
35.372142|81d7f36dec3926b2f37413a6bbc1cec678a939df|9.99|2014-11-04 19:58:00|80.779636304526477|3|8158401310|122|35.396821757261272|0|17|9959|-80.784334|887|35.384824|NFS-S/PREM-CHARDONNAY|0.0|13|CB-K. JACKSON V.R. CHARDONNAY|9a5f1aa555e720c95d43951b8c344ec1127592ac|1.705311640594015|35.392509581117899|00081584013105|SUPER PREMIUM ($11-$14.99)|WINE|-80.782849|80.782852783551135|476|1
35.372142|25d135fc5970370d0c618000e360e02a47d49b1a|3.99|2014-11-23 14:53:00|1.4102725052409182|3|4300095117|122|0.617360341382972|0|1|209|-80.782849|20|35.372142|POWDERED SOFT DRINKS|0.0|1|COUNTRY TIME LEMONADE (8QT)|9a5f1aa555e720c95d43951b8c344ec1127592ac|1.705311640594015|0.61833652052202714|00043000951170|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|c5cd0e6be2193e66f66fd40e64d8eb618fcb1e9a|4.49|2015-01-18 16:14:00|80.779636304526477|3|74759930652|122|35.396821757261272|0|17|62|-80.784334|7|35.384824|SPECIALTY BAR/BOX CHOCOLATE|0.0|1|GHIR MILK CHOC CARAMEL SQUARES|9a5f1aa555e720c95d43951b8c344ec1127592ac|1.705311640594015|35.392509581117899|00747599306518|CANDY|G1 GROCERY|-80.782849|80.782852783551135|476|1
35.372142|f11c9b7fce011203306f416e1232820958c7eeb9|1.97|2015-02-09 14:44:00|80.779636304526477|3|7203608134|122|35.396821753810428|0|17|82|-80.780702|11|35.318911|VINEGAR|0.0|1|HT VINEGAR WHITE DISTILLED 64|9a5f1aa555e720c95d43951b8c344ec1127592ac|1.705311640594015|35.392509581117899|00072036081346|CONDIMENTS|G1 GROCERY|-80.782849|80.782865449125907|167|1
35.372142|0c7f4f086d1f9efaa63bdaf2f70f182274c9230a|3.34|2015-02-17 14:55:00|80.779636304526477|3|7203610087|122|35.396821753810428|0|17|90|-80.780702|13|35.318911|SNACK CRACKERS|1.67|1|HT THIN WHEAT CRACKERS|9a5f1aa555e720c95d43951b8c344ec1127592ac|1.705311640594015|35.392509581117899|00072036100849|CRACKERS|G1 GROCERY|-80.782849|80.782865449125907|167|1
35.372142|28782d19560740865a24d7b82ef239d6154e861f|5.58|2015-01-26 16:15:00|80.779636304526477|3|5100014880|122|35.396821753810428|0|17|1499|-80.780702|33|35.318911|RTS MICROWAVE|0.0|1|CHUNKY MW PUB CHICKEN POT PIE|9a5f1aa555e720c95d43951b8c344ec1127592ac|1.705311640594015|35.392509581117899|00051000215864|SOUP|G1 GROCERY|-80.782849|80.782865449125907|167|2
35.372142|056e1c8ecd5d0ddadf797267dc84320b54b18ec8|19.99|2015-01-11 17:37:00|80.779636304526477|3|85122400201|122|35.396821757261272|0|17|458|-80.784334|82|35.384824|CRAFT BEER|0.0|16|REDOAK AMBER LAGER BEER 12PK|9a5f1aa555e720c95d43951b8c344ec1127592ac|1.705311640594015|35.392509581117899|00851224002017|DOMESTIC BEER|BEER|-80.782849|80.782852783551135|476|1
35.372142|871922c4291ea8e91aa170412a7847d031ef04a1|1.99|2014-12-22 16:42:00|1.4102725052409182|3|7127923100|122|0.617360341382972|0|1|555|-80.782849|64|35.372142|PACKAGED SALADS|0.0|4|F.E. BABY SPRING SALAD MIX|9a5f1aa555e720c95d43951b8c344ec1127592ac|1.705311640594015|0.61833652052202714|00071279231006|FRESH PRODUCE|PRODUCE|-80.782849|1.4099266941914086|122|1
35.372142|73ae6ab14228efd453b663f1401ceddbcd8ee83e|8.97|2015-01-20 22:10:00|80.779636304526477|3|63888200203|122|35.396821752305151|0|17|247|-80.746334|39|35.41832|VEGETABLES-FLANKER|0.3|1|FARMERS MKT ORG PUMPKIN|9a5f1aa555e720c95d43951b8c344ec1127592ac|1.705311640594015|35.392509581117899|00638882002005|VEGETABLES-CAN/JAR|G1 GROCERY|-80.782849|80.782868553894019|190|3
35.372142|4505b0116f08047042395bc76b03a70626a07b1d|9.99|2014-11-08 16:36:00|1.4102725052409182|3|8600387388|122|0.617360341382972|0|1|9934|-80.782849|885|35.372142|NFS POP CHARDONNAY|0.0|13|CB-WOODBRIDGE CHARDONNAY 1.5L|9a5f1aa555e720c95d43951b8c344ec1127592ac|1.705311640594015|0.61833652052202714|00086003873889|POPULAR (4-$7.99)|WINE|-80.782849|1.4099266941914086|122|1
35.372142|edc90768fd3327af8621f0f723ca055d734bb17c|9.99|2014-11-05 19:18:00|80.779636304526477|3|8600387388|122|35.396821757261272|0|17|9934|-80.784334|885|35.384824|NFS POP CHARDONNAY|0.0|13|CB-WOODBRIDGE CHARDONNAY 1.5L|9a5f1aa555e720c95d43951b8c344ec1127592ac|1.705311640594015|35.392509581117899|00086003873889|POPULAR (4-$7.99)|WINE|-80.782849|80.782852783551135|476|1
35.372142|522b9bfba5927f0f7be1cfeab2a302470e6f88f4|9.99|2014-09-14 17:33:00|80.779636304526477|3|1235407144|122|35.396821757261272|0|17|9957|-80.784334|886|35.384824|NFS-PREM-OTHER RED|0.0|13|PENFOLDS KOONUNGA SHIRAZ CAB|9a5f1aa555e720c95d43951b8c344ec1127592ac|1.705311640594015|35.392509581117899|00012354071445|PREMIUM ($8-$10.99)|WINE|-80.782849|80.782852783551135|476|1
35.372142|1bb1cc592875bbd54fb4de1e9987951e37fe2fb6|7.49|2014-12-22 14:23:00|80.779636304526477|3|1124620855|122|35.396821757261272|0|17|126|-80.784334|19|35.384824|PRESERVES/MARMALADE|0.0|1|D*ROTHS HOT PEP PEACH PRESERVE|9a5f1aa555e720c95d43951b8c344ec1127592ac|1.705311640594015|35.392509581117899|00011246208556|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.782849|80.782852783551135|476|1
35.372142|ee7fea40997ffdea19a6a8cb6c03f9b5242fdef2|3.95|2014-10-26 18:06:00|80.779636304526477|3||122|35.396821757261272|0|17|1405|-80.784334|21|35.384824|BULK NUTS|0.0|1|CHECKMATE MIX #309|9a5f1aa555e720c95d43951b8c344ec1127592ac|1.705311640594015|35.392509581117899|00094184110082|NUTS|G1 GROCERY|-80.782849|80.782852783551135|476|1
35.372142|81ab13d6155df014fecb70b189fba7c6793b2f58|1.69|2014-12-04 20:45:00|80.779636304526477|3|4900000044|122|35.396821757261272|0|17|54|-80.784334|8|35.384824|DIET|0.0|23|CB DIET COKE CONTOUR 20 OZ NR|9a5f1aa555e720c95d43951b8c344ec1127592ac|1.705311640594015|35.392509581117899|00049000000450|CARBONATED BEVERAGES|BEVERAGE|-80.782849|80.782852783551135|476|1
35.372142|81615191e395263dff3108eb0c39482014a2e0b5|8.49|2014-12-22 17:12:00|1.4102725052409182|3|7675320015|122|0.617360341382972|0|1|5879|-80.782849|1538|35.372142|FOOD PREPARATION|0.0|18|GOODCOOK MEAT TENDRZER 20015|9a5f1aa555e720c95d43951b8c344ec1127592ac|1.705311640594015|0.61833652052202714|00076753200158|KITCHEN GADGETS|GM|-80.782849|1.4099266941914086|122|1
35.667941|9ed8e70401cd998b177a3b97984964ae629dd954|5.79|2014-11-27 12:09:00|1.4057311447477159|2|2100060260|178|0.6225230078570788|0|52|315|-80.497332|52|35.667941|CHEESE-PROCESSED-SLICED|0.0|3|KRAFT DELI DELUXE SLICES|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00021000602605|CHEESE|DAIRY|-80.497332|1.4049434824709919|178|1
35.667941|7d4c2637335a522a2282695705db2ea784fc9796|0.99|2014-12-04 14:53:00|1.4057311447477159|2|2700038815|178|0.6225230078570788|0|52|257|-80.497332|39|35.667941|TOMATOES|0.0|1|HUNTS TOMATO PASTE BSL GAR ORE|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00027000388235|VEGETABLES-CAN/JAR|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|59ffc84f6315c29ce301b571b2726ec396e7de8e|10.79|2015-02-02 16:32:00|1.4057311447477159|2|2100060260|178|0.6225230078570788|0|52|315|-80.497332|52|35.667941|CHEESE-PROCESSED-SLICED|0.0|3|KRAFT DELI DELUXE SLICES|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00021000602605|CHEESE|DAIRY|-80.497332|1.4049434824709919|178|2
35.667941|5dedacea88651576f3c0302de2c2a3a132c20000|17.45|2014-10-20 16:23:00|1.4057311447477159|2|20138900000|178|0.6225230078570788|0|52|296|-80.497332|49|35.667941|RANCHER BEEF|4.85|2|BEEF TENDERLOIN FILET MIGNON|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00201389000005|BEEF|MEAT|-80.497332|1.4049434824709919|178|1
35.667941|e42d219d97ba636cd4d8376652ea97c90d69f4c8|14.57|2015-02-27 12:17:00|1.4057311447477159|2|20138900000|178|0.6225230078570788|0|52|296|-80.497332|49|35.667941|RANCHER BEEF|4.05|2|BEEF TENDERLOIN FILET MIGNON|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00201389000005|BEEF|MEAT|-80.497332|1.4049434824709919|178|1
35.667941|aa9ecadf0005d7ee68be16b0202f2a98a78b4512|2.86|2014-12-23 10:58:00|1.4057311447477159|2||178|0.6225230078570788|0|52|522|-80.497332|64|35.667941|FRESH TOMATOES|0.0|4|COO GREEN TOMATILLOS|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00204801000003|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|12f05961c707b4cb95532096751283625205f863|9.72|2015-01-23 15:27:00|1.4057311447477159|2|20193000000|178|0.6225230078570788|0|52|299|-80.497332|49|35.667941|ANGUS BEEF|0.0|2|ANGUS BEEF CHUCK TENDER ROAST|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00201930000003|BEEF|MEAT|-80.497332|1.4049434824709919|178|1
35.667941|454c3ad916340549195159720f9c47d2b549ffbd|15.29|2014-12-21 18:39:00|1.4057311447477159|2|20138900000|178|0.6225230078570788|0|52|296|-80.497332|49|35.667941|RANCHER BEEF|4.25|2|BEEF TENDERLOIN FILET MIGNON|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00201389000005|BEEF|MEAT|-80.497332|1.4049434824709919|178|1
35.667941|990ef82a0b8d495594dee794a46f00dd1f7ab36e|1.99|2014-12-27 16:31:00|80.497482303704658|2|3760023785|178|35.708501930169568|0|6|175|-80.66939|27|35.28326|CANNED MEATS|0.0|1|HORMEL CHILI NO BEANS|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|35.699188602026126|00037600237857|PREPARED FOODS-RTS|G1 GROCERY|-80.497332|80.497571076724597|46|1
35.667941|0f00b914cbf87f120af70a6ea8d2ad3efc6f7d01|11.99|2014-09-19 17:32:00|1.4057311447477159|2|78535710062|178|0.6225230078570788|0|52|35|-80.497332|10|35.667941|PREMIUM WHOLE BEAN|4.0|1|PEET'S SUMATRA WB|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00785357100909|COFFEE|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|020383bfaf19c6de2aa215842b8740b9480494b5|11.99|2014-10-24 14:55:00|1.4057311447477159|2|78535710062|178|0.6225230078570788|0|52|35|-80.497332|10|35.667941|PREMIUM WHOLE BEAN|4.0|1|PEET'S SUMATRA WB|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00785357100909|COFFEE|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|0dfe3320384dd13bdc1d0fcb5ebf05f550244d9f|2.29|2014-09-23 14:28:00|1.4057311447477159|2|930000044|178|0.6225230078570788|0|52|163|-80.497332|25|35.667941|RELISHES|0.0|1|MT OLV RELISH NO SUGAR|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00009300001069|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|34d577ea0c6bc081fe2a48d1b6a666763d8c20a1|2.19|2015-03-06 13:28:00|1.4057311447477159|2|930000044|178|0.6225230078570788|0|52|163|-80.497332|25|35.667941|RELISHES|0.0|1|MT OLV RELISH NO SUGAR|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00009300001069|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|e60605bcd3b2d5420df58b9073d0fe4cdba3fa06|4.99|2015-02-20 18:38:00|1.4057311447477159|2|78142152480|178|0.6225230078570788|0|52|1601|-80.497332|371|35.667941|BRANDED BREAD|1.5|14|LA BREA THREE CHEESE SEMOLINA|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00781421524800|BREAD|BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|cefd29f59e782e39ac4c79a54922efc892d167af|4.99|2015-01-16 14:10:00|1.4057311447477159|2|78142152480|178|0.6225230078570788|0|52|1601|-80.497332|371|35.667941|BRANDED BREAD|0.0|14|LA BREA THREE CHEESE SEMOLINA|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00781421524800|BREAD|BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|611e2e9865bf386c398b3af01ee8a3aa4af4d7f4|4.99|2014-10-29 19:17:00|1.4057311447477159|2|78142152480|178|0.6225230078570788|0|52|1601|-80.497332|371|35.667941|BRANDED BREAD|0.0|14|LA BREA THREE CHEESE SEMOLINA|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00781421524800|BREAD|BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|bb0070674ad4ed8095812f1b197a102a4a503b53|3.98|2014-10-13 13:33:00|1.4057311447477159|2||178|0.6225230078570788|0|52|561|-80.497332|64|35.667941|FR PROD ORGANIC PRODUCE|0.0|4|ORG CILANTRO|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00789622530019|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|2
35.667941|608af576ccff75f703fe0313838766265d29ed39|4.99|2014-10-02 18:02:00|1.4057311447477159|2|78142152480|178|0.6225230078570788|0|52|1601|-80.497332|371|35.667941|BRANDED BREAD|0.0|14|LA BREA THREE CHEESE SEMOLINA|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00781421524800|BREAD|BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|12bec72190165bba2c9b2df0decbfbd19de1a4fa|1.99|2015-01-19 13:35:00|1.4057311447477159|2||178|0.6225230078570788|0|52|561|-80.497332|64|35.667941|FR PROD ORGANIC PRODUCE|0.49|4|ORG CILANTRO|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00789622530019|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|ff742da6f9844b546136fc6ee35461a0d4883902|1.94|2015-01-24 19:11:00|1.4057311447477159|2|7203698757|178|0.6225230078570788|0|52|31|-80.497332|4|35.667941|NON CARBONATED WATER|0.0|1|HT PURIFIED WATER|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00072036987570|BOTTLED WATER|G1 GROCERY|-80.497332|1.4049434824709919|178|2
35.667941|bb236379696b34d87a8b352ce8241cf7c9a88376|1.94|2015-02-25 10:35:00|1.4057311447477159|2|7203698757|178|0.6225230078570788|0|52|31|-80.497332|4|35.667941|NON CARBONATED WATER|0.0|1|HT PURIFIED WATER|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00072036987570|BOTTLED WATER|G1 GROCERY|-80.497332|1.4049434824709919|178|2
35.667941|3bde8c9c0e1e71a2b5698e185ef90cde87c7aee3|1.94|2014-09-21 16:06:00|1.4057311447477159|2|7203698757|178|0.6225230078570788|0|52|31|-80.497332|4|35.667941|NON CARBONATED WATER|0.0|1|HT PURIFIED WATER|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00072036987570|BOTTLED WATER|G1 GROCERY|-80.497332|1.4049434824709919|178|2
35.667941|a42784a3f1486ceccf2400a90c902ff1c70d78ee|1.94|2014-11-28 15:39:00|1.4057311447477159|2|7203698757|178|0.6225230078570788|0|52|31|-80.497332|4|35.667941|NON CARBONATED WATER|0.0|1|HT PURIFIED WATER|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00072036987570|BOTTLED WATER|G1 GROCERY|-80.497332|1.4049434824709919|178|2
35.667941|773dfea650d6d33a0fcb857454cb354dc9202303|9.79|2014-11-12 19:19:00|1.4057311447477159|2|9955536128|178|0.6225230078570788|0|52|35|-80.497332|10|35.667941|PREMIUM WHOLE BEAN|0.0|1|NEWMAN'S ORG/COLOMBIAN W/B|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00099555361285|COFFEE|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|a6a7451c7e7786763d73216abeafc7240687717a|2.99|2014-11-12 21:21:00|1.4057311447477159|2|9396600091|178|0.6225230078570788|0|52|345|-80.497332|57|35.667941|ORGANIC MILK|0.0|3|ORGANIC VALLEY 2% LOW FAT MILK|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00093966000214|MILK|DAIRY|-80.497332|1.4049434824709919|178|1
35.667941|c8fe5dc443ae31fc04ca470ca36c7f02c52c9d21|3.59|2014-12-21 10:35:00|80.497482303704658|2|7225004319|178|35.708501930169568|0|6|1026|-80.66939|162|35.28326|WHEAT|0.0|7|NATOWN 100% WHEAT W/HNY  BRD|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|35.699188602026126|00072250043199|SLICED BREAD|COMMERCIAL BAKERY|-80.497332|80.497571076724597|46|1
35.667941|d34f0aebfb9313dbde47cda163f3902538cb5880|1.99|2014-11-18 10:46:00|1.4057311447477159|2|7203676415|178|0.6225230078570788|0|52|1465|-80.497332|42|35.667941|ORGANIC FROZEN FRUIT|0.0|5|HTO ORGANIC WHOLE MXED BERRIES|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00072036763846|FROZEN FRUIT|FROZEN|-80.497332|1.4049434824709919|178|1
35.667941|dcb38f367fae5734ef7b33aafc834f2a7cab5947|10.8|2015-02-06 12:40:00|1.4057311447477159|2|27085500000|178|0.6225230078570788|0|52|973|-80.497332|201|35.667941|FRESH PERDUE CHICKEN|0.0|2|PERDUE OVEN STUFFER ROASTER|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00270855000009|POULTRY|MEAT|-80.497332|1.4049434824709919|178|1
35.667941|d9b04291a366da42d5eed22030bb98982dac19a1|14.99|2015-01-08 12:43:00|1.4057311447477159|2|8500002028|178|0.6225230078570788|0|52|9957|-80.497332|886|35.667941|NFS-PREM-OTHER RED|0.0|13|BAREFOOT RED MOSCATO 1.5L|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00085000020289|PREMIUM ($8-$10.99)|WINE|-80.497332|1.4049434824709919|178|2
35.667941|9ef0bf63dde5d88baf11f1f02c31d4993e9ff79c|4.99|2014-12-20 08:23:00|80.497482303704658|2|1600027528|178|35.708501930169568|0|6|74|-80.66939|9|35.28326|RTE CEREAL ALL FAMILY|0.0|1|GM CHEERIOS 18 OZ|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|35.699188602026126|00016000275287|CEREAL|G1 GROCERY|-80.497332|80.497571076724597|46|1
35.667941|a825d833d7a68f1ae183d72095afdb84f0a76889|12.99|2014-12-26 17:42:00|1.4057311447477159|2|1440081400|178|0.6225230078570788|0|52|477|-80.497332|81|35.667941|NFS-CANNING JARS/LIDS|2.0|1|BALL CRYSTAL JELLY JARS 12OZ|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00014400814006|CANNING|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|99e7631ba0770fde3ee8fc45d344a426ac6f0221|4.19|2015-02-05 14:47:00|1.4057311447477159|2|4812110208|178|0.6225230078570788|0|52|1037|-80.497332|164|35.667941|ENGLISH MUFFINS|0.0|7|THOMAS ENG MUFFN ORIG 6 PK PP|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00048121102081|BREAKFAST|COMMERCIAL BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|9e04b7e430e6c58e1d8a5aecdc5efbd9fb7faff6|2.19|2015-01-22 13:07:00|1.4057311447477159|2|5410001870|178|0.6225230078570788|0|52|163|-80.497332|25|35.667941|RELISHES|1.1|1|VLASIC RELISH SWEET|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00054100018700|PICKLES/OLIVES/RELISHES|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|b336c7f93afe1ffbd7dac7182c0bcd8afa055a55|1.0|2014-11-04 16:17:00|1.4057311447477159|2|78352054321|178|0.6225230078570788|0|52|8598|-80.497332|1792|35.667941|NEWSPAPERS|0.0|18|DAILY  CHARLOTTE OBSERVER|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00783520543218|NEWSPAPERS|GM|-80.497332|1.4049434824709919|178|1
35.667941|8c6cb36c2d509aafddfae4a777417b52bfbfbe44|2.58|2014-11-22 15:25:00|1.4057311447477159|2|2904900602|178|0.6225230078570788|0|52|5619|-80.497332|1512|35.667941|RODENT/INSECT CONTROL|0.0|18|CM WOODEN 2PK MOUSE TRAPS|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00029049006026|BROOMS/MOPS & BRUSHES|GM|-80.497332|1.4049434824709919|178|2
35.667941|79fa696820df0f5f39e38e8854611ad4685c4164|0.84|2014-09-17 19:30:00|1.4057311447477159|2||178|0.6225230078570788|0|52|502|-80.497332|64|35.667941|FRESH BANANAS|0.0|4|BANANAS, YELLOW|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00204011000008|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|bbe63a766368cec0a77d9d9dcd53f2f8fdad5b91|4.99|2015-02-18 16:05:00|1.4057311447477159|2|7203695597|178|0.6225230078570788|0|52|1603|-80.497332|371|35.667941|PRIVATE LABEL BREAD|1.0|14|BAND OF BAKERS MERLOT BOULE|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00072036955975|BREAD|BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|a70fc192e118a6a33ff01c94df43ccd0be9a9a0b|3.29|2014-11-11 10:27:00|1.4057311447477159|2|7203698555|178|0.6225230078570788|0|52|427|-80.497332|72|35.667941|NFS-TOILET TISSUE|0.5|1|HT 1000 SHEET BATHTISSUE 4 RL|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00072036985552|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|683a7fb0b488bcafb588de5b7e3b06634c6ed15a|1.1|2014-09-11 17:02:00|1.4057311447477159|2||178|0.6225230078570788|0|52|526|-80.497332|64|35.667941|FRESH MUSHROOMS|0.0|4|USA WHITE MUSHROOMS, BULK|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00204085000003|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|a92d724855680d65689ec31465431970bc334823|0.54|2015-03-03 14:40:00|1.4057311447477159|2|7203641210|178|0.6225230078570788|0|52|257|-80.497332|39|35.667941|TOMATOES|0.0|1|HT TOMATO SAUCE 8|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00072036412102|VEGETABLES-CAN/JAR|G1 GROCERY|-80.497332|1.4049434824709919|178|2
35.667941|d7c35430871dbba5bdc9614d768cf6fe0f118342|18.99|2015-02-03 17:48:00|1.4057311447477159|2|20220200000|178|0.6225230078570788|0|52|299|-80.497332|49|35.667941|ANGUS BEEF|4.75|2|ANGUS BEEF FILET MIGNON|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00202204000002|BEEF|MEAT|-80.497332|1.4049434824709919|178|1
35.667941|fbf9cba1d1ea0a70bb0fe4e95483945826fbd80b|3.99|2014-11-19 21:34:00|1.4057311447477159|2|71514151464|178|0.6225230078570788|0|52|364|-80.497332|55|35.667941|ORGANIC AND CF EGGS|0.0|3|EGGLAND'S BEST CAGE FREE LARGE|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00715141514643|EGGS FRESH|DAIRY|-80.497332|1.4049434824709919|178|1
35.667941|5899d346e155062f63008dd3d24b4d9ac000d3ef|2.0|2014-11-07 15:58:00|1.4057311447477159|2||178|0.6225230078570788|0|52|512|-80.497332|64|35.667941|FRSH PROD FRSH FRUIT REM|0.0|4|MANGOS|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00204959000009|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|2
35.667941|94b54279ac0e492faa8030225e37a0ab1e703e83|1.79|2014-11-05 21:26:00|1.4057311447477159|2|7203663157|178|0.6225230078570788|0|52|1134|-80.497332|57|35.667941|CARTON MILK|0.0|3|HARRIS TEETER WHOLE MILK|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00072036631572|MILK|DAIRY|-80.497332|1.4049434824709919|178|1
35.667941|1d595f72d6d6b7913b2e7c8d4bbbe0a05041ef6e|6.99|2014-11-01 12:11:00|1.4057311447477159|2|73150956699|178|0.6225230078570788|0|52|3087|-80.497332|1000|35.667941|FALSE NAIL KIT-OTHER MANUF|0.0|17|KISS NAIL DRESS STRIP PUSHUP|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00731509567458|COSMETICS|HBC|-80.497332|1.4049434824709919|178|1
35.667941|6c5e1e39f91033cfb5bc7b79213a98c9ebf3b51d|5.69|2014-10-01 18:25:00|1.4057311447477159|2|4720015264|178|0.6225230078570788|0|52|312|-80.497332|51|35.667941|BUTTER|1.7|3|CHALLENGE UNSALTED BUTTER|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00047200152665|BUTTER & MARGARINE|DAIRY|-80.497332|1.4049434824709919|178|1
35.667941|cc19d917feed1f5c14f822be7d0fcac5b9381eab|4.59|2014-11-25 10:29:00|1.4057311447477159|2|78142100128|178|0.6225230078570788|0|52|1601|-80.497332|371|35.667941|BRANDED BREAD|0.0|14|LA BREA SOURDOUGH LOAF|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00781421001288|BREAD|BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|92d19302def3b74eb17aed7b6f9394f450b6eba6|4.59|2015-02-15 18:58:00|1.4057311447477159|2|78142100128|178|0.6225230078570788|0|52|1601|-80.497332|371|35.667941|BRANDED BREAD|0.0|14|LA BREA SOURDOUGH LOAF|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00781421001288|BREAD|BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|e71cd2ce5ef8cc5a17fc02b5fa9654f6b1b5c640|2.36|2014-09-13 13:58:00|1.4057311447477159|2||178|0.6225230078570788|0|52|522|-80.497332|64|35.667941|FRESH TOMATOES|0.0|4|RED H/H TOMATOES, BULK|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00204799000009|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|14a5bc538de2b26f242dc06b056cbc27cd17df29|3.47|2015-02-11 17:31:00|1.4057311447477159|2|7203659020|178|0.6225230078570788|0|52|312|-80.497332|51|35.667941|BUTTER|0.97|3|HARRIS TEETER BUTTER QUARTERS|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00072036590206|BUTTER & MARGARINE|DAIRY|-80.497332|1.4049434824709919|178|1
35.667941|fc95ea5fa0738dd715e49e739cd0d295708c3b3a|3.99|2014-09-30 14:30:00|1.4057311447477159|2|7203670719|178|0.6225230078570788|0|52|427|-80.497332|72|35.667941|NFS-TOILET TISSUE|0.0|1|YH BATH ULTRA STRONG 12DR|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00072036707192|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|6c6e96d577c5e0443384cecacadb326ceff44bf7|2.85|2014-12-23 16:06:00|80.497482303704658|2|7433610005|178|35.708501930169568|0|6|342|-80.66939|57|35.28326|FRESH MILK|0.0|3|HUNTER  WHOLE MILK|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|35.699188602026126|00074336100055|MILK|DAIRY|-80.497332|80.497571076724597|46|1
35.667941|9e67ba13a9ae93f0053edc3dfceeef208bde1c63|2.91|2014-10-17 20:41:00|1.4057311447477159|2|7203698757|178|0.6225230078570788|0|52|31|-80.497332|4|35.667941|NON CARBONATED WATER|0.0|1|HT PURIFIED WATER|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00072036987570|BOTTLED WATER|G1 GROCERY|-80.497332|1.4049434824709919|178|3
35.667941|65d32d57b67a03d7d85526f912221fc31697ad33|11.99|2014-11-01 15:32:00|1.4057311447477159|2|78535710062|178|0.6225230078570788|0|52|35|-80.497332|10|35.667941|PREMIUM WHOLE BEAN|4.0|1|PEET'S MAJOR DICKASON WB|9bc681da62f2e6d63421eb633bc66c99eab74b6d|2.802694439965691|0.6209993146566879|00785357100626|COFFEE|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.297134|11cb39857d1b1d12c6d2aec11c7eedc0617a238c|2.55|2014-11-09 13:48:00|80.728244613218536|3|4119601012|258|35.301281038748797|0|5|1201|-80.825175|33|35.152722|RTS CANNED|0.55|1|PROG VEG CLASSIC LENTIL|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|35.296297200616316|00041196010220|SOUP|G1 GROCERY|-80.737839|80.73784864545155|160|1
35.297134|b876bf78135e9350d34dbc7179c0dc02723f4978|12.99|2014-11-22 17:04:00|80.728244613218536|3|8254400904|258|35.301281041339649|0|5|9954|-80.80146|886|35.17739|NFS-PREM-ZINFANDEL|0.0|13|OAK RIDGE ZIN OLD VINES|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|35.296297200616316|00082544009046|PREMIUM ($8-$10.99)|WINE|-80.737839|80.737846795751622|208|1
35.297134|c765aab3e720f4569cf39f6de57a3bcedfac8b7c|5.49|2015-02-14 15:17:00|80.728244613218536|3|4900000548|258|35.301281035316919|0|5|54|-80.806073|8|35.106477|DIET|0.5|23|DTDR PEPPER 12OZ PET8PK BOTTLE|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|35.296297200616316|00078000083316|CARBONATED BEVERAGES|BEVERAGE|-80.737839|80.737850651939581|4|1
35.297134|4d83bb41e31942269c7b942729910ac64caa371a|44.69|2014-11-07 14:13:00|80.728244613218536|3|20221900000|258|35.301281039720365|0|5|299|-80.85013|49|35.175855|ANGUS BEEF|17.2|2|ANGUS STEAKHOUSE STRIP ROAST|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|35.296297200616316|00202105000002|BEEF|MEAT|-80.737839|80.737847996491638|218|1
35.297134|1e25398b14affc502b5cd7f180861f7550889b77|3.99|2014-10-12 14:33:00|80.728244613218536|3|20405400000|258|35.301281038748797|0|5|504|-80.825175|64|35.152722|FRESH BERRIES|0.2|4|RED RASPBERRIES 6 OZ|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|35.296297200616316|00812049004402|FRESH PRODUCE|PRODUCE|-80.737839|80.73784864545155|160|1
35.297134|f64d73b9a500d44e20f3607cc4bdd9b7659dba8c|8.99|2014-10-02 18:58:00|80.728244613218536|3|8130859187|258|35.301281039720365|0|5|9948|-80.85013|886|35.175855|NFS-PREM-CAB SAUVIGNON|0.0|13|CUPCAKE CAB SAUV|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|35.296297200616316|00081308591872|PREMIUM ($8-$10.99)|WINE|-80.737839|80.737847996491638|218|1
35.297134|f3025ae1c47446ad1a9bfb84e80f1783bc5753ed|1.59|2014-11-01 14:20:00|80.728244613218536|3|7152415913|258|35.301281038748797|0|5|1214|-80.825175|272|35.152722|AUTHENTIC HISPANIC|0.0|1|LA PREF ORG DICED GRN CHILIES.|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|35.296297200616316|00071524159130|HISPANIC PREP. FOODS|G1 GROCERY|-80.737839|80.73784864545155|160|1
35.297134|893d419e5ed69ea83fef7087af8f8e1cbcff85e7|9.29|2014-12-24 14:20:00|80.728244613218536|3|20606300000|258|35.301281041339649|0|5|2018|-80.80146|505|35.17739|PRESSED CHEESE|0.0|6|AFON CLEDDAU  CHEDDR (FC)|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|35.296297200616316|00206063000005|SPECIALTY CHEESE|DELI|-80.737839|80.737846795751622|208|1
35.297134|4ac63bfffd72e5cc94b6d6baa07e54a0bc3879c4|4.99|2014-11-02 12:15:00|80.728244613218536|3|78142100529|258|35.301281038748797|0|5|1601|-80.825175|371|35.152722|BRANDED BREAD|0.0|14|LA BREA SEEDED RYE BREAD|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|35.296297200616316|00781421005293|BREAD|BAKERY|-80.737839|80.73784864545155|160|1
35.297134|579ed2c6acca9d76026e4ca2a37893b5f613161b|2.78|2014-12-23 15:27:00|80.728244613218536|3|5210094269|258|35.301281038748797|0|5|80|-80.825175|34|35.152722|SEASONING PACKETS|0.78|1|E  MC CHILI SEASONING MIX|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|35.296297200616316|00052100091501|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.737839|80.73784864545155|160|2
35.297134|dd54f654eafc27a419199b68244ac76f24352490|13.99|2014-10-25 19:50:00|80.728244613218536|3|8600300165|258|35.30128104436286|0|5|9938|-80.661096|885|35.172688|NFS POP PINOT GRS/GRIGIO|0.0|13|WOODBRIDGE PINOT GRIGIO 1.5L|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|35.296297200616316|00086003001657|POPULAR (4-$7.99)|WINE|-80.737839|80.737843809288606|474|1
35.297134|78d960d980858d0f3b82e634d4d4449a77b0c293|9.99|2015-03-01 13:18:00|80.728244613218536|3|8500001222|258|35.301281041339649|0|5|9939|-80.80146|885|35.17739|NFS POP PINOT NOIR|0.0|13|REDWOOD CREEK PINOT NOIR 1.5L|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|35.296297200616316|00085000012222|POPULAR (4-$7.99)|WINE|-80.737839|80.737846795751622|208|1
35.297134|4b2f4467f73bce2379205dee2ad0d2e0825024bc|7.99|2015-03-08 14:32:00|80.728244613218536|3|7203676196|258|35.301281041339649|0|5|35|-80.80146|10|35.17739|PREMIUM WHOLE BEAN|2.42|1|HT TRADER COFFEE WB BRFST BLEN|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|35.296297200616316|00072036761965|COFFEE|G1 GROCERY|-80.737839|80.737846795751622|208|1
35.297134|ce67706aae8835510164e7b02330a618eac31447|0.79|2014-12-06 14:17:00|80.728244613218536|3|7203688001|258|35.301281038748797|0|5|527|-80.825175|64|35.152722|FRESH CARROTS|0.0|4|HT WHOLE CARROTS 1LB BAG|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|35.296297200616316|00072036880017|FRESH PRODUCE|PRODUCE|-80.737839|80.73784864545155|160|1
35.297134|9aa322a831995b59ed710c92d8518273758b2925|5.97|2014-10-11 17:06:00|80.728244613218536|3|7203676359|258|35.301281038748797|0|5|345|-80.825175|57|35.152722|ORGANIC MILK|0.0|3|HTO ORGANIC 2% MILK GAL|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|35.296297200616316|00072036763600|MILK|DAIRY|-80.737839|80.73784864545155|160|1
35.297134|e4f6da379d701b5ffcfca1242d009ac5ed9d9bed|1.19|2014-10-11 17:07:00|80.728244613218536|3|2620011700|258|35.301281038748797|0|5|206|-80.825175|31|35.152722|FRONT END SNACKS|0.0|1|SLIM JIM ORIGINAL GIANT|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|35.296297200616316|00026200117003|SNACKS|G1 GROCERY|-80.737839|80.73784864545155|160|1
35.297134|e650f3b276114307197ab55dc8c39087ed5ab387|4.99|2014-11-12 10:53:00|80.728244613218536|3|7203688137|258|35.301281039720365|0|5|500|-80.85013|64|35.175855|FRESH APPLES|0.0|4|HT BRAEBURN APPLE 3LB|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|35.296297200616316|00072036881373|FRESH PRODUCE|PRODUCE|-80.737839|80.737847996491638|218|1
35.297134|d7f946596f49567e2fce9d45c2be04b922e46fbc|1.77|2014-09-17 08:55:00|80.728244613218536|3|7009030410|258|35.301281041339649|0|5|225|-80.80146|35|35.17739|SUGAR-GRANULATED|0.0|1|CRYSTAL FINE GRANULATED SUGAR|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|35.296297200616316|00070090304104|SUGAR/SUBSTITUTES|G1 GROCERY|-80.737839|80.737846795751622|208|1
35.297134|b51af3270c1444e096413141a405b65ffac6092a|4.47|2014-09-20 14:30:00|80.728244613218536|3|519|258|35.301281038748797|0|5|1896|-80.825175|450|35.152722|SODA|0.0|6|24 OZ FOUNTAIN DRINK|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|35.296297200616316|00000000005190|BEVERAGES|DELI|-80.737839|80.73784864545155|160|3
35.297134|d1a0cce3b6d06dbf03cac766cf02632e5bd9f3b0|1.99|2014-11-09 13:22:00|80.728244613218536|3|78616200387|258|35.301281038748797|0|5|31|-80.825175|4|35.152722|NON CARBONATED WATER|1.0|1|FRUITWATER TROPICAL PINEAPPLE|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|35.296297200616316|00786162004444|BOTTLED WATER|G1 GROCERY|-80.737839|80.73784864545155|160|1
35.297134|b47d2cec64f571626d8cf4f9d8f519ccff5a0629|3.59|2014-10-11 12:28:00|80.728244613218536|3|7225003706|258|35.301281039720365|0|5|1026|-80.85013|162|35.175855|WHEAT|1.3|7|NATOWN HONEYWHEAT BRD|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|35.296297200616316|00072250037068|SLICED BREAD|COMMERCIAL BAKERY|-80.737839|80.737847996491638|218|1
35.297134|31b0615a48ee4cc706af8a5f28743a891ccaefb6|0.5|2014-09-10 15:28:00|1.4094857484078087|3|2840004176|258|0.6160512048176361|0|26|206|-80.737839|31|35.297134|FRONT END SNACKS|0.0|1|MUNCHIES SALTED PEANUTS|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|0.61471665291522548|00028400041768|SNACKS|G1 GROCERY|-80.737839|1.409141121495086|258|1
35.297134|45bc72cb73062da2aa584d9e4e991e8ba1ffcb89|7.99|2014-10-20 17:40:00|80.728244613218536|3|2210000288|258|35.301281035528916|0|5|454|-80.824767|82|35.116751|DOMESTIC ECONOMY 12PK&>|0.0|16|PABST 12PK 12OZ BTL|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|35.296297200616316|00022100002883|DOMESTIC BEER|BEER|-80.737839|80.737850538111246|294|1
35.297134|0427ed31f0a986b61b8e58946bab6de714570e57|16.82|2014-11-19 12:49:00|80.728244613218536|3|20812800000|258|35.301281039720365|0|5|664|-80.85013|145|35.175855|SHRIMP WILD CAUGHT|4.95|12|FRESH WILD CAUGHT 21/30 CT EAS|9cb3f9c671cd8bea0b6578f548b5afd83e88016c|0.2865508790685545|35.296297200616316|00208128000005|SHRIMP|SEAFOOD|-80.737839|80.737847996491638|218|1
35.17739|299c847fefd0212a173622d2376c02af06635027|5.29|2014-12-12 15:33:00|80.810069425230125|4|7203603031|208|35.236388386441149|0|23|4296|-80.810056|1205|35.219587|ACETAMINOPHEN|1.3|17|HT ACETAMINOPHEN CAPS 50CT|9de0a8e5c6b661ab1fc24b3e8a35c17c9655bd03|4.076646353405749|35.240679762029046|00072036030313|PAIN RELIEF|HBC|-80.80146|80.801488891276477|401|1
35.667941|8ed548999ae0b004042a9187a0462978f2bebd30|2.69|2014-12-01 15:20:00|80.497482303704658|1|70935100013|178|35.69150730682852|0|6|556|-80.860108|64|35.500972|PACKAGED VEGETABLES|0.0|4|APIO BROCCOLI & CAULIFLOWER|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00709351000263|FRESH PRODUCE|PRODUCE|-80.497332|80.497430447440678|268|1
35.667941|5b0485c7c22173e36827b88a0ce0dc79aa4a9348|4.99|2014-11-25 16:42:00|80.497482303704658|1|61300872592|178|35.69150730682852|0|6|99|-80.860108|32|35.500972|LIQUID TEA|0.0|1|ARNOLD PALMER LT HALF/HALF 12P|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00613008725921|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.497332|80.497430447440678|268|1
35.667941|e773f2b250da984d14e6c11e10f707d960a731c7|11.95|2015-02-02 18:42:00|80.497482303704658|1|76211101266|178|35.69150730682852|0|6|1583|-80.860108|370|35.500972|VIA|0.0|22|KCUP GUAT. ANT. BLEND 12 CT|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00762111012661|STARBUCKS|COFFEE SHOP|-80.497332|80.497430447440678|268|1
35.667941|d79973aeaadfc2752147e958c062ac1c2d8b999f|2.69|2014-12-11 09:56:00|80.497482303704658|1|70935100013|178|35.69150730682852|0|6|556|-80.860108|64|35.500972|PACKAGED VEGETABLES|0.0|4|APIO BROCCOLI & CAULIFLOWER|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00709351000263|FRESH PRODUCE|PRODUCE|-80.497332|80.497430447440678|268|1
35.667941|d480d09d8ffc89904c5c51dd287d1077330cee30|3.99|2015-02-12 11:24:00|1.4057311447477159|1|20405400000|178|0.6225230078570788|0|52|504|-80.497332|64|35.667941|FRESH BERRIES|0.0|4|RED RASPBERRIES 6 OZ|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00761635201605|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|934a95750af0048a1a3bb87ada2e129f280c2459|3.99|2015-02-20 12:44:00|1.4057311447477159|1|20405400000|178|0.6225230078570788|0|52|504|-80.497332|64|35.667941|FRESH BERRIES|0.0|4|RED RASPBERRIES 6 OZ|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00761635201605|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|4c8fb598efb0bdcba6b3e88528d75a74e95104a9|3.99|2015-02-01 14:42:00|1.4057311447477159|1|20405400000|178|0.6225230078570788|0|52|504|-80.497332|64|35.667941|FRESH BERRIES|0.0|4|RED RASPBERRIES 6 OZ|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00761635201605|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|8e7aaf92ac380432571f72c0b45f1a519b31268a|4.99|2015-01-01 14:13:00|80.497482303704658|1|61300872592|178|35.69150730682852|0|6|99|-80.860108|32|35.500972|LIQUID TEA|0.0|1|ARNOLD PALMER LT HALF/HALF 12P|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00613008725921|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.497332|80.497430447440678|268|1
35.667941|38d567584c1be5e2c07ca60b38aa3ca1cd748de2|3.66|2014-09-15 09:43:00|1.4057311447477159|1||178|0.6225230078570788|0|52|505|-80.497332|64|35.667941|FRESH SOFT FRUIT|2.21|4|EASTERN PEACHES|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00204403000005|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|11648b8b92d559bdac132132bd2489c44cad9722|2.29|2014-11-24 18:46:00|80.497482303704658|1||178|35.69150730682852|0|6|540|-80.860108|64|35.500972|FRESH CELERY|0.0|4|CELERY HEARTS (RPC)|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00204575000001|FRESH PRODUCE|PRODUCE|-80.497332|80.497430447440678|268|1
35.667941|a64b0c5432b015ce6d08814c84f2d9ebff7969a9|11.99|2014-11-20 14:35:00|1.4057311447477159|1|4300004648|178|0.6225230078570788|0|52|66|-80.497332|10|35.667941|GROUND CAN|6.0|1|MAXWELL HOUSE MASTER BLEND|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00043000046500|COFFEE|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|5a47369ce1bbc053e4d7cd21559cd0d8707ca299|6.58|2014-12-13 13:27:00|80.497482303704658|1|4300027678|178|35.69150730682852|0|6|20|-80.860108|3|35.500972|COCONUT|1.0|1|BAKERS COCONUT BAG|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00043000276785|BAKING SUPPLIES|G1 GROCERY|-80.497332|80.497430447440678|268|2
35.667941|d7f744120836bff67be3e8878b117518240873f0|2.99|2015-01-28 14:34:00|80.497482303704658|1|4119689107|178|35.691507255430857|0|6|120|-80.861571|15|35.444615|COATINGS & BREADERS|0.0|1|PROGRESSO BREAD CRUMBS ITALIAN|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00041196891072|FLOUR|G1 GROCERY|-80.497332|80.497447600120879|340|1
35.667941|9b96b0e5cda4a6287bd4dcba1bc8694572826856|3.0|2014-11-27 10:28:00|80.497482303704658|1|4023217761|178|35.691507293415832|0|6|8598|-80.762919|1792|35.442529|NEWSPAPERS|0.0|18|CHARLOTTE OBSERVER THANKGIVING|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00040232177613|NEWSPAPERS|GM|-80.497332|80.49743519887393|471|1
35.667941|ffda29b33cbf61264a1528aed68dd50e6b16fa13|8.97|2014-11-08 13:22:00|80.497482303704658|1|4150080502|178|35.69150730682852|0|6|76|-80.860108|11|35.500972|MEAT SAUCES|0.0|1|FRANKS RED HOT 12 SAUCE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00041500805023|CONDIMENTS|G1 GROCERY|-80.497332|80.497430447440678|268|3
35.667941|5d333ca0034c337d6ca5a698f9516826db9c133b|10.65|2015-01-13 13:35:00|80.497482303704658|1|4173601013|178|35.69150730682852|0|6|194|-80.860108|30|35.500972|OLIVE OIL|3.66|1|FILIPPO BERIO EX VIRGIN OLIVE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00041736010130|SHORTENING/OIL|G1 GROCERY|-80.497332|80.497430447440678|268|1
35.667941|a4b9f27fca81798442d70046b13bae160f4210f9|2.99|2014-11-20 15:26:00|80.497482303704658|1|4119689107|178|35.69150730682852|0|6|120|-80.860108|15|35.500972|COATINGS & BREADERS|0.0|1|PROGRESSO BREAD CRUMBS ITALIAN|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00041196891072|FLOUR|G1 GROCERY|-80.497332|80.497430447440678|268|1
35.667941|c8e60da2e928b9c339f1aa6b5380199ae1e5d9e0|1.69|2014-10-23 17:45:00|80.497482303704658|1|7680828073|178|35.69150730682852|0|6|149|-80.860108|23|35.500972|WHSE PASTA CORE|0.0|1|BARILLA PASTA PENNE RIGATE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00076808280739|PASTA|G1 GROCERY|-80.497332|80.497430447440678|268|1
35.667941|4e7c1bc2779bf4764950702da3ebcd4a357ed767|6.58|2015-02-24 12:11:00|1.4057311447477159|1|7265546007|178|0.6225230078570788|0|52|1278|-80.497332|48|35.667941|SINGLE SERVE NUTRITIONAL|0.0|5|HC FOUR CHS ZITI BAKE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00072655460010|FROZEN MEALS|FROZEN|-80.497332|1.4049434824709919|178|2
35.667941|c75588f489944c70b5bafa29c123a138213176b4|6.3|2014-09-26 16:21:00|1.4057311447477159|1|7265500105|178|0.6225230078570788|0|52|1278|-80.497332|48|35.667941|SINGLE SERVE NUTRITIONAL|1.15|5|HC CAFE STEAMERS BASIL CHICKEN|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00072655001145|FROZEN MEALS|FROZEN|-80.497332|1.4049434824709919|178|2
35.667941|76783661bb5ff3f800138e25b56faac5c1576c2e|2.99|2014-09-28 16:02:00|1.4057311447477159|1|7080004879|178|0.6225230078570788|0|52|978|-80.497332|202|35.667941|SMOKED MEATS|0.0|2|SMITHFIELD BONELESS HAM STEAK|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00070800048793|SMOKED HAMS|MEAT|-80.497332|1.4049434824709919|178|1
35.667941|ca57b46dbf6e4647929910b63518882920a681cd|3.99|2014-12-15 18:58:00|80.497482303704658|1|5150000163|178|35.69150730682852|0|6|123|-80.860108|19|35.500972|JELLY/JAMS|0.0|1|SMUCKER STRAWBERRY JAM|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00051500001639|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.497332|80.497430447440678|268|1
35.667941|23e363af6e01e7bd31adaca21ac687954fa3a97d|3.79|2014-09-14 12:52:00|1.4057311447477159|1|5160000001|178|0.6225230078570788|0|52|76|-80.497332|11|35.667941|MEAT SAUCES|0.0|1|LEA & PERRINS WORCESTERSHIRE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00051600000013|CONDIMENTS|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|3967e97c9eeb9ffce8e12862b3de9ecdfe6df363|4.59|2014-11-01 12:02:00|1.4057311447477159|1|5450019322|178|0.6225230078570788|0|52|484|-80.497332|101|35.667941|BEEF WIENERS|2.3|19|BALL PARK BEEF FRANKS|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00054500193229|WIENERS|CASE READY MEATS|-80.497332|1.4049434824709919|178|1
35.667941|1c2179d651790534e6a40d591565b5fc803a19ab|4.0|2014-09-13 17:51:00|80.497482303704658|1|7962501164|178|35.691507255430857|0|6|4171|-80.861571|1085|35.444615|TRAVEL SET|0.0|17|(JHK) 4PC 3OZ TRAVL BOTTLE SET|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00079625011647|TRIAL SIZE|HBC|-80.497332|80.497447600120879|340|1
35.667941|74e29abd790c77cfb1a6a2e2dcad26c629435ee7|8.22|2015-02-15 13:58:00|80.497482303704658|1|20165500000|178|35.691507293415832|0|6|297|-80.762919|49|35.442529|GROUND BEEF|0.0|2|HT PREMIUM GRND BEEF 80% LEAN|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00201655000005|BEEF|MEAT|-80.497332|80.49743519887393|471|2
35.667941|1faec844cf3fbaf76d2ebece84a4927344437e90|6.42|2014-12-22 15:30:00|80.497482303704658|1|20165500000|178|35.69150730682852|0|6|297|-80.860108|49|35.500972|GROUND BEEF|0.0|2|HT PREMIUM GRND BEEF 80% LEAN|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00201655000005|BEEF|MEAT|-80.497332|80.497430447440678|268|1
35.667941|d1c6a540701241a25c8177beef30a3fa3ff993f6|7.9|2014-10-23 16:04:00|80.497482303704658|1|20165500000|178|35.69150730682852|0|6|297|-80.860108|49|35.500972|GROUND BEEF|0.59|2|HT PREMIUM GRND BEEF 80% LEAN|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00201655000005|BEEF|MEAT|-80.497332|80.497430447440678|268|1
35.667941|2dfcb16b25770409840b07cf6657061910c7a3f1|4.29|2014-09-24 14:30:00|80.497482303704658|1|7797508217|178|35.69150730682852|0|6|202|-80.860108|31|35.500972|PRETZELS|0.3|1|SOH 100 CAL STICKS PRETZ LUNCH|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00077975082171|SNACKS|G1 GROCERY|-80.497332|80.497430447440678|268|1
35.667941|6713db1184e734978da44c7b65876ec333aae5c0|4.75|2015-02-04 13:13:00|80.497482303704658|1|20165500000|178|35.69150730682852|0|6|297|-80.860108|49|35.500972|GROUND BEEF|0.36|2|HT PREMIUM GRND BEEF 80% LEAN|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00201655000005|BEEF|MEAT|-80.497332|80.497430447440678|268|1
35.667941|88b12198639dc4001ed742f7f48f85a0f3de4c49|5.91|2014-10-01 12:25:00|80.497482303704658|1|20165500000|178|35.69150730682852|0|6|297|-80.860108|49|35.500972|GROUND BEEF|0.0|2|HT PREMIUM GRND BEEF 80% LEAN|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00201655000005|BEEF|MEAT|-80.497332|80.497430447440678|268|1
35.667941|69c7f6788ade4fcf0143eaba247e5094d68ce206|3.69|2015-01-22 14:36:00|80.497482303704658|1|7797508822|178|35.69150730682852|0|6|202|-80.860108|31|35.500972|PRETZELS|0.69|1|SOH CHEDDAR  PIECES|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00077975088210|SNACKS|G1 GROCERY|-80.497332|80.497430447440678|268|1
35.667941|f2d290f232f8273a8dee6063e5bee17c7a318ce9|6.98|2014-10-12 12:06:00|1.4057311447477159|1|3000001190|178|0.6225230078570788|0|52|60|-80.497332|9|35.667941|HOT CEREAL|1.98|1|QUAKER OATML REGULAR|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00030000012109|CEREAL|G1 GROCERY|-80.497332|1.4049434824709919|178|2
35.667941|1e59169e4d82a7301cadc1a473d0879949effea1|9.45|2014-12-03 11:55:00|1.4057311447477159|1|3000001190|178|0.6225230078570788|0|52|60|-80.497332|9|35.667941|HOT CEREAL|1.9500000000000002|1|QUAKER OATML REGULAR|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00030000012109|CEREAL|G1 GROCERY|-80.497332|1.4049434824709919|178|3
35.667941|fb7d9cf9a83c412e2050ce9fdf35893603536832|1.79|2015-01-13 15:11:00|1.4057311447477159|1|2120001023|178|0.6225230078570788|0|52|6648|-80.497332|1564|35.667941|HOME/OFFICE TAPE|0.0|18|SCOTCH MAGIC TAPE-01023|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00021200010231|SCHOOL & OFFICE SUPPLY|GM|-80.497332|1.4049434824709919|178|1
35.667941|1d2ca5d308c406b55a4760ab3ec5dbe3db350e7a|2.89|2014-12-23 17:56:00|80.497482303704658|1|2100065894|178|35.69150730682852|0|6|1441|-80.860108|274|35.500972|MAC AND CHEESE|0.0|1|KRAFT DIN MAC CHS FAMILY|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00021000658947|PREP FOODS DINNERS|G1 GROCERY|-80.497332|80.497430447440678|268|1
35.667941|a6d4d0737ad8801db28f5e8e7546973a17172e0b|5.7|2014-11-21 15:13:00|80.497482303704658|1|1800000401|178|35.69150730682852|0|6|327|-80.860108|54|35.500972|DINNER ROLLS-REFRIGERATED|1.7|3|PILLSBURY CRESCENT ROLLS|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00018000004010|DOUGH PRODUCTS|DAIRY|-80.497332|80.497430447440678|268|2
35.667941|1651434953f5902fa7fbd4c63063bfa2c3540def|1.69|2014-09-29 14:36:00|80.497482303704658|1|7680828073|178|35.69150730682852|0|6|149|-80.860108|23|35.500972|WHSE PASTA CORE|0.31|1|BARILLA PASTA RIGATONI|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00076808502947|PASTA|G1 GROCERY|-80.497332|80.497430447440678|268|1
35.667941|d35cce87fe73ee99cf7a0207a82aba5a325b3d9d|4.99|2014-10-30 12:06:00|1.4057311447477159|1|1111018700|178|0.6225230078570788|0|52|1647|-80.497332|379|35.667941|PACKAGED MUFFINS|2.5|14|FFM 4 CT CRAN ORANGE MUFFIN|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00011110187062|MUFFINS|BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|0502da36c2163cf2ff611bee6b5d0b22301a8d58|4.99|2014-10-24 11:42:00|1.4057311447477159|1|1111018700|178|0.6225230078570788|0|52|1647|-80.497332|379|35.667941|PACKAGED MUFFINS|1.02|14|FFM 4 CT CRAN ORANGE MUFFIN|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00011110187062|MUFFINS|BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|46e586b6dd3ac56fb03f92f513dc4ae4e2bc9d6f|4.99|2014-10-17 11:25:00|1.4057311447477159|1|1111018700|178|0.6225230078570788|0|52|1647|-80.497332|379|35.667941|PACKAGED MUFFINS|1.02|14|FFM 4 CT CRAN ORANGE MUFFIN|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00011110187062|MUFFINS|BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|151998c38adee3c2dfc17f38bf967aab4d110bd9|3.29|2014-11-26 15:40:00|80.497482303704658|1|1204403891|178|35.69150730682852|0|6|3816|-80.860108|1070|35.500972|INVISIBLE-MALE|0.0|17|OLD SPICE HE INV SOL PURE SPRT|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00012044000250|DEODORANT|HBC|-80.497332|80.497430447440678|268|1
35.667941|c70cfad65a727d3cf1a28f6321727c5a3b785c27|3.78|2014-10-02 13:54:00|80.497482303704658|1|1600027488|178|35.691507255430857|0|6|165|-80.861571|26|35.444615|DEHYDRATED POTATOES|0.0|1|BC POTATOES SCALLOPED CHEESE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00016000406704|PREPARED FOODS-DRY MIXES|G1 GROCERY|-80.497332|80.497447600120879|340|2
35.667941|fc7849f2cda0871aad086bff2e19c739d157a5e6|2.69|2014-12-22 11:01:00|1.4057311447477159|1|1480000179|178|0.6225230078570788|0|52|124|-80.497332|16|35.667941|APPLESAUCE MULTISERVE|0.0|1|MOTTS APPLESAUCE 23 ORIGINAL.|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00014800001792|FRUIT-CAN/JAR|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|654b9d273a358b3a6db9b253f76052308d838cff|19.99|2014-10-25 14:52:00|80.497482303704658|1|7203695592|178|35.691507293415832|0|6|1653|-80.762919|381|35.442529|CELEBRATION CAKES|0.0|14|1/4 SHT DL MARBLE CAK  W/BUTCR|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00072036955920|CAKES|BAKERY|-80.497332|80.49743519887393|471|1
35.667941|81de06d88626ada2e0bc47bd955a3db54dc580d1|3.99|2015-03-02 10:38:00|1.4057311447477159|1|7203695283|178|0.6225230078570788|0|52|1663|-80.497332|381|35.667941|CREME CAKE|0.0|14|FFM SLICED LEMON CAKE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00072036952950|CAKES|BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|59627070336cfdea4224f1268e91106c17589dcb|3.99|2014-11-25 10:43:00|1.4057311447477159|1|7203695283|178|0.6225230078570788|0|52|1663|-80.497332|381|35.667941|CREME CAKE|0.0|14|FFM SLICED POUND CAKE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00072036952752|CAKES|BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|5ea99de7d7b81b2fee0e6b9488c63b1312ee1178|12.99|2014-09-27 18:00:00|80.497482303704658|1|7203695587|178|35.69150730682852|0|6|1707|-80.860108|387|35.500972|MESSAGE|3.0|14|12 INCH MESSAGE COOKIE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00072036955876|COOKIES|BAKERY|-80.497332|80.497430447440678|268|1
35.667941|7ce6bcd50f21511e80c99d1fa25c7d2bc160f20e|3.99|2015-02-14 13:39:00|1.4057311447477159|1|7203695283|178|0.6225230078570788|0|52|1663|-80.497332|381|35.667941|CREME CAKE|1.0|14|FFM SLICED LEMON CAKE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00072036952950|CAKES|BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|64a244227093ad7376b52cce2d767e6b2ee5a5e0|3.99|2015-03-08 12:13:00|1.4057311447477159|1|7203695283|178|0.6225230078570788|0|52|1663|-80.497332|381|35.667941|CREME CAKE|0.0|14|FFM SLICED LEMON CAKE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00072036952950|CAKES|BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|627af745ed29d8b06798cbf2415cda1c38ae28ee|3.99|2015-01-24 11:56:00|1.4057311447477159|1|7203695283|178|0.6225230078570788|0|52|1663|-80.497332|381|35.667941|CREME CAKE|0.0|14|FFM SLICED LEMON CAKE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00072036952950|CAKES|BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|7558e3fc2ed83f0465cf29f24c19c600cbba90fd|4.39|2014-09-21 12:37:00|1.4057311447477159|1|1920083721|178|0.6225230078570788|0|52|404|-80.497332|69|35.667941|NFS-TOILET BOWL CLEANERS|0.0|1|LYSOL TOILET BWL CLNR LIME|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00019200882095|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|99a25c16250ccd72b85fc2efb3bebe61f719856b|3.99|2015-01-23 10:18:00|1.4057311447477159|1|1630016564|178|0.6225230078570788|0|52|335|-80.497332|56|35.667941|ORANGE JUICE-REGRIGERATED|0.0|3|FL NAT NO PULP W/CALCIUM OJ|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00016300165677|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.497332|1.4049434824709919|178|1
35.667941|8d7c5b0d4da63da423437cd61ebc9dbb2c8d2b1a|3.99|2014-12-27 13:50:00|1.4057311447477159|1|1630016564|178|0.6225230078570788|0|52|335|-80.497332|56|35.667941|ORANGE JUICE-REGRIGERATED|0.0|3|FL NAT NO PULP W/CALCIUM OJ|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00016300165677|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.497332|1.4049434824709919|178|1
35.667941|98dd6ded2d899eeb92b6bfc383b6b46ac1a89c87|2.99|2014-12-20 10:49:00|1.4057311447477159|1|81204900640|178|0.6225230078570788|0|52|504|-80.497332|64|35.667941|FRESH BERRIES|0.0|4|BLUEBERRIES 6 OZ|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00817621010109|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|af790c1806ae892768d33d0d341f45cf93c42fa3|1.1|2014-10-09 13:31:00|80.497482303704658|1||178|35.691507255430857|0|6|524|-80.861571|64|35.444615|FRESH PROD FRESH ONIONS|0.0|4|COO YELLOW ONIONS, LRG|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00204665000003|FRESH PRODUCE|PRODUCE|-80.497332|80.497447600120879|340|1
35.667941|afbdfa8c7d6fc2d651e7c94b8a0e047c35da1feb|2.39|2015-01-03 15:55:00|80.497482303704658|1|7203695175|178|35.691507255430857|0|6|1607|-80.861571|371|35.444615|FROZEN DOUGH (BREAD)|0.0|14|FRESH LRG FRENCH BREAD|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00072036951755|BREAD|BAKERY|-80.497332|80.497447600120879|340|1
35.667941|dd6b443fc91f356086e4a2e8607981edf1006161|4.19|2014-10-12 11:58:00|80.497482303704658|1|4812110208|178|35.69150730682852|0|6|1037|-80.860108|164|35.500972|ENGLISH MUFFINS|2.09|7|THOMAS ENG MUFFN ORIG 6 PK PP|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00048121102081|BREAKFAST|COMMERCIAL BAKERY|-80.497332|80.497430447440678|268|1
35.667941|f6694375f3c7cbb9933c1b56aa9ec3f6ba66913f|13.29|2014-12-09 12:41:00|80.497482303704658|1|3700013882|178|35.69150730682852|0|6|389|-80.860108|66|35.500972|NFS-LAUNDRY DETERGENTS|0.0|1|TIDE ORIGINAL W/BLEACH|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00037000875468|DETERGENTS|G1 GROCERY|-80.497332|80.497430447440678|268|1
35.667941|08082fa14b6da0abd7100229d2ec4382087bff16|13.29|2015-01-11 13:00:00|80.497482303704658|1|3700013882|178|35.691507293415832|0|6|389|-80.762919|66|35.442529|NFS-LAUNDRY DETERGENTS|0.0|1|TIDE ORIGINAL W/BLEACH|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00037000875468|DETERGENTS|G1 GROCERY|-80.497332|80.49743519887393|471|1
35.667941|bc65571bc7b72cc67e87b95b4ed0b839aa639388|13.29|2014-12-27 11:44:00|80.497482303704658|1|3700013882|178|35.69150730682852|0|6|389|-80.860108|66|35.500972|NFS-LAUNDRY DETERGENTS|0.0|1|TIDE ORIGINAL W/BLEACH|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00037000875468|DETERGENTS|G1 GROCERY|-80.497332|80.497430447440678|268|1
35.667941|2a8888242e208ac7623a58d211f594f72b3b58b7|2.39|2014-11-18 10:59:00|1.4057311447477159|1|4132100541|178|0.6225230078570788|0|52|184|-80.497332|28|35.667941|SALAD DRESSINGS-LIQUID|0.39|1|D WISHBONE DRS VIN ROMANO BAS|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00041000078354|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|d9a0643e1e1b9beae94921dfe38c500cf8bdcacb|2.19|2014-10-16 16:48:00|80.497482303704658|1|4300028543|178|35.691507363803225|0|6|28|-80.875654|26|35.585842|STUFFING PRODUCTS|0.0|1|STOVE TOP STUFFING CORNBREAD|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00043000285329|PREPARED FOODS-DRY MIXES|G1 GROCERY|-80.497332|80.497406980099072|99|1
35.667941|8f13e9e9ef7dc3b2e0737ddfeb6000dc884465b8|2.99|2015-01-29 14:50:00|1.4057311447477159|1|4667716832|178|0.6225230078570788|0|52|6133|-80.497332|1546|35.667941|BULB-CARD DECO-FLAME-SML BSE|0.0|18|PHILIP 25W DURAMAX SM FLAM CLR|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00046677168322|LIGHT BULBS/ELECTRICAL|GM|-80.497332|1.4049434824709919|178|1
35.667941|6b12b5cf6bc3330f35adee7c3d6a4ef8ebefab7f|5.49|2014-10-07 17:24:00|80.497482303704658|1|7203660022|178|35.69150730682852|0|6|355|-80.860108|104|35.500972|FRESH GRILLING SAUSAGE|0.0|19|HT HOT ITALIAN SAUSAGE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00072036600233|DINNER SAUSAGE|CASE READY MEATS|-80.497332|80.497430447440678|268|1
35.667941|098638d2326b7aa690fc9d3f765360dfdb244cab|2.19|2014-12-16 13:22:00|1.4057311447477159|1|7418226090|178|0.6225230078570788|0|52|722|-80.497332|73|35.667941|NFS-HAND SOAPS|0.0|1|SS HAND COUNTRY DESIGNS|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00074182260125|PERSONAL SOAP/BATH ADDITIVES|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|8ca94b5f97b00e1290ca87aad1ae1007f93596f8|3.99|2014-11-08 12:40:00|1.4057311447477159|1|4900005235|178|0.6225230078570788|0|52|55|-80.497332|8|35.667941|REGULAR|0.99|23|SCHWEPPES 7.5 OZ|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00078000009767|CARBONATED BEVERAGES|BEVERAGE|-80.497332|1.4049434824709919|178|1
35.667941|094b995bb492893396a0e050e25ecf69f5790f51|3.99|2014-10-28 15:27:00|80.497482303704658|1|4900005235|178|35.69150730682852|0|6|55|-80.860108|8|35.500972|REGULAR|1.0|23|SCHWEPPES 7.5 OZ|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00078000009767|CARBONATED BEVERAGES|BEVERAGE|-80.497332|80.497430447440678|268|1
35.667941|7265d40bb6bcad240efa8ad0d95860ba6cc07058|3.18|2015-03-04 17:48:00|80.497482303704658|1|8190000008|178|35.69150730682852|0|6|1218|-80.860108|273|35.500972|ASIAN OTHER|0.0|1|KOALA COOKIE CHOCOLATE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00081900000086|ASIAN PREP. FOODS|G1 GROCERY|-80.497332|80.497430447440678|268|2
35.667941|07b924bce5ae5a128967fad7b1464fa48eb97799|14.99|2014-12-12 17:28:00|80.497482303704658|1|8912128812|178|35.691507293415832|0|6|9960|-80.762919|887|35.442529|NFS-S/PREM-CAB SAUVIGNON|0.0|13|J  LOHR ESTATES CAB SAUV|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00089121288122|SUPER PREMIUM ($11-$14.99)|WINE|-80.497332|80.49743519887393|471|1
35.667941|8a87b6d0ee2d457866884e75aa444761a88482a9|11.99|2014-12-20 13:32:00|80.497482303704658|1|3700088206|178|35.69150730682852|0|6|426|-80.860108|72|35.500972|NFS-PAPER TOWELS|2.0|1|BOUNTY TOWEL 6 RL SAS WHITE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00037000882022|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.497332|80.497430447440678|268|1
35.667941|4bec550c00c8d662b0fafb6940ea9669c312f642|2.4|2015-03-02 17:11:00|80.497482303704658|1|3663203732|178|35.69150730682852|0|6|685|-80.860108|61|35.500972|GREEK|0.2|3|DANNON LNF GREEK KEY LIME|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00036632037381|YOGURT|DAIRY|-80.497332|80.497430447440678|268|2
35.667941|b242f4637719896202b9930117a8a35d7dedcc38|1.2|2014-12-27 11:38:00|80.497482303704658|1|3663203732|178|35.69150730682852|0|6|685|-80.860108|61|35.500972|GREEK|0.0|3|DANNON LNF GREEK KEY LIME|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00036632037381|YOGURT|DAIRY|-80.497332|80.497430447440678|268|1
35.667941|b9451e9b976d864d845fd5d94b5a71c60e1cc4b2|11.99|2014-10-09 15:58:00|1.4057311447477159|1|3700088206|178|0.6225230078570788|0|52|426|-80.497332|72|35.667941|NFS-PAPER TOWELS|2.0|1|BOUNTY TOWEL 6 RL SAS WHITE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00037000882022|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|a0f038644d00ce9fdc2cc26c9db9f871f13df520|11.99|2014-11-19 13:14:00|1.4057311447477159|1|3700088206|178|0.6225230078570788|0|52|426|-80.497332|72|35.667941|NFS-PAPER TOWELS|3.0|1|BOUNTY TOWEL 6 RL SAS WHITE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00037000882022|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|6a3ef10193f62a843d63a08b5e8f1f3de80b62c2|11.99|2014-10-15 15:59:00|1.4057311447477159|1|3700088206|178|0.6225230078570788|0|52|426|-80.497332|72|35.667941|NFS-PAPER TOWELS|6.0|1|BOUNTY TOWEL 6 RL SAS WHITE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00037000882022|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|372856980d49b6c4880258c2f053af12866997f9|2.4|2014-10-22 16:38:00|80.497482303704658|1|3663203732|178|35.691507293415832|0|6|685|-80.762919|61|35.442529|GREEK|0.4|3|DANNON LNF GREEK KEY LIME|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00036632037381|YOGURT|DAIRY|-80.497332|80.49743519887393|471|2
35.667941|dfef69c40ef255be3b5f56464e80ab550d2bc683|5.35|2015-02-27 14:10:00|80.497482303704658|1|3700040152|178|35.69150730682852|0|6|725|-80.860108|66|35.500972|NFS-DISHWASHING LIQUID|0.0|1|CASCADE GEL DAWN FRESH SCENT|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00037000401520|DETERGENTS|G1 GROCERY|-80.497332|80.497430447440678|268|1
35.667941|40b459098fd104a4e9560153aea8484ef1eb2adc|4.58|2014-11-14 15:49:00|80.497482303704658|1|4118804070|178|35.691507293415832|0|6|257|-80.762919|39|35.442529|TOMATOES|0.58|1|FURMANO TOMATO WHL 28|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00041188040662|VEGETABLES-CAN/JAR|G1 GROCERY|-80.497332|80.49743519887393|471|2
35.667941|30552e6023e62dea97d0064751bb8e3cb1de47e2|1.97|2015-02-05 17:57:00|80.497482303704658|1|7203697723|178|35.691507293415832|0|6|223|-80.762919|35|35.442529|SUGAR SUBSTITUTES|0.0|1|HT SWEETENER - SUCRALOSE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00072036977236|SUGAR/SUBSTITUTES|G1 GROCERY|-80.497332|80.49743519887393|471|1
35.667941|468477a4fa893aff6c969028cab7c2f2ad433d57|3.94|2014-11-08 13:26:00|80.497482303704658|1|7203697723|178|35.69150730682852|0|6|223|-80.860108|35|35.500972|SUGAR SUBSTITUTES|0.0|1|HT SWEETENER - SUCRALOSE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00072036977236|SUGAR/SUBSTITUTES|G1 GROCERY|-80.497332|80.497430447440678|268|2
35.667941|18f1d26c6b63e42d61189a244a8631df0dd20f42|1.97|2014-09-27 17:18:00|80.497482303704658|1|7203697723|178|35.69150730682852|0|6|223|-80.860108|35|35.500972|SUGAR SUBSTITUTES|0.0|1|HT SWEETENER - SUCRALOSE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00072036977236|SUGAR/SUBSTITUTES|G1 GROCERY|-80.497332|80.497430447440678|268|1
35.667941|98232e333f8abcb829b19cc7655daecee116345a|6.99|2014-09-18 15:12:00|1.4057311447477159|1|7203695357|178|0.6225230078570788|0|52|1295|-80.497332|383|35.667941|PIES PASTRY CASE TAX|0.0|14|"9"" KEY LIME PIE"|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00072036953575|PASTRY CASE|BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|b73eab674e242b73dcf315c927356c903b6e8149|2.59|2014-11-07 15:22:00|1.4057311447477159|1|7203695278|178|0.6225230078570788|0|52|1654|-80.497332|381|35.667941|DESSERT CAKES|0.0|14|DOUBLE FUDGE CAKE SLICE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00072036952783|CAKES|BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|e8de5c2258551241ae85dcfc6367bcedf5734fac|4.29|2015-02-14 15:21:00|80.497482303704658|1|4400003538|178|35.69150730682852|0|6|90|-80.860108|13|35.500972|SNACK CRACKERS|0.0|1|STONED WHEAT THINS|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00044000035389|CRACKERS|G1 GROCERY|-80.497332|80.497430447440678|268|1
35.667941|a6a29b30d9877a2742efcd01ed9d8d3c23725599|1.99|2014-12-23 16:58:00|80.497482303704658|1|4900004574|178|35.69150730682852|0|6|171|-80.860108|20|35.500972|ISOTONIC DRINKS|1.2|1|POWERADE LEMON LIME|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00049000045734|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.497332|80.497430447440678|268|1
35.667941|d968a17c16c3ef3773d740eccd10f9968fb0fce3|5.97|2014-12-20 08:22:00|80.497482303704658|1|7203676359|178|35.69150730682852|0|6|345|-80.860108|57|35.500972|ORGANIC MILK|0.0|3|HTO ORGANIC 2% MILK GAL|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00072036763600|MILK|DAIRY|-80.497332|80.497430447440678|268|1
35.667941|f42f0ee81fd4dde1b4aba381b9d0acb290f6f4b0|6.27|2015-02-23 17:05:00|80.497482303704658|1|7203676359|178|35.691507255430857|0|6|345|-80.861571|57|35.444615|ORGANIC MILK|0.0|3|HTO ORGANIC 2% MILK GAL|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00072036763600|MILK|DAIRY|-80.497332|80.497447600120879|340|1
35.667941|c02a593acd54e9f22d6597c2693c291320ea4c6c|6.47|2015-01-07 14:15:00|80.497482303704658|1|7203676359|178|35.691507293415832|0|6|345|-80.762919|57|35.442529|ORGANIC MILK|0.0|3|HTO ORGANIC 2% MILK GAL|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00072036763600|MILK|DAIRY|-80.497332|80.49743519887393|471|1
35.667941|fa38a56db98e978aacf5db4936bfc92473ca9497|5.97|2014-12-04 15:11:00|80.497482303704658|1|7203676359|178|35.691507255430857|0|6|345|-80.861571|57|35.444615|ORGANIC MILK|0.0|3|HTO ORGANIC 2% MILK GAL|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00072036763600|MILK|DAIRY|-80.497332|80.497447600120879|340|1
35.667941|2842e39f8ef7c301a1c12855252d85d7ad6fb07f|4.99|2014-12-01 10:30:00|1.4057311447477159|1|1111018700|178|0.6225230078570788|0|52|1647|-80.497332|379|35.667941|PACKAGED MUFFINS|1.02|14|FFM 4 CT BLUEBERRY MUFFIN|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00011110187000|MUFFINS|BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|97ace677d06990130250a8dd9cdcba871ea63fa1|6.49|2014-09-28 12:14:00|80.497482303704658|1|1480000039|178|35.69150730682852|0|6|128|-80.860108|20|35.500972|APPLE JUICE-SHELF|1.0|1|MOTTS APPLE JUICE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00014800000399|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.497332|80.497430447440678|268|1
35.667941|6b73ae4c75bc6e4779cf40b0be1376ca52e5fcc9|3.35|2015-01-17 16:15:00|80.497482303704658|1|1600042040|178|35.691507293415832|0|6|13|-80.762919|2|35.442529|ROLLS/BISCUIT MIXES|0.0|1|BC BISQUICK|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00016000420403|BAKING MIXES|G1 GROCERY|-80.497332|80.49743519887393|471|1
35.667941|e6693929d1adbc013434929766d7e3bcf1b480ac|2.69|2015-02-16 13:50:00|80.497482303704658|1|1600015110|178|35.691507255430857|0|6|205|-80.861571|31|35.444615|REMAINING SNACKS|0.0|1|CHEX SNACK MIX - PEANUT LOVERS|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00016000158108|SNACKS|G1 GROCERY|-80.497332|80.497447600120879|340|1
35.667941|6fa2b23fde97ade136b90700d97b122760f746ae|4.65|2014-12-05 15:47:00|80.497482303704658|1|95952|178|35.69150730682852|0|6|1596|-80.860108|369|35.500972|NFS OTHER|0.0|22|CARAMEL BRULEE LATTE GRANDE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00000000959520|NFS STARBUCKS|COFFEE SHOP|-80.497332|80.497430447440678|268|1
35.667941|1be485e244c54d48e69e3767370ddf5dd80ea03f|12.99|2015-02-09 12:17:00|1.4057311447477159|1|8500001658|178|0.6225230078570788|0|52|9963|-80.497332|887|35.667941|NFS-S/PREM-PINOT GRIS/GR|0.0|13|DA VINCI PINOT GRIGIO 750 ML|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00085000016589|SUPER PREMIUM ($11-$14.99)|WINE|-80.497332|1.4049434824709919|178|1
35.667941|848b0015084dc67b51f2644dd3687299c7d6dd99|12.99|2014-12-18 16:19:00|1.4057311447477159|1|8500001658|178|0.6225230078570788|0|52|9963|-80.497332|887|35.667941|NFS-S/PREM-PINOT GRIS/GR|0.0|13|DA VINCI PINOT GRIGIO 750 ML|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00085000016589|SUPER PREMIUM ($11-$14.99)|WINE|-80.497332|1.4049434824709919|178|1
35.667941|4dca8d9216c5e38d1ac2d4c8e138e649ec0fc542|5.49|2014-12-29 14:44:00|1.4057311447477159|1|827411111|178|0.6225230078570788|0|52|55|-80.497332|8|35.667941|REGULAR|1.5|23|VIRGILS BLACK CHERRY CREAM|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00090341231157|CARBONATED BEVERAGES|BEVERAGE|-80.497332|1.4049434824709919|178|1
35.667941|b9cf275fb662b97b53600da0f9b58ba974ace390|6.99|2014-10-04 12:30:00|1.4057311447477159|1|7255400153|178|0.6225230078570788|0|52|273|-80.497332|43|35.667941|PREMIUM NOVELTIES|0.0|5|NESTLE DRUMSTICK VANILLA 8 CT|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00072554001543|FROZEN NOVELTIES|FROZEN|-80.497332|1.4049434824709919|178|1
35.667941|71b77a1bac7cdc31dc6dcf8f50f44af445c5c085|8.79|2014-09-19 11:37:00|80.497482303704658|1|9955508520|178|35.691507255430857|0|6|37|-80.861571|10|35.444615|PODS/CUPS/SINGLES|0.0|1|CARIBOU BLEND K-CUPS|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00099555089929|COFFEE|G1 GROCERY|-80.497332|80.497447600120879|340|1
35.667941|5e2262a7ebe72a45395a51b9aa73194de1856c25|9.99|2014-10-26 14:52:00|1.4057311447477159|1|8500000843|178|0.6225230078570788|0|52|9951|-80.497332|886|35.667941|NFS-PREM-PINOT GRIS/GRIG|0.0|13|CB-ECCO DOMANI PINOT GRIGIO|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00085000008430|PREMIUM ($8-$10.99)|WINE|-80.497332|1.4049434824709919|178|1
35.667941|1a2dcbbfe5718c1d3e709d1d02ccc435c19229dc|2.78|2015-01-06 15:47:00|1.4057311447477159|1|4150005807|178|0.6225230078570788|0|52|80|-80.497332|34|35.667941|SEASONING PACKETS|0.0|1|FRENCH'S ORIGINAL CHILI-O|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00041500058078|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.497332|1.4049434824709919|178|2
35.667941|d620a78f2c6cfa1cc0fc8c3b61427a8fbfb19763|2.29|2015-01-04 12:27:00|1.4057311447477159|1|2670012915|178|0.6225230078570788|0|52|1267|-80.497332|53|35.667941|DIPS AND SPREADS|0.79|3|DEAN'S FRENCH ONION DIP|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00026700129155|CULTURES|DAIRY|-80.497332|1.4049434824709919|178|1
35.667941|069ea891da4273651e4300e4468a5dea3e1d5978|1.15|2014-09-12 13:36:00|80.497482303704658|1|4920005675|178|35.69150730682852|0|6|224|-80.860108|35|35.500972|SUGAR-BROWN|0.0|1|DOMINO LT BRWN SUGAR-BOX|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00049200056752|SUGAR/SUBSTITUTES|G1 GROCERY|-80.497332|80.497430447440678|268|1
35.667941|a31aedad7f5c66734388834d1b793689bbe7083d|3.99|2014-10-16 11:53:00|1.4057311447477159|1|7203688078|178|0.6225230078570788|0|52|523|-80.497332|64|35.667941|FRESH POTATOES|0.0|4|HT RED POTATO 3LB BAG|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00072036880789|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|5ad6b73ec68a56a2337b5668062c76e74310dd87|19.99|2015-02-27 17:07:00|80.497482303704658|1|20310300000|178|35.69150730682852|0|6|1153|-80.860108|87|35.500972|NFS-FRESH CUT ARRANGE|0.0|9|*CORSAGES|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00203103000001|FLORAL|FLORAL|-80.497332|80.497430447440678|268|1
35.667941|0ed6d527d467f377191f796c02b78a7efcaddfee|7.99|2014-11-12 15:21:00|1.4057311447477159|1|1380014333|178|0.6225230078570788|0|52|1280|-80.497332|48|35.667941|MULTI SERVE MEALS|1.0|5|STOUFFER FM/STYLE GRANDMA CHKN|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00013800190864|FROZEN MEALS|FROZEN|-80.497332|1.4049434824709919|178|1
35.667941|c7296fb25acb6c7d6ef1c4a1b80ff9d77641ab37|7.99|2015-02-21 17:46:00|80.497482303704658|1|30031872120|178|35.69150730682852|0|6|4236|-80.860108|1200|35.500972|DEX ADULT/CHILDREN|0.0|17|ROBITUSSIN DAY COLD+FLU CAPS|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00300318721209|COUGH/COLD/SINUS|HBC|-80.497332|80.497430447440678|268|1
35.667941|2bb22eb0c68e71ec4838a2cea41a388a93bdbe59|2.0|2014-11-13 13:15:00|80.497482303704658|1|7203663118|178|35.69150730682852|0|6|1262|-80.860108|57|35.500972|HALF N HALF WHIPPING CREAM|0.33|3|HT HALF & HALF|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00072036632043|MILK|DAIRY|-80.497332|80.497430447440678|268|1
35.667941|3a7a61949d4685583dbc97f2b71f839a8dd14225|3.99|2014-12-16 17:17:00|80.497482303704658|1|7203602701|178|35.691507293415832|0|6|1878|-80.762919|435|35.442529|HUMMUS|0.5|6|FFM ARTISAN PINE NUT HUMMUS|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00072036027054|SALADS|DELI|-80.497332|80.49743519887393|471|1
35.667941|21abaf397dcfe3787bc2ddac1543a0aa94663248|4.99|2014-10-07 11:24:00|1.4057311447477159|1|3917445141|178|0.6225230078570788|0|52|7221|-80.497332|1600|35.667941|WINTER GLOVES|1.0|18|I/O LADIES CHENILIE GLOVE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00039174451417|SEASONAL MERCHANDISE|GM|-80.497332|1.4049434824709919|178|1
35.667941|df868ff807baf63b1c504043ee10656d9dab0e98|4.49|2015-01-13 10:58:00|1.4057311447477159|1|4470003050|178|0.6225230078570788|0|52|840|-80.497332|102|35.667941|TUBS|0.99|19|OM DELI FRESH ROTISSERE CHCKEN|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00044700030998|LUNCHMEATS|CASE READY MEATS|-80.497332|1.4049434824709919|178|1
35.667941|2908bc234c1964dd7d36407fbff0b3bc8e275383|29.99|2014-11-26 11:12:00|1.4057311447477159|1|20960300000|178|0.6225230078570788|0|52|667|-80.497332|145|35.667941|PARTY PLATTERS|0.0|12|THE ORIGINAL SHRIMP PLATTER|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00209603000008|SHRIMP|SEAFOOD|-80.497332|1.4049434824709919|178|1
35.667941|f73efa78ef51454ac1046bf9e2914b2ba4a6e7ca|1.07|2014-11-23 13:22:00|1.4057311447477159|1||178|0.6225230078570788|0|52|502|-80.497332|64|35.667941|FRESH BANANAS|0.0|4|BANANAS, YELLOW|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00204011000008|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|6094c503138a84d17e7e5db6dbfd9313ffe5f077|1.09|2015-01-22 12:32:00|1.4057311447477159|1||178|0.6225230078570788|0|52|502|-80.497332|64|35.667941|FRESH BANANAS|0.0|4|BANANAS, YELLOW|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00204011000008|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|b120876348cb80e5c5640599428b1261c6e728ca|4.99|2015-02-07 14:03:00|1.4057311447477159|1|71575620002|178|0.6225230078570788|0|52|504|-80.497332|64|35.667941|FRESH BERRIES|1.49|4|STRAWBERRIES 1LB CLAM|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00850806002810|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|ad64a835a71a6446d81ed26ee357c11c2bc8e321|5.99|2015-02-03 16:49:00|1.4057311447477159|1|88831391490|178|0.6225230078570788|0|52|485|-80.497332|101|35.667941|PREMIUM WIENERS|0.0|19|NATHAN'S BUNSIZE BEEF FRANKS|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00888313914906|WIENERS|CASE READY MEATS|-80.497332|1.4049434824709919|178|1
35.667941|f33412d5a4e030359549b72af36b36d9cb9c597c|3.0|2014-10-19 11:58:00|1.4057311447477159|1|7203688157|178|0.6225230078570788|0|52|556|-80.497332|64|35.667941|PACKAGED VEGETABLES|0.0|4|HT RV FRENCH GREEN BEANS|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00072036881595|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.667941|7cc91961d355e4997d714eba90b8d784060d7fe2|1.89|2014-12-21 14:04:00|1.4057311447477159|1|7203695004|178|0.6225230078570788|0|52|1605|-80.497332|371|35.667941|PAR BAKED (BREAD)|0.0|14|SMALL FRENCH BREAD.|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00072036950048|BREAD|BAKERY|-80.497332|1.4049434824709919|178|1
35.667941|38f590ccbaba1463e57532ab4a47dd3d6730d2e5|5.82|2014-10-20 18:08:00|1.4057311447477159|1|20562000000|178|0.6225230078570788|0|52|1823|-80.497332|410|35.667941|BH HAM|0.0|6|BOARS HEAD VIRGINIA HAM|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00205620000007|BH MEAT|DELI|-80.497332|1.4049434824709919|178|1
35.667941|30fce3e6b511a0e2144c98b17cc812b8ee468db3|6.2|2015-01-26 15:17:00|1.4057311447477159|1|68954408130|178|0.6225230078570788|0|52|685|-80.497332|61|35.667941|GREEK|0.0|3|FAGE TOTAL 2% MIXED BERRIES|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00689544081777|YOGURT|DAIRY|-80.497332|1.4049434824709919|178|4
35.667941|6a6e72eb9b4b7755e0ceb28cbc62842f3321fa07|19.99|2015-02-28 17:28:00|80.497482303704658|1|7023666010|178|35.691507255430857|0|6|751|-80.861571|87|35.444615|NFS-BOUQUETS|0.0|9|$19.99  BUZZY BEES BQT|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00070236660101|FLORAL|FLORAL|-80.497332|80.497447600120879|340|1
35.667941|45bb0fc74b58ce4c9ad7c3b201ab2966c6e36de3|2.49|2014-09-17 10:51:00|1.4057311447477159|1|7203697799|178|0.6225230078570788|0|52|6859|-80.497332|1581|35.667941|RE USEABLE EVERYDAY|0.5|18|HT FOLD'NSNAP REUSABLE TOTE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00072036977991|SHOPPING BAGS|GM|-80.497332|1.4049434824709919|178|1
35.667941|578723a2d5e5a23fbd35851379c25d5a15a4fc0a|6.5|2014-11-02 14:49:00|80.497482303704658|1|7203656080|178|35.691507255430857|0|6|318|-80.861571|52|35.444615|SHREDDED/GRATED CHEESE|0.0|3|HT DOUBLE CHEDDAR SHRED|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00072036709271|CHEESE|DAIRY|-80.497332|80.497447600120879|340|2
35.667941|d40ef600bfaa38973f0184e599b762895cd43002|5.5|2015-03-08 17:24:00|80.497482303704658|1|20563200000|178|35.69150730682852|0|6|1823|-80.860108|410|35.500972|BH HAM|0.0|6|BOARS HEAD TAVERN HAM|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00205632000002|BH MEAT|DELI|-80.497332|80.497430447440678|268|1
35.667941|27599577fad0dd2789c2be33b18215433563cedc|2.4|2014-11-17 17:30:00|80.497482303704658|1|3663203732|178|35.69150730682852|0|6|685|-80.860108|61|35.500972|GREEK|0.4|3|DANNON LNF GREEK BLUEBERRY|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00036632037329|YOGURT|DAIRY|-80.497332|80.497430447440678|268|2
35.667941|c442e8efeba16a497259936ad56c7d2d3fde3298|4.39|2014-12-30 12:17:00|1.4057311447477159|1|4400003037|178|0.6225230078570788|0|52|90|-80.497332|13|35.667941|SNACK CRACKERS|2.2|1|WHEAT THINS ORIGINAL|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00044000030377|CRACKERS|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|06fdb0b5d4af59143a4f578c90622f8ff85a5639|7.99|2015-01-07 14:27:00|80.497482303704658|1|38151901250|178|35.691507293415832|0|6|3618|-80.762919|1055|35.442529|WOMEN-PERMANENT COLOR|0.0|17|NICE/EZ ROOT TCHUP 5 MD BROWN|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00381519012471|HAIR COLORING/PERM|HBC|-80.497332|80.49743519887393|471|1
35.667941|0ae4a1dff32f95599b41db3c72ceabdb3ec8aa3f|4.49|2015-02-22 16:36:00|80.497482303704658|1|5100002511|178|35.69150730682852|0|6|1221|-80.860108|275|35.500972|PASTA SC VALUE|0.0|1|PREGO SC 45 TRADITIONAL|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00051000025111|PASTA SAUCES|G1 GROCERY|-80.497332|80.497430447440678|268|1
35.667941|d9a3a4e6d992bbffa4f6432f76d826f0a09a60ee|5.99|2015-01-30 17:25:00|80.497482303704658|1|7055176104|178|35.691507363803225|0|6|2023|-80.875654|505|35.585842|GOAT CHEESE|0.0|6|CHAVRIE MINI GOAT LOG PLAIN|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00070551761040|SPECIALTY CHEESE|DELI|-80.497332|80.497406980099072|99|1
35.667941|6bc4fa1927a04070a7c37f3d73eb8021bce69379|6.99|2015-02-11 16:58:00|80.497482303704658|1|20496000000|178|35.69150730682852|0|6|755|-80.860108|87|35.500972|NFS-BALLOONS|0.0|9|*BALLOONS|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00204960000005|FLORAL|FLORAL|-80.497332|80.497430447440678|268|1
35.667941|26649b25700cc053eb7015f4130e900c80652575|10.3|2014-09-10 14:28:00|1.4057311447477159|1|7218063473|178|0.6225230078570788|0|52|254|-80.497332|892|35.667941|PREMIUM PIZZA|4.3|5|RED BARON THN CRUST 5 CHEESE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00072180633217|FROZEN PIZZA|FROZEN|-80.497332|1.4049434824709919|178|2
35.667941|da12193b48486d11399055ada91e9c78cc8be1c9|3.89|2014-12-09 14:39:00|80.497482303704658|1|4400003219|178|35.691507219599117|0|6|1249|-80.86175|12|35.40953|CHOCOLATE CHIP COOKIES|0.89|1|CHIPS AHOY CHEWY REESES CHOCO|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00044000033880|COOKIES|G1 GROCERY|-80.497332|80.497458186177482|209|1
35.667941|c2e06bb43e91d45c8596d29173288c9b26ab6ddf|7.59|2014-11-26 18:57:00|80.497482303704658|1|1583902020|178|35.691507293415832|0|6|204|-80.762919|31|35.442529|TORTILLA CHIPS|0.0|1|D GRDN OF EATIN CHIPS BLUE CRN|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|35.699188602026126|00015839020204|SNACKS|G1 GROCERY|-80.497332|80.49743519887393|471|1
35.667941|6aea62cf8efa30c566e15e88f1d708b06e277064|4.69|2015-01-18 13:29:00|1.4057311447477159|1|5100007620|178|0.6225230078570788|0|52|264|-80.497332|307|35.667941|DESSERT CAKES FROZEN|0.0|5|PEP FARM LEMON 3-LAYER CAKE|9e638964fad2e55f788801b57bf999fa9fbedc04|1.6283842662540275|0.6209993146566879|00051000174239|DESSERTS FROZEN|FROZEN|-80.497332|1.4049434824709919|178|1
35.17739|edf8225a3d3523eba6c342021b7ac94330d8688d|11.04|2014-10-21 18:23:00|80.801203185414451|4|20165700000|208|35.210562645413894|0|24|297|-80.739|49|35.141204|GROUND BEEF|1.31|2|HT GROUND BEEF CHUCK 80% LEAN|a22708a09b050e5283398c704e0e928cebc6de17|2.2921496990843884|35.194272495053255|00201657000003|BEEF|MEAT|-80.80146|80.801463802172094|171|2
35.17739|d7d3b6f1015f050212567548f101738e9a064c16|1.99|2015-02-11 13:54:00|80.801203185414451|4|7203648011|208|35.210562642904875|0|24|274|-80.810056|44|35.219587|ICE|0.0|5|HT BAGGED ICE 10LB (456)|a22708a09b050e5283398c704e0e928cebc6de17|2.2921496990843884|35.194272495053255|00000000004560|ICE|FROZEN|-80.80146|80.801476239345121|401|1
35.17739|f469a8540c1b6d66463c8457c417d254559ccf26|4.85|2014-12-31 15:47:00|80.801203185414451|4|7790011553|208|35.210562645413894|0|24|361|-80.739|105|35.141204|BREAKFAST SAUSAGE|1.51|19|JIMMY DEAN MILD SAUSAGE|a22708a09b050e5283398c704e0e928cebc6de17|2.2921496990843884|35.194272495053255|00077900115530|BREAKFAST SAUSAGE|CASE READY MEATS|-80.80146|80.801463802172094|171|1
35.17739|beb68d908a830888754e90960620e5b2f8ce1fbf|5.29|2014-10-22 18:57:00|80.801203185414451|4|31254742825|208|35.210562645413894|0|24|4030|-80.739|1080|35.141204|ORAL RINSE-ANTISEPTIC|0.0|17|LISTERINE ORIGINAL MW NB|a22708a09b050e5283398c704e0e928cebc6de17|2.2921496990843884|35.194272495053255|00312547701310|ORAL HYGIENE|HBC|-80.80146|80.801463802172094|171|1
35.17739|b870017f453e0d565bc057f6647e27a1fa0d90d6|4.39|2014-11-19 15:09:00|80.801203185414451|4|5480001008|208|35.210562645413894|0|24|239|-80.739|38|35.141204|RICE-PACKAGED & BULK|0.0|1|UNCLE BENS RICE CONVERTED 32|a22708a09b050e5283398c704e0e928cebc6de17|2.2921496990843884|35.194272495053255|00054800010080|RICE GRAINS AND BEANS|G1 GROCERY|-80.80146|80.801463802172094|171|1
35.17739|9a965e28eb92e510fe8959a9e143880501fda01f|16.29|2014-09-27 15:31:00|80.801203185414451|4|20188200000|208|35.210562645413894|0|24|299|-80.739|49|35.141204|ANGUS BEEF|0.0|2|ANGUS BEEF BNLS CHUCK STEAK|a22708a09b050e5283398c704e0e928cebc6de17|2.2921496990843884|35.194272495053255|00201882000007|BEEF|MEAT|-80.80146|80.801463802172094|171|2
35.17739|08fc6c2d2cc7a246438dc0633ae4af8b5c57f762|5.18|2014-10-13 17:52:00|80.801203185414451|4|5100013279|208|35.210562645413894|0|24|214|-80.739|33|35.141204|BROTH|0.59|1|SWANSON BROTH CHICKEN|a22708a09b050e5283398c704e0e928cebc6de17|2.2921496990843884|35.194272495053255|00051000121141|SOUP|G1 GROCERY|-80.80146|80.801463802172094|171|2
35.17739|cf315b2a3c99626857ea83dbe7304ee4bff1d008|4.99|2015-02-19 13:58:00|80.801203185414451|4|2840015282|208|35.210562645413894|0|24|203|-80.739|31|35.141204|CHEESE SNACKS|1.0|1|CHEETOS CRUNCHY PARTY SIZE|a22708a09b050e5283398c704e0e928cebc6de17|2.2921496990843884|35.194272495053255|00028400152822|SNACKS|G1 GROCERY|-80.80146|80.801463802172094|171|1
35.17739|25a396e7d7b6e7b4b2481e52a1838f6dd397df1f|15.19|2014-09-24 12:13:00|80.801203185414451|4|31284353642|208|35.210562645413894|0|24|4308|-80.739|1205|35.141204|ASPIRIN|0.0|17|BAYER ASPIRIN REGIMEN 81MG|a22708a09b050e5283398c704e0e928cebc6de17|2.2921496990843884|35.194272495053255|00312843536425|PAIN RELIEF|HBC|-80.80146|80.801463802172094|171|1
35.06858|892a0477ef433d4d3fa654bac34b7d155b8cd717|4.8|2014-11-17 14:31:00|80.700712769248256|4||273|35.089824597403002|0|42|529|-80.709466|64|35.124987|FRESH ASPARAGUS|2.67|4|GREEN  ASPARAGUS|a42e0ced139b2e34614eec497926445d050ab1ad|1.467950597192485|35.088667338853092|00204080000008|FRESH PRODUCE|PRODUCE|-80.7007|80.7007142291544|157|1
35.06858|a1dc27c0e9f7b807a2017b28f39377cf8eb5e859|1.55|2014-11-07 11:04:00|80.700712769248256|4|78616201000|273|35.089824600594206|0|42|31|-80.732725|4|35.082768|NON CARBONATED WATER|0.55|1|VIT WATER ZERO GLOW 20 OZ|a42e0ced139b2e34614eec497926445d050ab1ad|1.467950597192485|35.088667338853092|00786162003324|BOTTLED WATER|G1 GROCERY|-80.7007|80.700700073444651|147|1
35.06858|dc4dc0c2e4aeecfbf767abed0583bdc117fe4b1c|2.29|2014-10-03 13:27:00|80.700712769248256|4|5100000524|273|35.089824597403002|0|42|1201|-80.709466|33|35.124987|RTS CANNED|0.79|1|CHUNKY HR CHICKEN NOODLE|a42e0ced139b2e34614eec497926445d050ab1ad|1.467950597192485|35.088667338853092|00051000167750|SOUP|G1 GROCERY|-80.7007|80.7007142291544|157|1
35.06858|eb32a419d3d5f7586bd6c40e4f2aea2cc8b5eded|2.29|2014-09-18 16:59:00|80.700712769248256|4|88937912601|273|35.089824597403002|0|42|80|-80.709466|34|35.124987|SEASONING PACKETS|0.29|1|RED FORK SC LEM HERB ASPARAGUS|a42e0ced139b2e34614eec497926445d050ab1ad|1.467950597192485|35.088667338853092|00889379126012|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.7007|80.7007142291544|157|1
35.06858|71a7ba43cd1e0f73e8aa4889a44db7e71d54e62f|1.55|2014-09-19 15:53:00|80.700712769248256|4|7203663214|273|35.089824597403002|0|42|330|-80.709466|55|35.124987|EGGS|0.0|3|HT GRADE A    EX-LARGE EGGS|a42e0ced139b2e34614eec497926445d050ab1ad|1.467950597192485|35.088667338853092|00072036632142|EGGS FRESH|DAIRY|-80.7007|80.7007142291544|157|1
35.06858|391f8c20f114367e1928784dc748da1171a6d584|1.99|2014-12-10 16:23:00|80.700712769248256|4|7127923100|273|35.089824597403002|0|42|555|-80.709466|64|35.124987|PACKAGED SALADS|0.0|4|F.E. BABY SPRING SALAD MIX|a42e0ced139b2e34614eec497926445d050ab1ad|1.467950597192485|35.088667338853092|00071279231006|FRESH PRODUCE|PRODUCE|-80.7007|80.7007142291544|157|1
35.06858|574e9dea3fc057e81c77f385da3c994a621fdf08|3.49|2014-10-22 15:27:00|80.700712769248256|4|7341013546|273|35.089824597403002|0|42|1035|-80.709466|163|35.124987|SANDWICH ROLL|1.74|7|ARN FLX & FIBR SNDWCH THINS PP|a42e0ced139b2e34614eec497926445d050ab1ad|1.467950597192485|35.088667338853092|00073410135341|BUNS/ROLLS|COMMERCIAL BAKERY|-80.7007|80.7007142291544|157|1
35.06858|0f6017b1312f5587d173ba2f3dce58d07561aab3|1.77|2014-09-27 15:02:00|80.700712769248256|4|7203639031|273|35.089824597403002|0|42|228|-80.709466|36|35.124987|TABLE SYRUP|0.0|1|HT LITE SYRUP|a42e0ced139b2e34614eec497926445d050ab1ad|1.467950597192485|35.088667338853092|00072036390318|TABLE SYRUPS|G1 GROCERY|-80.7007|80.7007142291544|157|1
35.06858|fc9b4d033bc5bb04621a91b3ce702a3f86cdebd1|1.39|2014-10-13 17:25:00|80.700712769248256|4|1254661959|273|35.089824600592173|0|42|48|-80.64817|7|35.04711|REGISTER GUM|0.39|1|TRIDENT SPEARMINT|a42e0ced139b2e34614eec497926445d050ab1ad|1.467950597192485|35.088667338853092|00012546615310|CANDY|G1 GROCERY|-80.7007|80.700700367462787|129|1
35.06858|72452f0d39dfb9ea37d89a81d7b1a683805f8c1e|1.75|2014-09-24 13:13:00|80.700712769248256|4|2920000212|273|35.089824597403002|0|42|149|-80.709466|23|35.124987|WHSE PASTA CORE|0.87|1|MUELLER POT SZ WG THIN SPAG|a42e0ced139b2e34614eec497926445d050ab1ad|1.467950597192485|35.088667338853092|00029200908091|PASTA|G1 GROCERY|-80.7007|80.7007142291544|157|1
35.06858|2906d3cd7879457881afe2957fdda4b63b424bbd|3.39|2014-12-11 13:31:00|80.700712769248256|4|5000012734|273|35.089824597403002|0|42|341|-80.709466|57|35.124987|CREAMERS|0.89|3|COFFEEMATE FF HAZELNUT|a42e0ced139b2e34614eec497926445d050ab1ad|1.467950597192485|35.088667338853092|00050000127344|MILK|DAIRY|-80.7007|80.7007142291544|157|1
35.06858|cb3f565f9734cc260309ff2b426d6c0a1ee35d56|5.52|2014-12-31 18:26:00|80.700712769248256|4|20944900000|273|35.089824596982034|0|42|884|-80.739|145|35.141204|COOKED|1.38|12|SHRIMP CKD TAIL-ON 61/70 (TH)|a42e0ced139b2e34614eec497926445d050ab1ad|1.467950597192485|35.088667338853092|00209449000002|SHRIMP|SEAFOOD|-80.7007|80.700715138571013|171|1
35.06858|b7593463cf987f0fb272bfeb2250b92f90b106e1|1.27|2014-12-17 09:53:00|80.700712769248256|4|7203615012|273|35.089824597403002|0|42|119|-80.709466|17|35.124987|RAISINS|0.0|1|HT RAISINS 6PK|a42e0ced139b2e34614eec497926445d050ab1ad|1.467950597192485|35.088667338853092|00072036150127|FRUIT-DRIED|G1 GROCERY|-80.7007|80.7007142291544|157|1
35.06858|6d1d1ae62998a2f7c66ae3f51b51fac57d2bb2cc|2.0|2014-12-07 16:00:00|80.700712769248256|4|7203669026|273|35.089824597403002|0|42|4054|-80.709466|1080|35.124987|TOOTH BRUSH-PRIVATE LABEL|0.0|17|HT GEM GRIP SOFT TBRUSH|a42e0ced139b2e34614eec497926445d050ab1ad|1.467950597192485|35.088667338853092|00072036690265|ORAL HYGIENE|HBC|-80.7007|80.7007142291544|157|2
35.06858|27080152d6598a0b5a7faa61509d727877817eda|3.99|2014-10-07 13:08:00|80.700712769248256|4|7203663995|273|35.089824597403002|0|42|342|-80.709466|57|35.124987|FRESH MILK|0.0|3|HARRIS TEETER WHOLE MILK|a42e0ced139b2e34614eec497926445d050ab1ad|1.467950597192485|35.088667338853092|00072036639950|MILK|DAIRY|-80.7007|80.7007142291544|157|1
35.06858|6d18ab21cc22056bca793b6eead207e9445fd04b|3.99|2014-11-12 13:17:00|80.700712769248256|4|7203663995|273|35.089824597403002|0|42|342|-80.709466|57|35.124987|FRESH MILK|0.0|3|HARRIS TEETER WHOLE MILK|a42e0ced139b2e34614eec497926445d050ab1ad|1.467950597192485|35.088667338853092|00072036639950|MILK|DAIRY|-80.7007|80.7007142291544|157|1
35.06858|7e5ee2252e628a6381a3b4e58804d3363eb3b949|7.5|2014-11-03 14:52:00|80.700712769248256|4|7203697755|273|35.089824597403002|0|42|81|-80.709466|9|35.124987|RTE CEREAL KIDS|2.5|1|HT CER CINNI MINI CRUNCH|a42e0ced139b2e34614eec497926445d050ab1ad|1.467950597192485|35.088667338853092|00072036979896|CEREAL|G1 GROCERY|-80.7007|80.7007142291544|157|3
35.06858|b19d9770f9d82233fdebd918f4ca06f6bef9ce69|5.0|2014-10-08 13:36:00|80.700712769248256|4|7203697755|273|35.089824597403002|0|42|81|-80.709466|9|35.124987|RTE CEREAL KIDS|1.06|1|HT CER CINNI MINI CRUNCH|a42e0ced139b2e34614eec497926445d050ab1ad|1.467950597192485|35.088667338853092|00072036979896|CEREAL|G1 GROCERY|-80.7007|80.7007142291544|157|2
35.000049|2eb22e0f028dc96d3d4ea596b2f7f0b94cecdba0|3.0|2014-09-24 16:31:00|80.699698036522989|1||249|35.035225585294562|0|18|1617|-80.8062|373|35.037115|ROLLS BULK|0.0|14|BULK ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036955555|ROLLS|BAKERY|-80.699686|80.699690085658418|27|4
35.000049|23169dba1ca6fd4de330e0123c8aaffb16440437|3.0|2014-11-30 17:10:00|1.4091206135396188|1||249|0.6108660934093487|0|47|1617|-80.699686|373|35.000049|ROLLS BULK|0.0|14|BULK ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00072036955555|ROLLS|BAKERY|-80.699686|1.4084752260255726|249|4
35.000049|d6892c14e0923d7d468cb99700eda79d15a9b4ae|3.0|2014-09-28 14:42:00|1.4091206135396188|1||249|0.6108660934093487|0|47|1617|-80.699686|373|35.000049|ROLLS BULK|0.0|14|BULK ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00072036955555|ROLLS|BAKERY|-80.699686|1.4084752260255726|249|4
35.000049|ee13bc809522d0b1d267f171cc6ad640f49aa094|3.0|2015-02-15 18:03:00|80.699698036522989|1||249|35.035225576227809|0|18|1617|-80.64817|373|35.04711|ROLLS BULK|0.0|14|BULK ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036955555|ROLLS|BAKERY|-80.699686|80.699717108215381|129|4
35.000049|78ed389340789d13d76177d6ead45e7ac02d2186|1.5|2015-02-16 14:23:00|80.699698036522989|1||249|35.035225578015265|0|18|1617|-80.824767|373|35.116751|ROLLS BULK|0.0|14|BULK ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036955555|ROLLS|BAKERY|-80.699686|80.699713932630658|294|2
35.000049|4d7fde199d29d6d5bde0504a82f065baffbd5368|3.0|2014-09-13 15:37:00|80.699698036522989|1||249|35.035225576227809|0|18|1617|-80.64817|373|35.04711|ROLLS BULK|0.0|14|BULK ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036955555|ROLLS|BAKERY|-80.699686|80.699717108215381|129|4
35.000049|2eb7ad30a2d9b81c0c5d66785380cb1fce38db1d|4.5|2014-10-02 16:18:00|80.699698036522989|1||249|35.035225585294562|0|18|1617|-80.8062|373|35.037115|ROLLS BULK|0.0|14|BULK ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036955555|ROLLS|BAKERY|-80.699686|80.699690085658418|27|6
35.000049|ddd71631182e4fb9d87712945f7023c7c5ac7ab8|4.5|2014-10-20 16:11:00|80.699698036522989|1||249|35.035225585294562|0|18|1617|-80.8062|373|35.037115|ROLLS BULK|0.0|14|BULK ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036955555|ROLLS|BAKERY|-80.699686|80.699690085658418|27|6
35.000049|3718d01faeef006033f3b003e45c5c66a45c87fd|2.59|2015-01-06 16:12:00|80.699698036522989|1|7203695278|249|35.035225585443811|0|18|1654|-80.760919|381|35.024332|DESSERT CAKES|0.0|14|DOUBLE FUDGE CAKE SLICE|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036952783|CAKES|BAKERY|-80.699686|80.699687018251439|343|1
35.000049|11b84ec9fa7c79c065895290b828175c2dfc52b0|6.0|2015-03-02 17:25:00|80.699698036522989|1||249|35.035225585294562|0|18|1617|-80.8062|373|35.037115|ROLLS BULK|0.41|14|BULK ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036955555|ROLLS|BAKERY|-80.699686|80.699690085658418|27|8
35.000049|c4fa800e006bb439bba0fd558f6adad4523725f5|3.0|2014-12-02 16:50:00|80.699698036522989|1||249|35.035225576227809|0|18|1617|-80.64817|373|35.04711|ROLLS BULK|0.0|14|BULK ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036955555|ROLLS|BAKERY|-80.699686|80.699717108215381|129|4
35.000049|d0d62b8b3d776cd953282dba09f1f2a832fd2992|4.5|2014-11-09 09:40:00|1.4091206135396188|1||249|0.6108660934093487|0|47|1617|-80.699686|373|35.000049|ROLLS BULK|0.0|14|BULK ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00072036955555|ROLLS|BAKERY|-80.699686|1.4084752260255726|249|6
35.000049|b34aa3f31da336227eec6afbe7e943cd33090251|3.0|2015-02-02 17:20:00|80.699698036522989|1||249|35.035225585294562|0|18|1617|-80.8062|373|35.037115|ROLLS BULK|0.0|14|BULK ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036955555|ROLLS|BAKERY|-80.699686|80.699690085658418|27|4
35.000049|5c188cdb101dcf599c5d7db4914276b67ee4fac4|2.25|2015-01-27 15:50:00|80.699698036522989|1||249|35.035225585294562|0|18|1617|-80.8062|373|35.037115|ROLLS BULK|0.0|14|BULK ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036955555|ROLLS|BAKERY|-80.699686|80.699690085658418|27|3
35.000049|6cb2d3cf00063cc76e7d1355a5dcb7dfaf249715|3.0|2014-09-18 16:23:00|1.4091206135396188|1||249|0.6108660934093487|0|47|1617|-80.699686|373|35.000049|ROLLS BULK|0.0|14|BULK ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00072036955555|ROLLS|BAKERY|-80.699686|1.4084752260255726|249|4
35.000049|2cda157d0e6ec4aeaff74cbbfe75b5856d4431ec|2.59|2014-10-05 16:38:00|1.4091206135396188|1|7203695278|249|0.6108660934093487|0|47|1654|-80.699686|381|35.000049|DESSERT CAKES|0.0|14|DOUBLE FUDGE CAKE SLICE|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00072036952783|CAKES|BAKERY|-80.699686|1.4084752260255726|249|1
35.000049|a0837ab0dc93e4a496955c695ceafc6bbb7645b9|6.0|2015-02-23 12:41:00|80.699698036522989|1||249|35.035225578015265|0|18|1617|-80.824767|373|35.116751|ROLLS BULK|0.0|14|BULK ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036955555|ROLLS|BAKERY|-80.699686|80.699713932630658|294|8
35.000049|0c08ba9b45e12bfa06d07896afa3a6eea06f9e6c|2.59|2015-01-15 15:59:00|80.699698036522989|1|7203695298|249|35.035225585443811|0|18|1654|-80.760919|381|35.024332|DESSERT CAKES|0.0|14|OLD FASHION FUDGE CAKE SLICE|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036952981|CAKES|BAKERY|-80.699686|80.699687018251439|343|1
35.000049|5c1290b67b06ed7cc27d58797a5f4efd0820b353|5.99|2014-12-12 18:52:00|80.699698036522989|1|7203695897|249|35.035225585443811|0|18|1654|-80.760919|381|35.024332|DESSERT CAKES|0.0|14|2 CT. TIRAMISU|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036958976|CAKES|BAKERY|-80.699686|80.699687018251439|343|1
35.000049|98b8dda1645ca75a3ec4df5a9fb3ed53b435033b|1.5|2014-09-29 16:20:00|80.699698036522989|1||249|35.035225585294562|0|18|1617|-80.8062|373|35.037115|ROLLS BULK|0.0|14|BULK ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036955555|ROLLS|BAKERY|-80.699686|80.699690085658418|27|2
35.000049|6c2221bdfa19230e50c712703ad0240fe665e5ba|3.0|2015-02-12 16:46:00|80.699698036522989|1||249|35.035225585294562|0|18|1617|-80.8062|373|35.037115|ROLLS BULK|0.0|14|BULK ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036955555|ROLLS|BAKERY|-80.699686|80.699690085658418|27|4
35.000049|7318a1d04202c14792438ca6d05e63d3fdaa2b98|3.0|2014-11-23 18:07:00|80.699698036522989|1||249|35.035225576227809|0|18|1617|-80.64817|373|35.04711|ROLLS BULK|0.0|14|BULK ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036955555|ROLLS|BAKERY|-80.699686|80.699717108215381|129|4
35.000049|9ccbe1b508ebbe188da31415866f09e61b33a018|6.0|2015-02-07 17:38:00|80.699698036522989|1||249|35.035225585294562|0|18|1617|-80.8062|373|35.037115|ROLLS BULK|0.0|14|BULK ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036955555|ROLLS|BAKERY|-80.699686|80.699690085658418|27|8
35.000049|5131da3dc3d72df637db6aa8d8d8f3cc5eb4d11f|2.59|2014-10-26 10:06:00|80.699698036522989|1|7203695298|249|35.035225576584935|0|18|1654|-80.7007|381|35.06858|DESSERT CAKES|0.0|14|OLD FASHION FUDGE CAKE SLICE|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036952981|CAKES|BAKERY|-80.699686|80.699716500181339|273|1
35.000049|2c996199a42fd124b0fa963cc9370a8406bcce53|3.0|2014-11-02 13:15:00|80.699698036522989|1||249|35.035225585294562|0|18|1617|-80.8062|373|35.037115|ROLLS BULK|0.0|14|BULK ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036955555|ROLLS|BAKERY|-80.699686|80.699690085658418|27|4
35.000049|4264d0d3c77c528921f01b0dfffb9e90ec6ab7d0|1.5|2014-10-13 16:51:00|1.4091206135396188|1||249|0.6108660934093487|0|47|1617|-80.699686|373|35.000049|ROLLS BULK|0.0|14|BULK ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00072036955555|ROLLS|BAKERY|-80.699686|1.4084752260255726|249|2
35.000049|0414aed584a84c864a3dd850c53088ac629dcb70|3.0|2014-09-21 15:50:00|1.4091206135396188|1||249|0.6108660934093487|0|47|1617|-80.699686|373|35.000049|ROLLS BULK|0.0|14|BULK ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00072036955555|ROLLS|BAKERY|-80.699686|1.4084752260255726|249|4
35.000049|9312856393fc6be4403f6d62a63250501216a7f5|9.99|2015-01-10 13:38:00|80.699698036522989|1|85877000245|249|35.035225585443811|0|18|458|-80.760919|82|35.024332|CRAFT BEER|0.0|16|OMB CAPT JACK 12OZ 6PACK|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00858770002454|DOMESTIC BEER|BEER|-80.699686|80.699687018251439|343|1
35.000049|54d8e2eb690dbbbce2a0edc9423ca254751dc609|3.99|2014-12-16 16:36:00|80.699698036522989|1|81767001048|249|35.035225585443811|0|18|62|-80.760919|7|35.024332|SPECIALTY BAR/BOX CHOCOLATE|0.0|1|ALTER ECO DARK SEA SALT BAR|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00817670010488|CANDY|G1 GROCERY|-80.699686|80.699687018251439|343|1
35.000049|4026d60ca65dca15b4c8c6a9a8f45752544cbaee|9.99|2015-01-25 15:50:00|80.699698036522989|1|85877000245|249|35.035225585443811|0|18|458|-80.760919|82|35.024332|CRAFT BEER|0.0|16|OMB CAPT JACK 12OZ 6PACK|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00858770002454|DOMESTIC BEER|BEER|-80.699686|80.699687018251439|343|1
35.000049|440577ed40d32fab76ebac6369a68df125e3961f|10.49|2014-09-16 16:41:00|80.699698036522989|1|79849310320|249|35.035225585443811|0|18|36|-80.760919|10|35.024332|PREMIUM GROUND|2.5|1|CARIBOU BLEND  GROUND COFFEE|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00798493103659|COFFEE|G1 GROCERY|-80.699686|80.699687018251439|343|1
35.000049|2a0706fc3335943ad43720d7a983ffcc1337a351|3.69|2015-01-05 16:50:00|1.4091206135396188|1|1410007412|249|0.6108660934093487|0|47|1253|-80.699686|12|35.000049|ALL OTHER COOKIES|0.5|1|PF MILANO MILK CHOCOLATE|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00014100099970|COOKIES|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|9580b68fe8b3be3f98aeb086ccceaf488d0b88ab|2.99|2014-11-16 16:00:00|80.699698036522989|1|1380016610|249|35.035225585443811|0|18|1278|-80.760919|48|35.024332|SINGLE SERVE NUTRITIONAL|0.0|5|LC CAFE CLSSC SESAME CHICKEN|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00013800654557|FROZEN MEALS|FROZEN|-80.699686|80.699687018251439|343|1
35.000049|5a3834470bbe9c4620c5906f1ee61427cefc7693|3.69|2015-02-11 16:21:00|80.699698036522989|1|7518500003|249|35.035225585443811|0|18|1033|-80.760919|163|35.024332|HAMBURGER|0.0|7|MARTIN'S POTATO SANDWICH ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00075185000039|BUNS/ROLLS|COMMERCIAL BAKERY|-80.699686|80.699687018251439|343|1
35.000049|57bca6260c463337dda436249844ddc4ed796a3b|2.89|2015-03-08 16:12:00|80.699698036522989|1|7203695917|249|35.035225585294562|0|18|1625|-80.8062|373|35.037115|FROZEN DOUGH (ROLLS)|0.0|14|FRESH CHICAGO ROLL|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036959171|ROLLS|BAKERY|-80.699686|80.699690085658418|27|1
35.000049|2f1da4eb628a26300957510c631b06d126e06388|2.69|2015-02-25 13:22:00|80.699698036522989|1|7203670627|249|35.035225578015265|0|18|1213|-80.824767|272|35.116751|HISP DINNERS/SHELLS|0.69|1|HT TACO DINNER KIT HARD|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036706270|HISPANIC PREP. FOODS|G1 GROCERY|-80.699686|80.699713932630658|294|1
35.000049|b6441445ea88edc53c4b0fc5a23481279e251572|2.89|2014-12-08 17:14:00|1.4091206135396188|1|7203695917|249|0.6108660934093487|0|47|1625|-80.699686|373|35.000049|FROZEN DOUGH (ROLLS)|0.0|14|FRESH CHICAGO ROLL|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00072036959171|ROLLS|BAKERY|-80.699686|1.4084752260255726|249|1
35.000049|38e03996a3e37154f59f1c8047c6555ac43b58bd|3.69|2015-02-26 16:54:00|80.699698036522989|1|7518500003|249|35.035225585294562|0|18|1033|-80.8062|163|35.037115|HAMBURGER|0.0|7|MARTIN'S POTATO SANDWICH ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00075185000039|BUNS/ROLLS|COMMERCIAL BAKERY|-80.699686|80.699690085658418|27|1
35.000049|ea0a0ae93826142cd2df4e37f349f7888b27b318|3.69|2015-02-21 17:46:00|80.699698036522989|1|7518500003|249|35.035225585443811|0|18|1033|-80.760919|163|35.024332|HAMBURGER|0.0|7|MARTIN'S POTATO SANDWICH ROLLS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00075185000039|BUNS/ROLLS|COMMERCIAL BAKERY|-80.699686|80.699687018251439|343|1
35.000049|6c4fdb913c58933a96e89a2fb6251492d32d4226|10.88|2014-10-23 16:36:00|80.699698036522989|1|20596200000|249|35.035225585443811|0|18|1821|-80.760919|410|35.024332|BH TURKEY|1.98|6|BOARS HEAD MAPLE HONEY TURKEY|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00205962000000|BH MEAT|DELI|-80.699686|80.699687018251439|343|1
35.000049|bdc55f0d825047db65cc1ea3ef445469407a8163|11.21|2015-01-11 15:22:00|80.699698036522989|1|20596200000|249|35.035225585443811|0|18|1821|-80.760919|410|35.024332|BH TURKEY|0.0|6|BOARS HEAD MAPLE HONEY TURKEY|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00205962000000|BH MEAT|DELI|-80.699686|80.699687018251439|343|1
35.000049|ae0da2fb36cf740acc000183e9f8df674aa193b6|10.88|2014-10-27 17:37:00|1.4091206135396188|1|20596200000|249|0.6108660934093487|0|47|1821|-80.699686|410|35.000049|BH TURKEY|1.98|6|BOARS HEAD MAPLE HONEY TURKEY|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00205962000000|BH MEAT|DELI|-80.699686|1.4084752260255726|249|1
35.000049|ba79bacf9b917192c1a70b5d86370302f8978c74|11.21|2014-12-21 17:10:00|80.699698036522989|1|20596200000|249|35.035225585443811|0|18|1821|-80.760919|410|35.024332|BH TURKEY|0.0|6|BOARS HEAD MAPLE HONEY TURKEY|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00205962000000|BH MEAT|DELI|-80.699686|80.699687018251439|343|1
35.000049|e26d0190bc5b67ddd0ae26fb85319cbebd159283|13.3|2014-11-12 15:53:00|80.699698036522989|1|20596200000|249|35.035225585443811|0|18|1821|-80.760919|410|35.024332|BH TURKEY|0.0|6|BOARS HEAD MAPLE HONEY TURKEY|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00205962000000|BH MEAT|DELI|-80.699686|80.699687018251439|343|1
35.000049|aba005255814017b92ebf509b02cf329e0851cfe|10.99|2014-11-25 17:47:00|80.699698036522989|1|20596200000|249|35.035225585443811|0|18|1821|-80.760919|410|35.024332|BH TURKEY|0.0|6|BOARS HEAD MAPLE HONEY TURKEY|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00205962000000|BH MEAT|DELI|-80.699686|80.699687018251439|343|1
35.000049|7b39a4f645a0e69003b8894b6f0de46ea0b9aed9|11.1|2014-12-07 15:31:00|80.699698036522989|1|20596200000|249|35.035225585443811|0|18|1821|-80.760919|410|35.024332|BH TURKEY|0.0|6|BOARS HEAD MAPLE HONEY TURKEY|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00205962000000|BH MEAT|DELI|-80.699686|80.699687018251439|343|1
35.000049|5bc326b6d2d5d59b0303443c209d3c0cef79196e|11.21|2015-01-08 16:21:00|80.699698036522989|1|20596200000|249|35.035225585443811|0|18|1821|-80.760919|410|35.024332|BH TURKEY|0.0|6|BOARS HEAD MAPLE HONEY TURKEY|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00205962000000|BH MEAT|DELI|-80.699686|80.699687018251439|343|1
35.000049|d458ed2ab967cbd30460fa5603dea6979fa4e680|5.93|2014-12-28 15:00:00|80.699698036522989|1|20596200000|249|35.035225585443811|0|18|1821|-80.760919|410|35.024332|BH TURKEY|0.0|6|BOARS HEAD MAPLE HONEY TURKEY|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00205962000000|BH MEAT|DELI|-80.699686|80.699687018251439|343|1
35.000049|baf498e090d0aa8a0949aa035c91c4df8de484f9|11.43|2014-11-20 16:06:00|80.699698036522989|1|20596200000|249|35.035225585443811|0|18|1821|-80.760919|410|35.024332|BH TURKEY|0.0|6|BOARS HEAD MAPLE HONEY TURKEY|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00205962000000|BH MEAT|DELI|-80.699686|80.699687018251439|343|1
35.000049|542ca5ff7a10159a4961caad45d878d763d1e133|9.79|2014-11-06 15:49:00|80.699698036522989|1|20596200000|249|35.035225585294562|0|18|1821|-80.8062|410|35.037115|BH TURKEY|0.0|6|BOARS HEAD MAPLE HONEY TURKEY|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00205962000000|BH MEAT|DELI|-80.699686|80.699690085658418|27|1
35.000049|df8c8da66568bd0ee6dac9d210e88f69eee6c3c2|10.09|2014-10-30 16:51:00|80.699698036522989|1|20596200000|249|35.035225575853595|0|18|1821|-80.758228|410|34.95459|BH TURKEY|0.0|6|BOARS HEAD MAPLE HONEY TURKEY|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00205962000000|BH MEAT|DELI|-80.699686|80.699717732842998|182|1
35.000049|36b08a55063f9c22d1b928d3ae32f57d11cf5c17|11.87|2014-10-09 16:36:00|80.699698036522989|1|20596200000|249|35.035225585443811|0|18|1821|-80.760919|410|35.024332|BH TURKEY|0.0|6|BOARS HEAD MAPLE HONEY TURKEY|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00205962000000|BH MEAT|DELI|-80.699686|80.699687018251439|343|1
35.000049|3226de8931bc9dd9742b5eeefc1d0d540d78e51c|11.21|2015-01-17 15:24:00|80.699698036522989|1|20596200000|249|35.035225576584935|0|18|1821|-80.7007|410|35.06858|BH TURKEY|0.0|6|BOARS HEAD MAPLE HONEY TURKEY|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00205962000000|BH MEAT|DELI|-80.699686|80.699716500181339|273|1
35.000049|b79a3c0b055bda6202c6084d2e7e68ce47ee46d4|10.99|2015-02-10 13:39:00|80.699698036522989|1|20596200000|249|35.035225581038794|0|18|1821|-80.85753|410|35.116638|BH TURKEY|0.0|6|BOARS HEAD MAPLE HONEY TURKEY|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00205962000000|BH MEAT|DELI|-80.699686|80.699707519466116|204|1
35.000049|0a37847744e10fc50f4e742377c8ba73075558f1|10.88|2015-01-04 14:21:00|80.699698036522989|1|20596200000|249|35.035225585443811|0|18|1821|-80.760919|410|35.024332|BH TURKEY|0.0|6|BOARS HEAD MAPLE HONEY TURKEY|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00205962000000|BH MEAT|DELI|-80.699686|80.699687018251439|343|1
35.000049|2ff403fab9d1a2319a8902ec44f2c9a713606289|11.43|2015-01-29 16:09:00|80.699698036522989|1|20596200000|249|35.035225585443811|0|18|1821|-80.760919|410|35.024332|BH TURKEY|0.0|6|BOARS HEAD MAPLE HONEY TURKEY|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00205962000000|BH MEAT|DELI|-80.699686|80.699687018251439|343|1
35.000049|a0f0d419a42cfa91ce8f94fa98261080ebb1f506|10.99|2015-03-01 14:46:00|80.699698036522989|1|20596200000|249|35.035225585443811|0|18|1821|-80.760919|410|35.024332|BH TURKEY|0.0|6|BOARS HEAD MAPLE HONEY TURKEY|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00205962000000|BH MEAT|DELI|-80.699686|80.699687018251439|343|1
35.000049|0cd9c07265b1adb5efb31d1c3e9f30cbe8c6b6a3|3.49|2014-11-01 09:11:00|1.4091206135396188|1|4812127620|249|0.6108660934093487|0|47|1037|-80.699686|164|35.000049|ENGLISH MUFFINS|1.75|7|THOMAS 100% WHEAT ENG MUFN PP|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00048121184070|BREAKFAST|COMMERCIAL BAKERY|-80.699686|1.4084752260255726|249|1
35.000049|6b3e1ad3bd526badc53e81b4e184f9bd80ac9670|4.19|2014-10-12 11:16:00|80.699698036522989|1|4812127620|249|35.035225585443811|0|18|1037|-80.760919|164|35.024332|ENGLISH MUFFINS|2.1|7|THOMAS 100% WHEAT ENG MUFN PP|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00048121184070|BREAKFAST|COMMERCIAL BAKERY|-80.699686|80.699687018251439|343|1
35.000049|f498bc429b993597a5fd7280c7a276bd7330149b|5.29|2014-11-07 18:07:00|1.4091206135396188|1|5150024177|249|0.6108660934093487|0|47|125|-80.699686|19|35.000049|PEANUT BUTTER|1.3|1|JIF CREAMY PEANUT BUTTER|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00051500241776|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|ecde298e94da26a2e32819fa5bdee5df43b62c19|5.29|2014-11-26 17:27:00|80.699698036522989|1|5150024177|249|35.035225585443811|0|18|125|-80.760919|19|35.024332|PEANUT BUTTER|1.3|1|JIF CREAMY PEANUT BUTTER|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00051500241776|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.699686|80.699687018251439|343|1
35.000049|7ac573c9e2e2a6ca7964ed7f46596da8ffbd9b8f|5.29|2014-12-09 15:41:00|80.699698036522989|1|5150024177|249|35.035225585290299|0|18|125|-80.816172|19|35.059823|PEANUT BUTTER|1.3|1|JIF CREAMY PEANUT BUTTER|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00051500241776|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.699686|80.699690139960765|66|1
35.000049|66676a7191facb80a482faf12620c03d52d62a97|1.99|2014-12-30 17:13:00|80.699698036522989|1|7127923100|249|35.035225585443811|0|18|555|-80.760919|64|35.024332|PACKAGED SALADS|0.0|4|F.E. BABY SPRING SALAD MIX|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00071279231006|FRESH PRODUCE|PRODUCE|-80.699686|80.699687018251439|343|1
35.000049|1965942035487bafb9bff49ee4a8608671766cb8|1.99|2014-11-21 18:10:00|1.4091206135396188|1|7127923100|249|0.6108660934093487|0|47|555|-80.699686|64|35.000049|PACKAGED SALADS|0.0|4|F.E. BABY SPRING SALAD MIX|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00071279231006|FRESH PRODUCE|PRODUCE|-80.699686|1.4084752260255726|249|1
35.000049|72600a2540dcbc432cd50f96be979c5ae0ea5743|1.99|2015-01-19 11:52:00|1.4091206135396188|1|7127923100|249|0.6108660934093487|0|47|555|-80.699686|64|35.000049|PACKAGED SALADS|0.0|4|F.E. BABY SPRING SALAD MIX|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00071279231006|FRESH PRODUCE|PRODUCE|-80.699686|1.4084752260255726|249|1
35.000049|d21f46a57c8b4b88d35768edaa67556947ad920b|2.79|2014-10-06 16:06:00|80.699698036522989|1|7020059601|249|35.035225585443811|0|18|22|-80.760919|28|35.024332|CROUTONS|1.0|1|TEXAS TORT STRIP CHILI LIME|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00070200596009|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.699686|80.699687018251439|343|1
35.000049|d25ca1d66bcad7db975f27f4b07ed4555002fa83|4.99|2015-01-12 13:25:00|1.4091206135396188|1|7203688077|249|0.6108660934093487|0|47|523|-80.699686|64|35.000049|FRESH POTATOES|1.5|4|HT RED POTATO 5LB BAG|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00072036880772|FRESH PRODUCE|PRODUCE|-80.699686|1.4084752260255726|249|1
35.000049|14753148825ac486721cb581a029486a5167fb54|5.99|2014-12-20 07:32:00|1.4091206135396188|1|7203688215|249|0.6108660934093487|0|47|500|-80.699686|64|35.000049|FRESH APPLES|0.0|4|HT GALA APPLE 5LB|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00072036882158|FRESH PRODUCE|PRODUCE|-80.699686|1.4084752260255726|249|1
35.000049|92d6d23a843eb016f3d2e4726c45f33438468cf3|4.99|2014-12-18 16:43:00|1.4091206135396188|1|7203688077|249|0.6108660934093487|0|47|523|-80.699686|64|35.000049|FRESH POTATOES|0.0|4|HT RED POTATO 5LB BAG|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00072036880772|FRESH PRODUCE|PRODUCE|-80.699686|1.4084752260255726|249|1
35.000049|19aaa7f51379aec508087f3375a2f9d27f906725|3.99|2015-02-26 16:17:00|1.4091206135396188|1|7203688077|249|0.6108660934093487|0|47|523|-80.699686|64|35.000049|FRESH POTATOES|0.0|4|HT RED POTATO 5LB BAG|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00072036880772|FRESH PRODUCE|PRODUCE|-80.699686|1.4084752260255726|249|1
35.000049|2f323870ce704f8026d4cec330fe7e9ca83cf077|17.98|2015-02-23 13:59:00|1.4091206135396188|1|7203697794|249|0.6108660934093487|0|47|6903|-80.699686|1582|35.000049|DOG RAWHIDE CHEW|6.0|18|YP 1LB WHITE CHIPS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00072036977946|PET NEEDS|GM|-80.699686|1.4084752260255726|249|2
35.000049|919e55a0f25956f244934cb603fcabb468464c94|0.79|2014-11-18 16:11:00|80.699698036522989|1||249|35.035225585443811|0|18|532|-80.760919|64|35.024332|FRESH CUCUMBERS|0.0|4|COO CUCUMBERS S/S|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00204062000002|FRESH PRODUCE|PRODUCE|-80.699686|80.699687018251439|343|1
35.000049|b348f174810b583837fd139d5b3a2c1a450fc3ad|2.49|2014-09-22 16:26:00|80.699698036522989|1||249|35.035225585294562|0|18|544|-80.8062|64|35.037115|FRESH PRODUCE FRSH HERBS|0.0|4|BUNCHED ARUGULA (RPC)|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00204884000006|FRESH PRODUCE|PRODUCE|-80.699686|80.699690085658418|27|1
35.000049|e0a4c87103b51e67b1d2199d30afc718c783ee54|1.29|2014-12-24 17:00:00|1.4091206135396188|1|7203657030|249|0.6108660934093487|0|47|322|-80.699686|53|35.000049|SOUR CREAM|0.0|3|HT LIGHT SOUR CREAM|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00072036600349|CULTURES|DAIRY|-80.699686|1.4084752260255726|249|1
35.000049|0836b6d938fe919a122ab156eb4a590f8a8bc032|4.99|2014-09-10 15:47:00|80.699698036522989|1|4242101480|249|35.035225585443811|0|18|482|-80.760919|100|35.024332|PRECOOKED BACON|0.7|19|BOARS HEAD FULLY COOKED BACON|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00042421014808|BACON|CASE READY MEATS|-80.699686|80.699687018251439|343|1
35.000049|6d3892588f27516930dece8dceee756b9a68a456|8.79|2014-09-20 12:19:00|80.699698036522989|1||249|35.035225585443811|0|18|503|-80.760919|64|35.024332|FRESH GRAPES|5.33|4|GREEN GRAPES, SEEDLESS 12/16|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00204022000004|FRESH PRODUCE|PRODUCE|-80.699686|80.699687018251439|343|1
35.000049|7ad3e43d812c4392d1f39d7ab66e264a51033c88|7.59|2014-09-25 15:50:00|80.699698036522989|1|4667716908|249|35.035225585443811|0|18|6140|-80.760919|1546|35.024332|BULB-CLEAR|0.0|18|DURAMAX VANITY CLEAR 40W|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00046677169084|LIGHT BULBS/ELECTRICAL|GM|-80.699686|80.699687018251439|343|1
35.000049|2af0f38cdbeb2fa97ece9c8150a2c2bb70281678|6.49|2015-02-01 11:28:00|1.4091206135396188|1|4698501674|249|0.6108660934093487|0|47|4237|-80.699686|1200|35.000049|MEDICATED LIP CARE|0.0|17|LYSINE+LIPCLEAR CLD SR TRTMNT|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00046985016742|COUGH/COLD/SINUS|HBC|-80.699686|1.4084752260255726|249|1
35.000049|9fc578116a3a52e1868144232f0309cf0b6fab8a|16.99|2014-12-29 16:11:00|80.699698036522989|1|7203698131|249|35.035225575853595|0|18|6903|-80.758228|1582|34.95459|DOG RAWHIDE CHEW|0.0|18|YP 2LB NATURAL CHIPS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036981318|PET NEEDS|GM|-80.699686|80.699717732842998|182|1
35.000049|201dcefb3a1e0484256e86b3b3c388fc2d768c41|2.49|2014-12-24 13:36:00|80.699698036522989|1|7203688130|249|35.035225585443811|0|18|556|-80.760919|64|35.024332|PACKAGED VEGETABLES|0.0|4|HT DICED ROMA TOMATOES|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036881328|FRESH PRODUCE|PRODUCE|-80.699686|80.699687018251439|343|1
35.000049|5280dd7da52c668beb1bd6a51b23a1319e1d0c13|8.5|2014-10-15 16:50:00|80.699698036522989|1|4400000488|249|35.035225576584935|0|18|89|-80.7007|12|35.06858|GRAHAM CRACKERS|1.5|1|HONEYMAID GRAHAMS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00044000004637|COOKIES|G1 GROCERY|-80.699686|80.699716500181339|273|2
35.000049|0260e10efc7a4ee1d9e243e64644f74c836e37c1|2.0|2014-12-19 18:41:00|80.699698036522989|1|4000000435|249|35.035225575853595|0|18|47|-80.758228|7|34.95459|REGISTER BARS|0.2|1|(FE)TWIX CARAMEL COOKIE BAR|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00040000004356|CANDY|G1 GROCERY|-80.699686|80.699717732842998|182|2
35.000049|075960461af30d66f7b8ee7e629fc2f46e4d0f66|1.49|2015-01-07 16:15:00|80.699698036522989|1|7203653022|249|35.035225575853595|0|18|1273|-80.758228|50|34.95459|BAG VEG NON STEAM|0.49|5|HT CUT OKRA|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036537522|VEGETABLES-FROZEN|FROZEN|-80.699686|80.699717732842998|182|1
35.000049|dff8d8115bf76d870f0fc34503aa15dad0ba85fe|2.69|2015-02-19 17:22:00|80.699698036522989|1|1380016610|249|35.035225585443811|0|18|1271|-80.760919|41|35.024332|PROTEIN BREAKFAST|0.0|5|LEAN CUIS TKY SAUS EGG SCRAM|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00013800872326|BREAKFAST FOODS FROZEN|FROZEN|-80.699686|80.699687018251439|343|1
35.000049|17a40f3977149c550e2fc00d4027d87a2770c318|3.98|2014-09-11 15:59:00|80.699698036522989|1|7203688096|249|35.035225585290299|0|18|526|-80.816172|64|35.059823|FRESH MUSHROOMS|0.4|4|HT SLICED WHITE MUSHROOMS|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036880963|FRESH PRODUCE|PRODUCE|-80.699686|80.699690139960765|66|2
35.000049|d44905de1b28fb7134122f097adb1b3b38345d64|8.99|2014-10-10 17:59:00|1.4091206135396188|1|8769230050|249|0.6108660934093487|0|47|458|-80.699686|82|35.000049|CRAFT BEER|0.0|16|SAM ADAMS SEASONAL 6PK|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00087692300502|DOMESTIC BEER|BEER|-80.699686|1.4084752260255726|249|1
35.000049|c5221f34cf9d8c39f79ea9d6c68184e52a0a3f2d|1.49|2014-12-22 11:39:00|80.699698036522989|1|3084900006|249|35.035225585443811|0|18|577|-80.760919|136|35.024332|OTHER MERCH FR MSC JUICE|0.0|4|SICILIA LIME JUICE 4OZ|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00030849000060|OTHER MERCHANDISE|PRODUCE|-80.699686|80.699687018251439|343|1
35.000049|c4b367b4690edd993a05bca1054091529935d67d|3.29|2014-12-16 12:47:00|80.699698036522989|1|1410008786|249|35.035225578015265|0|18|1033|-80.824767|163|35.116751|HAMBURGER|0.0|7|PEP GOLDEN POTATO HAMS PP|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00014100091417|BUNS/ROLLS|COMMERCIAL BAKERY|-80.699686|80.699713932630658|294|1
35.000049|c566f9d6819a45c6fa8fe972aba5bce7ea0f6e96|4.59|2015-02-19 17:30:00|1.4091206135396188|1|67811225415|249|0.6108660934093487|0|47|4928|-80.699686|1245|35.000049|EYE-ARTIFICAL TEARS|1.0|17|CLEAR EYES DROPS MAX RELIEF|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00678112665778|EYE & EAR CARE|HBC|-80.699686|1.4084752260255726|249|1
35.000049|ecdb8d381c4a9c38d8a4a57634c09bf2843ad650|5.25|2014-10-03 17:53:00|80.699698036522989|1|7203633086|249|35.035225585443811|0|18|1148|-80.760919|21|35.024332|ALMONDS|1.75|1|HT ROASTED ALMONDS LIGHT SALT|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00072036979537|NUTS|G1 GROCERY|-80.699686|80.699687018251439|343|1
35.000049|8b7219eeaa5eca6154993c1cba91ef49ed5e9de4|5.25|2014-12-15 17:18:00|1.4091206135396188|1|7203633086|249|0.6108660934093487|0|47|1148|-80.699686|21|35.000049|ALMONDS|1.75|1|HT ROASTED ALMONDS LIGHT SALT|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00072036979537|NUTS|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|19d505118463ab3bea984018866bf1181699832a|2.29|2015-02-28 19:35:00|1.4091206135396188|1|7046203598|249|0.6108660934093487|0|47|50|-80.699686|7|35.000049|PEG CANDY|0.29|1|SOUR PATCH KIDS EXPLODERZ|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00070462433517|CANDY|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|5fd4564f2e3a6b19da648bf661b09cbefb8a382a|3.99|2014-09-20 12:21:00|80.699698036522989|1|7127927100|249|35.035225585443811|0|18|555|-80.760919|64|35.024332|PACKAGED SALADS|0.99|4|F.E. BABY SPINACH|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00071279271002|FRESH PRODUCE|PRODUCE|-80.699686|80.699687018251439|343|1
35.000049|5bc99a1418410a4d53c48cf07b8d0a3612ea1360|1.19|2015-01-08 15:17:00|80.699698036522989|1|4000000419|249|35.035225575853595|0|18|727|-80.758228|7|34.95459|SEASONAL CANDY-SINGLE FAC|0.6|1|I/O(C14)TWIX PEANUT BUTTER BAR|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|35.030887098939942|00040000004196|CANDY|G1 GROCERY|-80.699686|80.699717732842998|182|1
35.000049|76ef76a12e3e334f95b6461d9974aff84abd6624|1.79|2014-11-29 16:43:00|1.4091206135396188|1|7203620122|249|0.6108660934093487|0|47|139|-80.699686|20|35.000049|REMAINING SHELF STABLE JUICES|0.0|1|HT LEMON JUICE|a6fe77a48a3764d8616b0eae8ab9bf50a23d31e3|2.430617106437779|0.61242566243833529|00072036201225|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.43259|2a65f394968c476d6737e3ac78200203070b64a0|5.49|2015-01-19 11:42:00|1.4057311447477159|4|2301290134|202|0.6184153580092175|0|52|1477|-80.605588|485|35.43259|SUSHI HYBRID|0.0|6|VEGETABLE COMBO SP|a8929b5735c3eaa61fa457b4fcbfdf9fd7f63cc9|3.332402133592992|0.6209993146566879|00023012901349|SUSHI|DELI|-80.605588|1.406832906106031|202|1
35.124987|d5f20caf1a68555e2b496bd45f10cec30d8c0024|7.19|2014-12-20 08:30:00|80.7095026033777|4|3760048620|157|35.157870607009791|0|51|358|-80.654118|100|35.123768|REGULAR BACON|0.0|19|HORMEL BLACK LABEL LOW SALT|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00037600486200|BACON|CASE READY MEATS|-80.709466|80.709475587267946|473|1
35.124987|ec5ca237731024e3316c71cc75ca52bfa7c2909d|2.0|2014-12-23 17:51:00|80.7095026033777|4||157|35.157870607009791|0|51|512|-80.654118|64|35.123768|FRSH PROD FRSH FRUIT REM|0.0|4|MANGOS|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00204959000009|FRESH PRODUCE|PRODUCE|-80.709466|80.709475587267946|473|2
35.124987|8ff6c3fd550eca14bb44dcc1c9c164d5e078fb5a|6.0|2014-10-04 14:02:00|80.7095026033777|4||157|35.157870607009791|0|51|512|-80.654118|64|35.123768|FRSH PROD FRSH FRUIT REM|0.0|4|MANGOS|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00204959000009|FRESH PRODUCE|PRODUCE|-80.709466|80.709475587267946|473|6
35.124987|5a9e0035e08f8e3d0d28e087ac0f2f72a16fcfea|3.0|2014-10-12 19:23:00|80.7095026033777|4||157|35.157870607009791|0|51|512|-80.654118|64|35.123768|FRSH PROD FRSH FRUIT REM|0.0|4|MANGOS|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00204959000009|FRESH PRODUCE|PRODUCE|-80.709466|80.709475587267946|473|3
35.124987|49eeaaa288586a404350e59efcef73d6f932d9f6|2.0|2014-09-30 14:41:00|80.7095026033777|4||157|35.157870607009791|0|51|512|-80.654118|64|35.123768|FRSH PROD FRSH FRUIT REM|0.0|4|MANGOS|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00204959000009|FRESH PRODUCE|PRODUCE|-80.709466|80.709475587267946|473|2
35.124987|42573ea0d83a50e03b8035f1bf9fda2db5d21be0|1.34|2015-01-01 11:05:00|80.7095026033777|4|7203660058|157|35.157870607009791|0|51|325|-80.654118|54|35.123768|BISCUITS-REFRIGERATED|0.0|3|HT TEXAS STYLE BUTTERMILK BIS|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00072036600608|DOUGH PRODUCTS|DAIRY|-80.709466|80.709475587267946|473|1
35.124987|3b0c955ee763722e435452f3abc73c21e109dd47|14.99|2014-11-26 20:47:00|80.7095026033777|4|8834510053|157|35.157870607009791|0|51|459|-80.654118|83|35.123768|IMPORT BEER|0.0|16|NEWCASTLE 12PK 12OZ BTL|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00088345100531|IMPORT BEER|BEER|-80.709466|80.709475587267946|473|1
35.124987|e35ca2439008dce27bdc9d4c90f7a6f7f5b1873a|3.5|2014-11-08 19:40:00|80.7095026033777|4|7203698425|157|35.157870607009791|0|51|254|-80.654118|892|35.123768|PREMIUM PIZZA|0.5|5|HT THIN CRUST PEPP/SAUS PIZZA|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00072036984265|FROZEN PIZZA|FROZEN|-80.709466|80.709475587267946|473|1
35.124987|b937a382779c4967640e35ba6bd9af539c5616dd|7.16|2014-11-26 20:50:00|80.7095026033777|4|8079380770|157|35.157870607009791|0|51|99|-80.654118|32|35.123768|LIQUID TEA|2.16|1|D FUZE SLENDERIZE PEACH MANGO|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00080793807826|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.709466|80.709475587267946|473|4
35.124987|c5ffce95fe7c61a736cfc8353386625ca6036af0|4.98|2015-01-10 11:38:00|80.7095026033777|4|70935100016|157|35.157870607009791|0|51|556|-80.654118|64|35.123768|PACKAGED VEGETABLES|0.0|4|APIO BROCCOLI COLE SLAW|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00709351000164|FRESH PRODUCE|PRODUCE|-80.709466|80.709475587267946|473|2
35.124987|b1950c01ec5ab6bbd753b4698a252844e67a4965|1.19|2014-11-20 12:20:00|80.7095026033777|4|7247001725|157|35.157870607009791|0|51|1641|-80.654118|377|35.123768|PACKAGED DONUTS|0.0|14|KK GLAZED FRUIT PIE- APPLE PP|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00072470017253|DONUTS|BAKERY|-80.709466|80.709475587267946|473|1
35.124987|727fe070ae6687a9b65a6d31821a2880eb1fad25|0.5|2014-10-27 19:53:00|80.7095026033777|4||157|35.157870607009791|0|51|543|-80.654118|64|35.123768|FRESH GARLIC|0.0|4|COO GARLIC, WHITE, BULK|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00204608000008|FRESH PRODUCE|PRODUCE|-80.709466|80.709475587267946|473|1
35.124987|e6730371fc04025bfa6831f56a16aecd259c9f4a|3.29|2014-12-29 16:39:00|80.7095026033777|4|4144930140|157|35.157870607009791|0|51|9|-80.654118|2|35.123768|DESSERT MIXES|0.3|1|KRUSTEAZ CINN. CRUMB CAKE MIX|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00041449111407|BAKING MIXES|G1 GROCERY|-80.709466|80.709475587267946|473|1
35.124987|dad92749115963fdda2bdb6def3bee28a72f7c63|3.19|2014-10-19 10:18:00|80.7095026033777|4|3760019991|157|35.157870607009791|0|51|175|-80.654118|27|35.123768|CANNED MEATS|1.52|1|HORMEL MAR KTC ROAST BEEF HASH|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00037600199919|PREPARED FOODS-RTS|G1 GROCERY|-80.709466|80.709475587267946|473|1
35.124987|d5658336ba28959155b31407ccb7c383bfcb1dbf|1.4|2014-11-22 16:46:00|80.7095026033777|4||157|35.157870607009791|0|51|502|-80.654118|64|35.123768|FRESH BANANAS|0.0|4|BANANAS, YELLOW|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00204011000008|FRESH PRODUCE|PRODUCE|-80.709466|80.709475587267946|473|1
35.124987|1d4e909f2cb7042f3bff19e5d1167c0904c026dc|4.49|2014-12-19 19:15:00|80.7095026033777|4|70897111893|157|35.157870601314983|0|51|1703|-80.78468|387|35.096737|SEASONAL COOKIES|1.5|14|HOLIDAY WHT FRSTD SUGAR COOKIE|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00708971118938|COOKIES|BAKERY|-80.709466|80.709491534591407|30|1
35.124987|d679276f77cc5002465816490620ad3b4589e9a4|2.58|2014-09-14 17:07:00|80.7095026033777|4|8379152001|157|35.157870603736932|0|51|1981|-80.70901|480|35.17335|CHIPS|0.0|6|CALIFORNIA SEA SALT CHIPS|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00705845015201|DRY GOODS|DELI|-80.709466|80.709486342334188|174|2
35.124987|e52c34dbfa24b21dd3a969c97efd136653ddda53|9.38|2014-09-13 20:02:00|80.7095026033777|4|7347200123|157|35.157870607009791|0|51|1462|-80.654118|40|35.123768|FROZEN GLUTEN FREE BREAD|0.0|5|EZEKIEL 4:9 SPROUTED GRAIN ORG|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00073472001202|FROZEN DOUGH|FROZEN|-80.709466|80.709475587267946|473|2
35.124987|ee11d6af6666c22ce3ad4c89503a8ffe18214e67|9.38|2014-11-16 16:39:00|80.7095026033777|4|7347200123|157|35.157870607009791|0|51|1462|-80.654118|40|35.123768|FROZEN GLUTEN FREE BREAD|0.0|5|EZEKIEL 4:9 SPROUTED GRAIN ORG|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00073472001202|FROZEN DOUGH|FROZEN|-80.709466|80.709475587267946|473|2
35.124987|2683a19cf6e17fc2b4777ccf5b3a961546467420|12.99|2015-02-01 17:06:00|1.4091206135396188|4|1820005990|157|0.6130466728702054|0|47|456|-80.709466|82|35.124987|DOMESTIC SUPER PREM 12PK&>|0.0|16|MICHELOB ULTRA 12PK 12OZ BTL|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|0.61242566243833529|00018200059902|DOMESTIC BEER|BEER|-80.709466|1.4086459192264178|157|1
35.124987|48d68c61f21b4e8192d37ca01167b81f710be5a7|12.5|2015-02-04 12:11:00|80.7095026033777|4|7218063979|157|35.157870607009791|0|51|284|-80.654118|892|35.123768|SUPER PREMIUM PIZZA|2.5|5|FRESCHETTA 12 PEPPERONI PIZZA|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00072180639790|FROZEN PIZZA|FROZEN|-80.709466|80.709475587267946|473|2
35.124987|ad6691545080a6ff96ae2fe95e618d5bc7c71252|7.0|2014-09-24 14:44:00|80.7095026033777|4|7203698425|157|35.157870607009791|0|51|254|-80.654118|892|35.123768|PREMIUM PIZZA|1.0|5|HT THIN CRUST PEPPERONI PIZZA|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00072036984241|FROZEN PIZZA|FROZEN|-80.709466|80.709475587267946|473|2
35.124987|976c973356821e147365a1052da607aef3a8a21b|4.29|2014-10-18 20:27:00|80.7095026033777|4|5100007519|157|35.157870607009791|0|51|270|-80.654118|307|35.123768|DESSERTS FROZEN|0.0|5|PEP FARM APPLE TURNOVER|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00051000075017|DESSERTS FROZEN|FROZEN|-80.709466|80.709475587267946|473|1
35.124987|c18fe0bf741f189300cc818b1d420b90e95b15db|4.29|2014-09-13 00:01:00|1.4091206135396188|4|5100007519|157|0.6130466728702054|0|47|270|-80.709466|307|35.124987|DESSERTS FROZEN|0.0|5|PEP FARM APPLE TURNOVER|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|0.61242566243833529|00051000075017|DESSERTS FROZEN|FROZEN|-80.709466|1.4086459192264178|157|1
35.124987|513f01d9b12f20bce6b791e6a17a38e09b25800f|6.79|2014-12-16 08:42:00|1.4091206135396188|4|4850001833|157|0.6130466728702054|0|47|335|-80.709466|56|35.124987|ORANGE JUICE-REGRIGERATED|0.8|3|TROPICANA CALCIUM ORANGE JUICE|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|0.61242566243833529|00048500018309|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.709466|1.4086459192264178|157|1
35.124987|82eecb64eb7797913489758039595e1ff6c5d405|4.65|2015-01-29 19:21:00|80.7095026033777|4|7218063473|157|35.157870607009791|0|51|254|-80.654118|892|35.123768|PREMIUM PIZZA|1.31|5|RED BARON THN CRUST PEPPERONI|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00072180633224|FROZEN PIZZA|FROZEN|-80.709466|80.709475587267946|473|1
35.124987|030a829ab81368722c915792d21b69eaabc23ba8|4.65|2015-01-09 13:59:00|80.7095026033777|4|7218063473|157|35.157870607009791|0|51|254|-80.654118|892|35.123768|PREMIUM PIZZA|0.0|5|RED BARON THN CRUST PEPPERONI|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00072180633224|FROZEN PIZZA|FROZEN|-80.709466|80.709475587267946|473|1
35.124987|28907c4169b40bda4ca2841643a32dadc8ee382c|2.19|2015-01-03 12:13:00|80.7095026033777|4|2900001546|157|35.157870607009791|0|51|1244|-80.654118|21|35.123768|OTHER NUTS|0.0|1|PLANTERS SUNFLOWER KERNEL|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00029000015463|NUTS|G1 GROCERY|-80.709466|80.709475587267946|473|1
35.124987|9d775f3790627875eaa04bfb9eb5a0ff431045a1|1.69|2015-02-01 10:11:00|80.7095026033777|4|4900000044|157|35.157870607009791|0|51|54|-80.654118|8|35.123768|DIET|0.0|23|CB DIET COKE CONTOUR 20 OZ NR|b067a9094f24513fb682e3e5e70348f0b4c25456|2.272177897884649|35.154129163572591|00049000000450|CARBONATED BEVERAGES|BEVERAGE|-80.709466|80.709475587267946|473|1
35.444064|24478e99c057f38d7fe7af24a896b97b393ffc5c|10.99|2014-09-17 16:32:00|1.4102725052409182|4|7203663048|121|0.6186156170875914|0|1|297|-80.995484|49|35.444064|GROUND BEEF|0.0|2|93% LEAN GROUND BEEF 2 LB|b1b1b77bb6ceb4d7f9f7b622cb35bbcf22d04f3c|1.5825730080851959|0.61833652052202714|00072036630483|BEEF|MEAT|-80.995484|1.413637875046387|121|1
35.444064|4be5c27c40f4ae11c40d545632f2511bdd720e08|4.59|2014-09-14 15:05:00|1.4102725052409182|4|7203663117|121|0.6186156170875914|0|1|1262|-80.995484|57|35.444064|HALF N HALF WHIPPING CREAM|0.0|3|HT HALF & HALF|b1b1b77bb6ceb4d7f9f7b622cb35bbcf22d04f3c|1.5825730080851959|0.61833652052202714|00072036631176|MILK|DAIRY|-80.995484|1.413637875046387|121|1
35.444064|30f67c85fa36c03b9baf3b78bdd1b6b54097e7d5|31.98|2015-01-30 16:50:00|1.4102725052409182|4|20220200000|121|0.6186156170875914|0|1|299|-80.995484|49|35.444064|ANGUS BEEF|8.0|2|ANGUS BEEF FILET MIGNON CUSTOM|b1b1b77bb6ceb4d7f9f7b622cb35bbcf22d04f3c|1.5825730080851959|0.61833652052202714|00202209000007|BEEF|MEAT|-80.995484|1.413637875046387|121|1
35.444064|19bb79edfe3b4f6bc7e66d4df1193b58f041b2cd|17.97|2014-10-11 12:37:00|1.4102725052409182|4|1834175101|121|0.6186156170875914|0|1|9935|-80.995484|885|35.444064|NFS POP CAB SAUV|2.02|13|BAREFOOT CAB SAUV|b1b1b77bb6ceb4d7f9f7b622cb35bbcf22d04f3c|1.5825730080851959|0.61833652052202714|00018341751017|POPULAR (4-$7.99)|WINE|-80.995484|1.413637875046387|121|3
35.444064|ebd17190b1f9fa3797ebf1c3660b64d863db3e40|9.38|2015-01-21 16:20:00|1.4102725052409182|4|71514111357|121|0.6186156170875914|0|1|330|-80.995484|55|35.444064|EGGS|1.19|3|EGGLAND BEST 18 GRADE A LARGE|b1b1b77bb6ceb4d7f9f7b622cb35bbcf22d04f3c|1.5825730080851959|0.61833652052202714|00715141113570|EGGS FRESH|DAIRY|-80.995484|1.413637875046387|121|2
35.444064|12d52e960d4a995fa7b4b667b2b12a4b269c1677|1.38|2014-10-13 16:34:00|1.4102725052409182|4||121|0.6186156170875914|0|1|523|-80.995484|64|35.444064|FRESH POTATOES|0.0|4|"COO RED POTATO ""A""SIZE, BULK"|b1b1b77bb6ceb4d7f9f7b622cb35bbcf22d04f3c|1.5825730080851959|0.61833652052202714|00204073000008|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|c5840ff2d2f6f85e52b9483fc6f65b589894e8a4|2.49|2014-11-02 11:32:00|1.4102725052409182|4|7878351001|121|0.6186156170875914|0|1|527|-80.995484|64|35.444064|FRESH CARROTS|0.0|4|CARROT CHIPS, PKG|b1b1b77bb6ceb4d7f9f7b622cb35bbcf22d04f3c|1.5825730080851959|0.61833652052202714|00078783510016|FRESH PRODUCE|PRODUCE|-80.995484|1.413637875046387|121|1
35.444064|56dd96985fc7b64a36bc9fdedf48f40e50ea3881|7.78|2014-11-15 11:02:00|1.4102725052409182|4|2100012277|121|0.6186156170875914|0|1|320|-80.995484|53|35.444064|COTTAGE CHEESE|1.78|3|BREAKSTONE 2% COTTAGE CHEESE|b1b1b77bb6ceb4d7f9f7b622cb35bbcf22d04f3c|1.5825730080851959|0.61833652052202714|00021000123544|CULTURES|DAIRY|-80.995484|1.413637875046387|121|2
35.444064|c03c780ce905b850805d7ca42124a13f8694d116|5.98|2014-09-18 16:35:00|1.4102725052409182|4|2484201121|121|0.6186156170875914|0|1|1887|-80.995484|440|35.444064|PASTA CUTS|0.0|6|BUITONI FETTUCINE|b1b1b77bb6ceb4d7f9f7b622cb35bbcf22d04f3c|1.5825730080851959|0.61833652052202714|00024842011215|PASTA|DELI|-80.995484|1.413637875046387|121|2
35.444064|3ee775def1c00133e3151b2719e27c282bc647f3|6.99|2014-11-24 17:01:00|1.4102725052409182|4|3114200011|121|0.6186156170875914|0|1|2021|-80.995484|505|35.444064|FRESH CHEESE|0.0|6|BELGIOIOSO MASCARPONE|b1b1b77bb6ceb4d7f9f7b622cb35bbcf22d04f3c|1.5825730080851959|0.61833652052202714|00031142000115|SPECIALTY CHEESE|DELI|-80.995484|1.413637875046387|121|1
35.444064|5db85d3731a059e75c5e51e9ff0a6120fc39d8cf|3.99|2014-11-01 16:48:00|1.4102725052409182|4|7835470843|121|0.6186156170875914|0|1|317|-80.995484|52|35.444064|CHUNK AND BAR CHEESE|1.49|3|CABOT 75% LIGHT WHITE CHEDDAR|b1b1b77bb6ceb4d7f9f7b622cb35bbcf22d04f3c|1.5825730080851959|0.61833652052202714|00078354707272|CHEESE|DAIRY|-80.995484|1.413637875046387|121|1
35.053394|2805f3107c7165523ff8b8ddba676fdd4dc172a1|6.29|2014-12-05 16:54:00|80.848351720559364|4|4369507143|11|35.091845859777088|0|25|1276|-80.847383|279|35.024464|FROZEN SANDWICHES|1.3|5|HOT POCKETS 5PK PEPP PIZZA|b43e43bd71d22e54b77bb1759ac94f3e2dda3d9f|2.656930769193146|35.082633588753836|00043695071436|FROZEN SANDWICH AND SNACKS|FROZEN|-80.848528|80.848541914011989|317|1
35.053394|b72ad982f0fcbcd6c989276838be3945ad7deec7|1.0|2014-10-08 16:26:00|80.848351720559364|4|812|11|35.091845859777088|0|25|1639|-80.847383|377|35.024464|BULK (DONUTS)|0.5|14|NEW BULK DONUT CODE|b43e43bd71d22e54b77bb1759ac94f3e2dda3d9f|2.656930769193146|35.082633588753836|00000000008120|DONUTS|BAKERY|-80.848528|80.848541914011989|317|1
35.053394|cc585a105e7c8f7ef07d076b8fdefd506353be40|2.0|2015-01-05 16:31:00|80.848351720559364|4|812|11|35.091845859777088|0|25|1639|-80.847383|377|35.024464|BULK (DONUTS)|0.0|14|NEW BULK DONUT CODE|b43e43bd71d22e54b77bb1759ac94f3e2dda3d9f|2.656930769193146|35.082633588753836|00000000008120|DONUTS|BAKERY|-80.848528|80.848541914011989|317|2
35.053394|2b3e3c662ee353fa79463a53a0804ec4da092f88|2.99|2014-12-31 18:12:00|80.848351720559364|4|7433610102|11|35.091845859777088|0|25|342|-80.847383|57|35.024464|FRESH MILK|0.0|3|HIGHLAND CREST WHOLE MILK|b43e43bd71d22e54b77bb1759ac94f3e2dda3d9f|2.656930769193146|35.082633588753836|00074336879203|MILK|DAIRY|-80.848528|80.848541914011989|317|1
35.053394|be7f554a52dfd2fc4610cbee1e45ed4aeee7b5c8|3.75|2014-09-14 14:32:00|80.848351720559364|4|7433610102|11|35.091845859777088|0|25|342|-80.847383|57|35.024464|FRESH MILK|0.0|3|HIGHLAND CREST WHOLE MILK|b43e43bd71d22e54b77bb1759ac94f3e2dda3d9f|2.656930769193146|35.082633588753836|00074336879203|MILK|DAIRY|-80.848528|80.848541914011989|317|1
35.053394|1afd5fb60bb264523742e6898f78c9ef3c2fd191|1.97|2014-11-09 11:21:00|80.848351720559364|4|7203642077|11|35.091845859777088|0|25|236|-80.847383|38|35.024464|DRY BEANS|0.0|1|HT PEAS DRY BLACKEYE|b43e43bd71d22e54b77bb1759ac94f3e2dda3d9f|2.656930769193146|35.082633588753836|00072036429964|RICE GRAINS AND BEANS|G1 GROCERY|-80.848528|80.848541914011989|317|1
35.053394|52ce4ccb1dafb2254f03f11a9b99fc94f1270a43|1.79|2014-12-31 12:22:00|80.848351720559364|4|7203663158|11|35.091845859777088|0|25|495|-80.847383|108|35.024464|NON REFRIGERATED|0.8|19|HT CORN TORTILLA 30CT|b43e43bd71d22e54b77bb1759ac94f3e2dda3d9f|2.656930769193146|35.082633588753836|00072036631589|TORTILLAS|CASE READY MEATS|-80.848528|80.848541914011989|317|1
35.053394|75e7ea63c96990e733147a8817b22fcd86e47889|2.29|2014-11-08 17:39:00|80.848351720559364|4|7800023046|11|35.091845859777088|0|25|55|-80.847383|8|35.024464|REGULAR|1.29|23|CANADA DRY CBRY G/ALE 2LTR|b43e43bd71d22e54b77bb1759ac94f3e2dda3d9f|2.656930769193146|35.082633588753836|00078000156461|CARBONATED BEVERAGES|BEVERAGE|-80.848528|80.848541914011989|317|1
35.053394|e6b85ea2f3131b2bfaa655c508cc2d51265ce52a|1.77|2014-11-07 16:05:00|80.848351720559364|4|7203657031|11|35.091845859777088|0|25|322|-80.847383|53|35.024464|SOUR CREAM|0.52|3|HT SOUR CREAM|b43e43bd71d22e54b77bb1759ac94f3e2dda3d9f|2.656930769193146|35.082633588753836|00072036570314|CULTURES|DAIRY|-80.848528|80.848541914011989|317|1
35.053394|f37e4dad1a9a74ae2c5878efd6c9a3c8989c15a5|5.61|2014-12-11 17:51:00|80.848351720559364|4|20227900000|11|35.091845860281175|0|25|299|-80.850065|49|35.030252|ANGUS BEEF|0.0|2|ANGUS BEEF BOTTOM ROUND ROAST|b43e43bd71d22e54b77bb1759ac94f3e2dda3d9f|2.656930769193146|35.082633588753836|00202279000006|BEEF|MEAT|-80.848528|80.848539650048323|470|1
35.053394|2830812de095bb860a8134dbcd9d4da3cad99d05|7.18|2015-02-21 18:08:00|80.848351720559364|4|20328400000|11|35.091845859777088|0|25|641|-80.847383|137|35.024464|PREMIUM PORK|3.78|2|PORK LOIN RIB END ROAST|b43e43bd71d22e54b77bb1759ac94f3e2dda3d9f|2.656930769193146|35.082633588753836|00203284000005|PORK|MEAT|-80.848528|80.848541914011989|317|1
35.053394|7022fd0817fe8a97ca507c5f1cd58ae6f83db5dd|3.49|2015-01-07 15:47:00|80.848351720559364|4|664|11|35.091845859777088|0|25|1639|-80.847383|377|35.024464|BULK (DONUTS)|0.5|14|PICK 6  DONUTS|b43e43bd71d22e54b77bb1759ac94f3e2dda3d9f|2.656930769193146|35.082633588753836|00000000006640|DONUTS|BAKERY|-80.848528|80.848541914011989|317|1
35.053394|598df4edde017e1f8d16dfeb0e027881dbf14712|2.27|2015-03-02 17:13:00|80.848351720559364|4|20229600000|11|35.091845859777088|0|25|299|-80.847383|49|35.024464|ANGUS BEEF|0.0|2|ANGUS BEEF EYE OF ROUND STEAK|b43e43bd71d22e54b77bb1759ac94f3e2dda3d9f|2.656930769193146|35.082633588753836|00202296000003|BEEF|MEAT|-80.848528|80.848541914011989|317|1
35.053394|d963cffd313518f831a08902cb7a1115a8441f05|4.0|2014-09-17 18:44:00|80.848351720559364|4||11|35.091845859777088|0|25|565|-80.847383|64|35.024464|REDUCED PRODUCE|0.0|4|PRODUCE REWRAP BY CT|b43e43bd71d22e54b77bb1759ac94f3e2dda3d9f|2.656930769193146|35.082633588753836|00204845000007|FRESH PRODUCE|PRODUCE|-80.848528|80.848541914011989|317|4
35.053394|9cf73869188be7ae4a20eafac49a19aaba409825|2.0|2015-02-06 16:48:00|80.848351720559364|4||11|35.091845859777088|0|25|565|-80.847383|64|35.024464|REDUCED PRODUCE|0.0|4|PRODUCE REWRAP BY CT|b43e43bd71d22e54b77bb1759ac94f3e2dda3d9f|2.656930769193146|35.082633588753836|00204845000007|FRESH PRODUCE|PRODUCE|-80.848528|80.848541914011989|317|2
35.053394|6012f5f3d22bda2225d71d1d45cf3b8d98b08052|1.0|2014-11-16 12:24:00|80.848351720559364|4||11|35.091845859777088|0|25|565|-80.847383|64|35.024464|REDUCED PRODUCE|0.0|4|PRODUCE REWRAP BY CT|b43e43bd71d22e54b77bb1759ac94f3e2dda3d9f|2.656930769193146|35.082633588753836|00204845000007|FRESH PRODUCE|PRODUCE|-80.848528|80.848541914011989|317|1
35.053394|493296aab5f478300d641394775680e67ab2a3ee|3.39|2014-09-12 16:04:00|80.848351720559364|4|7203661037|11|35.091845859777088|0|25|840|-80.847383|102|35.024464|TUBS|0.0|19|HT DELI THIN HONEY HAM|b43e43bd71d22e54b77bb1759ac94f3e2dda3d9f|2.656930769193146|35.082633588753836|00072036610379|LUNCHMEATS|CASE READY MEATS|-80.848528|80.848541914011989|317|1
35.053394|9d8e33c93ddd0df1add48623b28462ba4a8bd57d|4.99|2015-01-15 15:31:00|80.848351720559364|4|5200033776|11|35.091845859777088|0|25|171|-80.847383|20|35.024464|ISOTONIC DRINKS|1.02|1|GATORADE FRUIT PUNCH|b43e43bd71d22e54b77bb1759ac94f3e2dda3d9f|2.656930769193146|35.082633588753836|00052000337754|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.848528|80.848541914011989|317|1
35.053394|7bd3dcdca946b4156ed7e87a536d4f0ed4c20f41|23.49|2014-12-05 16:55:00|80.848351720559364|4|1901461081|11|35.091845859777088|0|25|156|-80.847383|24|35.024464|NFS-DOG FOOD-DRY|0.0|1|IAM HLTHY NATRALS CHCK BRL|b43e43bd71d22e54b77bb1759ac94f3e2dda3d9f|2.656930769193146|35.082633588753836|00019014703579|PET FOOD/SUPPLIES|G1 GROCERY|-80.848528|80.848541914011989|317|1
35.43259|c365f52caaaf656507dd927cea7c5d0a61e96dc4|7.3|2015-01-27 10:56:00|80.606823361882718|4|3800059663|202|35.555289190594081|0|57|61|-80.497332|9|35.667941|RTE CEREAL ADULT|2.3|1|KELLOGG RAISIN BRAN 18|b8d4ad366402ceecc9b9744e4067e6a68ff1def5|8.478254505908305|35.500309569604553|00038000596636|CEREAL|G1 GROCERY|-80.605588|80.606031688625322|178|2
35.43259|64ee2500e4acfafa86b1c4f8a4ba8793b39d5e50|3.78|2015-02-19 12:13:00|1.4057311447477159|4|5100002457|202|0.6184153580092175|0|52|212|-80.605588|33|35.43259|CONDENSED SOUP|1.28|1|CAMP COND 98% FF CREAM MSHROOM|b8d4ad366402ceecc9b9744e4067e6a68ff1def5|8.478254505908305|0.6209993146566879|00051000115515|SOUP|G1 GROCERY|-80.605588|1.406832906106031|202|2
35.43259|b3f984b29e766a8668fbed7187c527a39e37b4f9|2.69|2015-03-09 10:51:00|80.606823361882718|4|7203663217|202|35.555289190594081|0|57|330|-80.497332|55|35.667941|EGGS|0.69|3|HT GRADE A LARGE EGGS 18 CT|b8d4ad366402ceecc9b9744e4067e6a68ff1def5|8.478254505908305|35.500309569604553|00072036632173|EGGS FRESH|DAIRY|-80.605588|80.606031688625322|178|1
35.43259|332fb844fef9246f6e82b2f9a6c00a74021cc09e|2.39|2014-11-15 12:01:00|1.4057311447477159|4|7203663217|202|0.6184153580092175|0|52|330|-80.605588|55|35.43259|EGGS|0.39|3|HT GRADE A LARGE EGGS 18 CT|b8d4ad366402ceecc9b9744e4067e6a68ff1def5|8.478254505908305|0.6209993146566879|00072036632173|EGGS FRESH|DAIRY|-80.605588|1.406832906106031|202|1
35.43259|551fef594658309dc67b517999ea6478c8f6ea5d|2.79|2014-09-25 15:20:00|1.4057311447477159|4|7203698295|202|0.6184153580092175|0|52|81|-80.605588|9|35.43259|RTE CEREAL KIDS|1.29|1|HT CER APPLE CINNAMON|b8d4ad366402ceecc9b9744e4067e6a68ff1def5|8.478254505908305|0.6209993146566879|00072036159977|CEREAL|G1 GROCERY|-80.605588|1.406832906106031|202|1
35.323246|b6541df8ea3b6a69bf75512e1c4bde0c29444e64|0.97|2014-12-08 21:00:00|80.8939826282094|4|3100010903|166|35.500315685183345|0|2|1279|-80.992182|48|35.103409|SINGLE SERVE FLAVOR|0.0|5|BANQUET SALISBURY STEAK MEAL|bbf7c786890668b7a563a972b697d80accbe2130|12.235125820953641|35.490689277687849|00031000109059|FROZEN MEALS|FROZEN|-80.945176|80.945718785088175|88|1
35.323246|515d5e480b8e1fadadabcf06a63f1012fd9d7a58|0.65|2014-12-24 14:01:00|80.8939826282094|4|5000042264|166|35.500315470728218|0|2|154|-80.994596|24|35.061685|NFS-CAT FOOD WET|0.1|1|FSK TST PATE CHK&OCNFSH W/CHS|bbf7c786890668b7a563a972b697d80accbe2130|12.235125820953641|35.490689277687849|00050000582082|PET FOOD/SUPPLIES|G1 GROCERY|-80.945176|80.945815494055552|475|1
35.037115|47cc3a7e436125eaa1174f6393840a46fbbf8f98|3.99|2014-11-25 18:16:00|80.805842308733688|1|3425600064|27|35.050830289023082|0|49|577|-80.848528|136|35.053394|OTHER MERCH FR MSC JUICE|0.49|4|HT APPLE CIDER, 64 OZ|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00072036880888|OTHER MERCHANDISE|PRODUCE|-80.8062|80.806200361802553|11|1
35.037115|23fede30327c716a08c34335ab1d5a2703d13244|6.94|2015-01-07 09:06:00|80.805842308733688|1|7203659020|27|35.050830286185757|0|49|312|-80.758228|51|34.95459|BUTTER|0.0|3|HARRIS TEETER UNSALTED BUTTER|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00072036590213|BUTTER & MARGARINE|DAIRY|-80.8062|80.806210781648971|182|2
35.037115|ba3802aee52dfe1e78902f10fd5993b57bf5b441|6.57|2014-12-09 09:17:00|80.805842308733688|1|8000000672|27|35.050830286185757|0|49|190|-80.758228|29|34.95459|TUNA-CANNED|1.57|1|STARKIST TUNA SOLID WHT ALB|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00080000006721|SEAFOOD-CANNED|G1 GROCERY|-80.8062|80.806210781648971|182|3
35.037115|9774d5ce1f4acb1a4cbff090d4ab9965760b0837|3.99|2014-11-24 12:28:00|80.805842308733688|1|8390000649|27|35.050830286185757|0|49|365|-80.758228|56|34.95459|REFRIGERATED TEAS|0.99|3|GOLD PEAK SWEET BLACK TEA|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00083900006495|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.8062|80.806210781648971|182|1
35.037115|c18400d663b69b6ef46d1f460fa451722ab9f1c3|2.99|2015-01-03 15:09:00|1.4091206135396188|1|8186422116|27|0.611513017149893|0|47|583|-80.8062|136|35.037115|NUTS|0.0|4|SALTED PEANUTS IN-SHELL|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00081864221169|OTHER MERCHANDISE|PRODUCE|-80.8062|1.4103342460250419|27|1
35.037115|ce186dc49e33d6c960f7f95483d6e66bf7825c39|5.59|2015-02-10 13:52:00|1.4091206135396188|1|9830800202|27|0.611513017149893|0|47|211|-80.8062|33|35.037115|BOUILLON|1.6|1|BETTER THAN BOUILLON BEEF|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00098308002031|SOUP|G1 GROCERY|-80.8062|1.4103342460250419|27|1
35.037115|8f1d1c0520c5030a6a1d0a4375a438ddb416da95|6.39|2015-02-21 12:31:00|1.4091206135396188|1|7403000003|27|0.611513017149893|0|47|2017|-80.8062|505|35.037115|STRETCHED CURD CHEESE|0.0|6|SORRENTO WHOLE MILK MOZZARELA|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00074030000033|SPECIALTY CHEESE|DELI|-80.8062|1.4103342460250419|27|1
35.037115|de15be4743b722408d1d4dec97815f4fe59404d6|3.34|2015-02-25 18:02:00|1.4091206135396188|1|7110000407|27|0.611513017149893|0|47|183|-80.8062|28|35.037115|SALAD DRESSINGS-DRY|0.0|1|HVR DIP MIX RANCH|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00071100004038|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.8062|1.4103342460250419|27|2
35.037115|4b402507c46a9c484d746d58a5b2b771e424189e|4.69|2014-12-04 16:31:00|1.4091206135396188|1|7468309950|27|0.611513017149893|0|47|1220|-80.8062|275|35.037115|PASTA SC PREMIUM|0.0|1|EMERIL PASTA SC VODKA|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00074683099477|PASTA SAUCES|G1 GROCERY|-80.8062|1.4103342460250419|27|1
35.037115|42e3de253029735c15b484e693d23905eb7bdbb5|4.97|2014-09-29 16:51:00|80.805842308733688|1|7229000227|27|35.050830288299345|0|49|1271|-80.770346|41|35.052812|PROTEIN BREAKFAST|0.0|5|TENN PRIDE CHKN&BTTRMLK BISC|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00072290022406|BREAKFAST FOODS FROZEN|FROZEN|-80.8062|80.806205454227992|40|1
35.037115|133fb61b271613149c511294e88777547141fbbb|4.99|2015-01-22 14:44:00|80.805842308733688|1|7468309950|27|35.050830288299345|0|49|1220|-80.770346|275|35.052812|PASTA SC PREMIUM|1.0|1|EMERIL PASTA SC VODKA|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00074683099477|PASTA SAUCES|G1 GROCERY|-80.8062|80.806205454227992|40|1
35.037115|2b173f9f7bd833bd0eb573c9624df4e2f493ea8f|0.79|2015-01-28 11:52:00|80.805842308733688|1||27|35.050830286185757|0|49|532|-80.758228|64|34.95459|FRESH CUCUMBERS|0.0|4|COO CUCUMBERS S/S|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00204062000002|FRESH PRODUCE|PRODUCE|-80.8062|80.806210781648971|182|1
35.037115|8068a65499118fc9750cc7c90c8949336f16cfc2|0.79|2015-02-24 18:00:00|1.4091206135396188|1||27|0.611513017149893|0|47|532|-80.8062|64|35.037115|FRESH CUCUMBERS|0.0|4|COO CUCUMBERS S/S|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00204062000002|FRESH PRODUCE|PRODUCE|-80.8062|1.4103342460250419|27|1
35.037115|2c620cbe776949c1ddb77ce9d8d154b92ac62cdd|0.79|2015-03-01 14:31:00|1.4091206135396188|1||27|0.611513017149893|0|47|532|-80.8062|64|35.037115|FRESH CUCUMBERS|0.0|4|COO CUCUMBERS S/S|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00204062000002|FRESH PRODUCE|PRODUCE|-80.8062|1.4103342460250419|27|1
35.037115|6d3af103d2371c030f70a07616011786819f6220|0.89|2014-12-17 10:42:00|80.805842308733688|1||27|35.050830286185757|0|49|532|-80.758228|64|34.95459|FRESH CUCUMBERS|0.0|4|COO CUCUMBERS S/S|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00204062000002|FRESH PRODUCE|PRODUCE|-80.8062|80.806210781648971|182|1
35.037115|a7619c86aac1fb0825f052d3948de3424f37e39e|9.42|2014-12-13 18:15:00|1.4091206135396188|1||27|0.611513017149893|0|47|562|-80.8062|64|35.037115|FRESH CUT FRUIT|0.0|4|PINEAPPLE RING SLICES|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00204347000000|FRESH PRODUCE|PRODUCE|-80.8062|1.4103342460250419|27|2
35.037115|7ee567464f01c8cd982d2cba81ed2b4026b2db3c|3.29|2014-12-23 16:09:00|1.4091206135396188|1|60502177400|27|0.611513017149893|0|47|192|-80.8062|30|35.037115|COOKING SPRAYS|0.79|1|BAKERS JOY BAKING SPRAY|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00605021774000|SHORTENING/OIL|G1 GROCERY|-80.8062|1.4103342460250419|27|1
35.037115|79133ea2af6f4c4d15795fe44f6496a1ce7318fa|1.99|2015-01-17 09:44:00|1.4091206135396188|1|5849672304|27|0.611513017149893|0|47|168|-80.8062|24|35.037115|NFS-CAT TREATS|0.32|1|TEMPTATIONS TMBLR SALMN/TURKY|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00023100109282|PET FOOD/SUPPLIES|G1 GROCERY|-80.8062|1.4103342460250419|27|1
35.037115|2e0b2c3a796dd66edca840280cde97e72e6c1374|1.29|2015-03-01 21:00:00|1.4091206135396188|1|2200000488|27|0.611513017149893|0|47|48|-80.8062|7|35.037115|REGISTER GUM|0.0|1|(FE)ORBIT PEPPERMINT GUM 14PC|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00022000004864|CANDY|G1 GROCERY|-80.8062|1.4103342460250419|27|1
35.037115|51540cb59059f9796598d1ee7ba351d88f36080a|3.78|2015-01-26 14:03:00|1.4091206135396188|1|2000000065|27|0.611513017149893|0|47|1275|-80.8062|50|35.037115|BOX VEG|0.78|5|GG BROCCOLI SPEAR NO SAUCE|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00020000174839|VEGETABLES-FROZEN|FROZEN|-80.8062|1.4103342460250419|27|2
35.037115|229b688fcc96d7a72dd52063ca613a7f302c6b55|3.29|2014-12-14 14:41:00|1.4091206135396188|1|2840014741|27|0.611513017149893|0|47|205|-80.8062|31|35.037115|REMAINING SNACKS|0.0|1|SUNCHIPS REGULAR|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00028400147415|SNACKS|G1 GROCERY|-80.8062|1.4103342460250419|27|1
35.037115|7b95d46115baa527fe8b96d40c685d48608df13d|2.49|2015-01-05 17:11:00|1.4091206135396188|1|2840005658|27|0.611513017149893|0|47|206|-80.8062|31|35.037115|FRONT END SNACKS|0.0|1|LAYS CLASSIC SINGLES|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00028400056588|SNACKS|G1 GROCERY|-80.8062|1.4103342460250419|27|1
35.037115|9e45000f0b06c7a77452b41c24df7939a0308f8b|8.98|2014-11-11 17:01:00|80.805842308733688|1|2840009217|27|35.050830288299345|0|49|1981|-80.770346|480|35.052812|CHIPS|0.0|6|STACY'S PITA CHIPS NAKED|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00028400092173|DRY GOODS|DELI|-80.8062|80.806205454227992|40|2
35.037115|f9b348e00f3fd9f87a6a5b008ef2fd449545a7f5|3.0|2015-02-06 19:08:00|1.4091206135396188|1||27|0.611513017149893|0|47|1635|-80.8062|375|35.037115|BULK (BAGELS)|0.0|14|BULK  BAGELS|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00072036955500|BAGELS|BAKERY|-80.8062|1.4103342460250419|27|4
35.037115|e7d1101347f2b9fecfda33bb0121ab4de31a80d5|3.99|2015-02-01 14:05:00|1.4091206135396188|1|7203695451|27|0.611513017149893|0|47|2003|-80.8062|495|35.037115|FFM GREEN SALADS|1.0|6|GARDEN SALAD|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00072036954510|GREEN SALADS|DELI|-80.8062|1.4103342460250419|27|1
35.037115|5622f558074b79a6648e26621cb375f5c1c051b8|3.69|2014-09-16 14:59:00|1.4091206135396188|1|7203695783|27|0.611513017149893|0|47|1631|-80.8062|373|35.037115|THAW & SELL (ROLLS)|0.0|14|RICH & BUTTERY BRIOCHE ROLLS|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00072036957832|ROLLS|BAKERY|-80.8062|1.4103342460250419|27|1
35.037115|ba517d03d9d5516858d311fb2a092bea522f20c9|13.96|2014-12-18 08:56:00|80.805842308733688|1|74759961422|27|35.050830286185757|0|49|727|-80.758228|7|34.95459|SEASONAL CANDY-SINGLE FAC|1.96|1|I/O(C14)GHIR PEPP BARK BARS|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00747599614224|CANDY|G1 GROCERY|-80.8062|80.806210781648971|182|4
35.037115|23e59268f58f2a60d7dd5310c6816206b8bc451f|5.99|2014-10-30 18:01:00|1.4091206135396188|1|79285001444|27|0.611513017149893|0|47|3272|-80.8062|1023|35.037115|NATURAL/ORGANIC PRODUCT|1.2|17|BURTS B TOWELETTES PEACH|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00792850018167|NATURAL PERSONAL CARE|HBC|-80.8062|1.4103342460250419|27|1
35.037115|153bdee693c22a5dd8591a4281775d5ae21bed5f|3.95|2014-10-24 16:12:00|1.4091206135396188|1|1410007467|27|0.611513017149893|0|47|1025|-80.8062|162|35.037115|WHITE|0.0|7|PEP FH SOURDOUGH WP BRD PP|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00014100074670|SLICED BREAD|COMMERCIAL BAKERY|-80.8062|1.4103342460250419|27|1
35.037115|30b49617641115225efb1417ca00bbdb9baafe6a|3.49|2014-10-27 16:30:00|1.4091206135396188|1|7146426040|27|0.611513017149893|0|47|577|-80.8062|136|35.037115|OTHER MERCH FR MSC JUICE|0.0|4|BOLTHOUSE AMAZING MANGO|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00071464309503|OTHER MERCHANDISE|PRODUCE|-80.8062|1.4103342460250419|27|1
35.037115|33a9fa0282fce75981697bf9b107fb4a266a6127|6.79|2014-10-09 14:23:00|80.805842308733688|1|4900002890|27|35.05083028877484|0|49|55|-80.816172|8|35.059823|REGULAR|1.8|23|CLASSIC 12OZ 12PK FRIDGE CAN|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00049000028904|CARBONATED BEVERAGES|BEVERAGE|-80.8062|80.806203207767311|66|1
35.037115|d9d3d6266e51e48986bf6d8b41111e584c34aee3|6.79|2014-10-15 10:40:00|80.805842308733688|1|4900002890|27|35.050830286185757|0|49|55|-80.758228|8|34.95459|REGULAR|1.8|23|CLASSIC 12OZ 12PK FRIDGE CAN|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00049000028904|CARBONATED BEVERAGES|BEVERAGE|-80.8062|80.806210781648971|182|1
35.037115|60a72b516f1bf8ef70325a003b20c285d1a95294|6.99|2015-01-13 14:38:00|1.4091206135396188|1|4900002890|27|0.611513017149893|0|47|55|-80.8062|8|35.037115|REGULAR|2.0|23|CLASSIC 12OZ 12PK FRIDGE CAN|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00049000028904|CARBONATED BEVERAGES|BEVERAGE|-80.8062|1.4103342460250419|27|1
35.037115|c8bf65e2411f918dd8b7e139e79ecdf67b82df82|6.79|2014-11-22 16:44:00|1.4091206135396188|1|4900002890|27|0.611513017149893|0|47|55|-80.8062|8|35.037115|REGULAR|1.8|23|CLASSIC 12OZ 12PK FRIDGE CAN|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00049000028904|CARBONATED BEVERAGES|BEVERAGE|-80.8062|1.4103342460250419|27|1
35.037115|33cd5c4a13fb09a131a614db9c3fdd302dfc2e64|1.99|2014-09-16 10:20:00|80.805842308733688|1|5849672304|27|35.050830286185757|0|49|168|-80.758228|24|34.95459|NFS-CAT TREATS|0.2|1|WHISKAS TEMPTATIONS SAVORY SAL|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00058496723040|PET FOOD/SUPPLIES|G1 GROCERY|-80.8062|80.806210781648971|182|1
35.037115|b0ebcf2e0612dc8e7034a18e900c655c9a8356f5|2.79|2015-02-15 15:42:00|80.805842308733688|1|4200061045|27|35.050830287558419|0|49|423|-80.771677|72|35.066546|NFS-DISPOSE PLATES/BOWLS|0.0|1|DIXIE HVY DUTY 8 1/2 PLT 45CT|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00042000610452|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.8062|80.806207750487758|45|1
35.037115|708c4a88de5f4dab68084e664be087d894e00056|2.59|2014-12-26 15:01:00|1.4091206135396188|1|1480000034|27|0.611513017149893|0|47|128|-80.8062|20|35.037115|APPLE JUICE-SHELF|0.0|1|MOTTS NATURAL APPLE JUICE|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00014800316568|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.8062|1.4103342460250419|27|1
35.037115|04cce1073e556bf8e609c57293cd1f4025559987|6.98|2014-12-13 08:50:00|80.805842308733688|1|88513178282|27|35.050830286185757|0|49|5151|-80.758228|1300|34.95459|FEEDING ACCESSORIES|0.0|17|GERBER SOFT BITE SPOON|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00885131782823|BABY ACCESSORY|HBC|-80.8062|80.806210781648971|182|2
35.037115|db29d4535f621c3e125665923f2f7deb33ec77f4|3.99|2014-10-03 17:16:00|1.4091206135396188|1|64767100014|27|0.611513017149893|0|47|581|-80.8062|136|35.037115|FRESH SALSA|0.0|4|GFG JACKS SPECIAL MILD SALSA|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00647671000153|OTHER MERCHANDISE|PRODUCE|-80.8062|1.4103342460250419|27|1
35.037115|98bcbdd785b69d967a622f86608fe2e1d6fa36c4|6.49|2015-01-10 13:31:00|80.805842308733688|1|63256500009|27|35.050830286185757|0|49|31|-80.758228|4|34.95459|NON CARBONATED WATER|1.0|1|FIJI WATER 16.9OZ 6PK|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00632565000098|BOTTLED WATER|G1 GROCERY|-80.8062|80.806210781648971|182|1
35.037115|12769ca0a51fe6fba5d18c83a49a55268fa01d3c|3.69|2014-12-16 12:31:00|80.805842308733688|1|73599509111|27|35.050830286185757|0|49|71|-80.758228|11|34.95459|GROC CONDIMENTS MARINADE|0.7|1|MOORES MARINADE TERIYAKI|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00735995091121|CONDIMENTS|G1 GROCERY|-80.8062|80.806210781648971|182|1
35.037115|7c6b458d6434be78e1ee777840793ace90a4d119|2.5|2014-09-22 15:59:00|80.805842308733688|1|81851201703|27|35.050830288299345|0|49|43|-80.770346|6|35.052812|INSTANT BREAKFAST-POWDERED|0.51|1|SPROUT RSE PEACH ORG YOG SMOTH|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00818512017047|BREAKFAST FOODS|G1 GROCERY|-80.8062|80.806205454227992|40|1
35.037115|5a8f1867facf2f2d9f5163460022acbb994bca16|4.29|2014-10-19 18:07:00|80.805842308733688|1|74236526405|27|35.050830288299345|0|49|345|-80.770346|57|35.052812|ORGANIC MILK|0.0|3|HORIZON ORGANIC 2% MILK.|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00742365264252|MILK|DAIRY|-80.8062|80.806205454227992|40|1
35.037115|e1e5255e95be0deea34889630dc876f88ae01606|4.97|2015-01-21 12:00:00|80.805842308733688|1|31015808504|27|35.050830286185757|0|49|4086|-80.758228|1080|34.95459|TOOTHPASTE-SENSITIVE|0.0|17|SENSODYNE TARTAR CONTRL TPASTE|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00310158085041|ORAL HYGIENE|HBC|-80.8062|80.806210781648971|182|1
35.037115|2ec59cb2a6734fb58d68f0a4dbdbfbe484ab3573|5.99|2014-11-13 18:29:00|80.805842308733688|1|81034700605|27|35.050830286185757|0|49|1074|-80.758228|219|34.95459|INDIAN-SPEC|0.0|1|KOHINOOR MADRAS CURRY PWDR|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00810347006050|SPECIALTY-ETHNIC FOODS|G1 GROCERY|-80.8062|80.806210781648971|182|1
35.037115|1b7459b5bb2d815046a13c48218fc46e7ffd07c9|3.99|2014-09-21 18:23:00|1.4091206135396188|1|1906301228|27|0.611513017149893|0|47|31|-80.8062|4|35.037115|NON CARBONATED WATER|2.0|1|VYFINE FRUIT 2 O LEMON 6PK|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00019063232310|BOTTLED WATER|G1 GROCERY|-80.8062|1.4103342460250419|27|1
35.037115|f241172cda2fba309e995531b555f11aabb22533|3.99|2014-12-24 12:47:00|80.805842308733688|1|1862753422|27|35.05083028877484|0|49|1269|-80.816172|41|35.059823|BREAKFAST SYRUP CARRIER|0.0|5|KASHI BLUEBERRY WAFFLE|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00018627534228|BREAKFAST FOODS FROZEN|FROZEN|-80.8062|80.806203207767311|66|1
35.037115|725897e4c517ea6f771dbd669e8747f49f3dbdca|2.79|2015-01-12 19:56:00|80.805842308733688|1|1600015110|27|35.050830288334097|0|49|205|-80.847383|31|35.024464|REMAINING SNACKS|0.0|1|BUGLES ORIGINAL|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00016000283701|SNACKS|G1 GROCERY|-80.8062|80.806205322259999|317|1
35.037115|8d41587e1508b92eb1d533f6a54a11da83506c2d|12.99|2014-11-01 17:20:00|80.805842308733688|1|7203695587|27|35.05083028877484|0|49|1707|-80.816172|387|35.059823|MESSAGE|3.0|14|12 INCH MESSAGE COOKIE|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00072036955876|COOKIES|BAKERY|-80.8062|80.806203207767311|66|1
35.037115|5b725c45da69a1735750229e558ad8e29217f694|4.99|2014-12-12 20:42:00|1.4091206135396188|1|4850002141|27|0.611513017149893|0|47|1407|-80.8062|57|35.037115|ICED COFFEE|0.5|3|I/OSTARBUCKS PEPPERMINT MOCHA|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00048500022450|MILK|DAIRY|-80.8062|1.4103342460250419|27|1
35.037115|3086bc49fc1bdc525538fd308a3861ce49e0c551|0.6|2015-01-26 17:40:00|1.4091206135396188|1||27|0.611513017149893|0|47|502|-80.8062|64|35.037115|FRESH BANANAS|0.0|4|BANANAS, YELLOW|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00204011000008|FRESH PRODUCE|PRODUCE|-80.8062|1.4103342460250419|27|1
35.037115|1f5ab2111114f222d5e94174b5a71a137dff974f|3.99|2014-10-21 17:29:00|1.4091206135396188|1|8259272215|27|0.611513017149893|0|47|577|-80.8062|136|35.037115|OTHER MERCH FR MSC JUICE|0.0|4|NAKED PROTEIN DOUBLE BERRY|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00082592631954|OTHER MERCHANDISE|PRODUCE|-80.8062|1.4103342460250419|27|1
35.037115|119ef671ae070d4d1985c3d58054fcb22b9dedfe|12.98|2014-12-13 08:54:00|80.805842308733688|1|3160066801|27|35.050830286185757|0|49|5519|-80.758228|1506|34.95459|SHOE CARE-ACCESSORIES|0.0|18|SMALL FEET HEEL LINERS|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00031600668048|SHOE CARE/LACES/SEWING|GM|-80.8062|80.806210781648971|182|2
35.037115|75a4a0e8448192c7bccb60d15b3d7284efc66aaa|3.49|2015-02-18 17:24:00|1.4091206135396188|1|81989801902|27|0.611513017149893|0|47|1251|-80.8062|12|35.037115|WHOLESOME COOKIES|0.0|1|SNACKWELL DEVIL CAKE COOKIE|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00819898019007|COOKIES|G1 GROCERY|-80.8062|1.4103342460250419|27|1
35.037115|ae98d73077f0bf162c96fad98bde2a7bbf6d1d07|6.99|2015-02-14 12:47:00|1.4091206135396188|1|7403008182|27|0.611513017149893|0|47|2017|-80.8062|505|35.037115|STRETCHED CURD CHEESE|0.0|6|SORRENTO FRESH MOZZARELLA|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00074030081827|SPECIALTY CHEESE|DELI|-80.8062|1.4103342460250419|27|1
35.037115|9b92d79e3fd73db9b6f3532e9b8eb65aec3d6716|19.77|2014-12-23 16:10:00|1.4091206135396188|1|7478037743|27|0.611513017149893|0|47|30|-80.8062|4|35.037115|CARBONATED WATER|1.7999999999999998|1|PERRIER SPARK LIME 10PK|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00074780333566|BOTTLED WATER|G1 GROCERY|-80.8062|1.4103342460250419|27|3
35.037115|010b6827984d336b7704bb5833a00dbb20e8d0b9|7.08|2014-11-18 16:51:00|80.805842308733688|1|7203676122|27|35.050830288299345|0|49|1218|-80.770346|273|35.052812|ASIAN OTHER|0.0|1|HT TRADER COCONUT MILK|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00072036761224|ASIAN PREP. FOODS|G1 GROCERY|-80.8062|80.806205454227992|40|4
35.037115|8fc93248c075d0d1b6301be76632908c96e86143|12.6|2014-10-01 10:55:00|80.805842308733688|1|4132100541|27|35.050830286185757|0|49|184|-80.758228|28|34.95459|SALAD DRESSINGS-LIQUID|1.58|1|D  WISHBONE DRS LT RANCH|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00041000005732|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.8062|80.806210781648971|182|4
35.037115|3eb82ba96dd3de744b3d7a657c7b72008cccb075|24.950000000000003|2014-12-11 09:03:00|80.805842308733688|1|4082201114|27|35.050830286185757|0|49|1878|-80.758228|435|34.95459|HUMMUS|0.0|6|CLASSIC HUMMUS|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00040822011143|SALADS|DELI|-80.8062|80.806210781648971|182|5
35.037115|1ded7434ef42f9ebc6ba5bb1d53698819cd1c58d|8.78|2015-01-15 14:01:00|80.805842308733688|1|1356211105|27|35.05083028877484|0|49|1200|-80.816172|6|35.059823|FRUIT SNACKS|2.78|1|ANNIES FRT SNACK BERRY PATCH|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00013562111053|BREAKFAST FOODS|G1 GROCERY|-80.8062|80.806203207767311|66|2
35.037115|d389847929b9b81eb134211a7b2fd681f7d60427|3.99|2014-12-10 20:14:00|80.805842308733688|1|60659701012|27|35.05083028877484|0|49|312|-80.816172|51|35.059823|BUTTER|0.49|3|I/OKELLER'S CHRISTMAS TREE BTR|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00606597010127|BUTTER & MARGARINE|DAIRY|-80.8062|80.806203207767311|66|1
35.037115|d9ad920ac1213a66ccea2efa5901844de5700f22|1.94|2014-11-26 17:32:00|1.4091206135396188|1|7203604053|27|0.611513017149893|0|47|51|-80.8062|7|35.037115|MARSHMALLOWS|0.2|1|HT MINI MARSHMALLOW|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00072036040534|CANDY|G1 GROCERY|-80.8062|1.4103342460250419|27|2
35.037115|d5a65055cba70a53a367ecc3bab233f9887c6097|1.39|2014-11-01 11:35:00|80.805842308733688|1|5210094269|27|35.050830286185757|0|49|80|-80.758228|34|34.95459|SEASONING PACKETS|0.39|1|CHILI SEASONING LESS SODIUM|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00052100942698|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.8062|80.806210781648971|182|1
35.037115|c02c168e5f4d845ebfbce2ec85e5c1296523cc48|9.02|2015-02-27 15:59:00|80.805842308733688|1|20165700000|27|35.050830285488026|0|49|297|-80.78468|49|35.096737|GROUND BEEF|1.0|2|HT GRND BF CHUCK 80% LEAN CUST|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|35.053350220983141|00201693000005|BEEF|MEAT|-80.8062|80.806212033196402|30|2
35.037115|54ee9b26374ee974b80c8022e0280b62462c7c14|2.75|2014-12-09 16:06:00|1.4091206135396188|1|2500001309|27|0.611513017149893|0|47|121|-80.8062|20|35.037115|ASEPTIC JUICES|0.76|1|HI-C FLASHIN FRUIT PUNCH 10 PK|bcca3d8377d8ff21c65703d1c6a43a1b84c5a4e7|0.9476933504786241|0.61242566243833529|00025000010804|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.8062|1.4103342460250419|27|1
35.43259|d0130e3a7062a6d0744895f2213f8270b60fde6d|7.97|2015-01-07 08:17:00|80.607132136635443|4|3700009614|202|35.466994523635648|0|9|3774|-80.762919|1070|35.442529|CLINICAL-FEMALE|0.0|17|SECRET CLINICAL INV LVND|c4f8fb422152b734a332c81f57277bfa5d7b2c01|2.3772699485782804|35.47365851958088|00037000885191|DEODORANT|HBC|-80.605588|80.605613965965063|471|1
35.43259|729589b03a0b479009bb51412d24e58662293eee|26.25|2015-01-08 19:57:00|80.607132136635443|4|4650075362|202|35.466994526308127|0|9|393|-80.662946|68|35.412407|NFS-AIR FRESHENERS|1.5|1|GLADE CANDLE CUSTRD & APPLE|c4f8fb422152b734a332c81f57277bfa5d7b2c01|2.3772699485782804|35.47365851958088|00046500753664|FRESHENERS/DEODORIZERS|G1 GROCERY|-80.605588|80.60560792803318|68|7
35.43259|0482350008bb3afc94702bf7ca6c3df8e682e6d1|1.06|2015-01-12 13:24:00|80.607132136635443|4||202|35.466994523635648|0|9|502|-80.762919|64|35.442529|FRESH BANANAS|0.0|4|BANANAS, YELLOW|c4f8fb422152b734a332c81f57277bfa5d7b2c01|2.3772699485782804|35.47365851958088|00204011000008|FRESH PRODUCE|PRODUCE|-80.605588|80.605613965965063|471|1
35.43259|e2e01a5251665c773d4fd409065f6d918228e396|0.99|2015-02-07 19:16:00|1.4057311447477159|4|1780014597|202|0.6184153580092175|0|52|154|-80.605588|24|35.43259|NFS-CAT FOOD WET|0.0|1|ONE PREMIUM PATE TENDER CHICKN|c4f8fb422152b734a332c81f57277bfa5d7b2c01|2.3772699485782804|0.6209993146566879|00017800145978|PET FOOD/SUPPLIES|G1 GROCERY|-80.605588|1.406832906106031|202|1
35.43259|c0217c7693824e98f73cd19719eabc9619360794|2.19|2015-01-08 19:18:00|1.4057311447477159|4|3760003895|202|0.6184153580092175|0|52|659|-80.605588|103|35.43259|CHILDRENS LUNCH SNACKS|0.0|19|HORMEL REV BACON CLUB|c4f8fb422152b734a332c81f57277bfa5d7b2c01|2.3772699485782804|0.6209993146566879|00037600207706|LUNCH SNACKS|CASE READY MEATS|-80.605588|1.406832906106031|202|1
35.03469|c99b31c3c77189750af542f06b274e2c64da2c25|7.99|2014-10-14 17:42:00|1.4132775322775095|3|8378322822|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|SIERRA NEVADA SEASONAL 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00083783228229|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|7f53d08ad4765711018c1fc175fb1437101190bd|9.99|2015-01-30 18:51:00|1.4132775322775095|3|8769200004|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|SAM ADAMS WINTER SEASONAL 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00087692000044|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|52c67d9a22f8f394d68a1b9caa397a3f9dacf832|7.99|2015-01-01 16:42:00|1.4132775322775095|3|8130859187|82|0.6114706929155321|0|58|9948|-80.97058|886|35.03469|NFS-PREM-CAB SAUVIGNON|0.0|13|CUPCAKE CAB SAUV|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00081308591872|PREMIUM ($8-$10.99)|WINE|-80.97058|1.4132032182494703|82|1
35.03469|533e7d2a17c83e4117b83bf57a3d3b50df200403|9.99|2015-01-22 18:59:00|1.4132775322775095|3|8769200004|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|SAM ADAMS WINTER SEASONAL 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00087692000044|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|d816dd177bd5f1c69c7d874aebc2ea7935d9a87f|7.99|2015-01-09 19:15:00|1.4132775322775095|3|8130859187|82|0.6114706929155321|0|58|9948|-80.97058|886|35.03469|NFS-PREM-CAB SAUVIGNON|0.0|13|CUPCAKE CAB SAUV|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00081308591872|PREMIUM ($8-$10.99)|WINE|-80.97058|1.4132032182494703|82|1
35.03469|e7ccb400eab818d44a97f2e12d73a07447990267|9.99|2015-03-06 18:51:00|1.4132775322775095|3|8769200004|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|SAM ADAMS WINTER SEASONAL 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00087692000044|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|18f1274d2cb98e6ebbf7803eb834f8ef4430a061|9.99|2015-02-11 18:29:00|1.4132775322775095|3|8769200004|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|SAM ADAMS WINTER SEASONAL 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00087692000044|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|5281fd28582ea354fb407b4cb9b28efb4357fe74|9.99|2015-02-07 10:28:00|1.4132775322775095|3|8769200004|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|SAM ADAMS WINTER SEASONAL 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00087692000044|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|179a22ba8891dce3d4785469faa80be364b7bccd|9.99|2015-01-20 18:50:00|1.4132775322775095|3|8769200004|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|SAM ADAMS WINTER SEASONAL 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00087692000044|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|6ddee6971ec769412807aeaf5599eceecbf6afc0|9.99|2015-02-14 13:34:00|1.4132775322775095|3|8769200004|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|SAM ADAMS WINTER SEASONAL 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00087692000044|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|5f36c601db000a912618b481364b8b5051c0a63b|9.99|2015-02-24 19:21:00|1.4132775322775095|3|8769200004|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|SAM ADAMS WINTER SEASONAL 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00087692000044|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|dbf270f174e894b99a3309c33df70b84d06ef709|9.99|2015-01-28 19:24:00|1.4132775322775095|3|8769200004|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|SAM ADAMS WINTER SEASONAL 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00087692000044|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|f92095bd7d924085da1c3bebf0f12ba9eb6e54a5|9.99|2015-02-26 18:46:00|1.4132775322775095|3|8769200004|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|SAM ADAMS WINTER SEASONAL 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00087692000044|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|da20b8de8a2a784197cb12da2ea93c78655dee2b|9.99|2015-03-04 19:28:00|1.4132775322775095|3|8769200004|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|SAM ADAMS WINTER SEASONAL 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00087692000044|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|58ab4694998aa44ab71bc566c5b5e1b67e985ad7|9.99|2015-01-24 12:59:00|1.4132775322775095|3|8769200004|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|SAM ADAMS WINTER SEASONAL 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00087692000044|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|e334c43b8dad183f9ba5e0d3bb7980dd75538c89|7.99|2015-01-26 19:25:00|1.4132775322775095|3|8069611122|82|0.6114706929155321|0|58|9935|-80.97058|885|35.03469|NFS POP CAB SAUV|0.0|13|BV COASTAL CAB SAUV|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00080696111228|POPULAR (4-$7.99)|WINE|-80.97058|1.4132032182494703|82|1
35.03469|1e4ccc01ab151893b63d753e617d2600a707dd2e|7.99|2015-01-07 18:41:00|1.4132775322775095|3|8069611122|82|0.6114706929155321|0|58|9935|-80.97058|885|35.03469|NFS POP CAB SAUV|0.0|13|BV COASTAL CAB SAUV|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00080696111228|POPULAR (4-$7.99)|WINE|-80.97058|1.4132032182494703|82|1
35.03469|cae82a9c2a71c1c82203bb9ddda993c1d7cbf8f6|9.99|2014-12-20 13:44:00|1.4132775322775095|3|71280824276|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|HIGHLAND BLK MOCHA STOUT 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00712808242765|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|630436de4dcdffc2083ad246a52c9b015eddc595|8.99|2014-10-28 18:43:00|1.4132775322775095|3|71280824276|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|HIGHLAND BLK MOCHA STOUT 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00712808242765|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|7d109992515d3756f615022a80b32ec33c1212a5|9.99|2015-01-13 18:26:00|1.4132775322775095|3|71280824276|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|HIGHLAND BLK MOCHA STOUT 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00712808242765|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|62da95c011de61b41df56803a199fa97b4511404|9.99|2015-02-02 17:47:00|1.4132775322775095|3|71280824276|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|HIGHLAND BLK MOCHA STOUT 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00712808242765|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|edbf2e07be408a23d7a8ccc34da1a9349f52ef30|8.99|2014-11-03 19:17:00|1.4132775322775095|3|71280824276|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|HIGHLAND BLK MOCHA STOUT 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00712808242765|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|ca1855bbe25169a06485610db53141b0559e8ae3|8.99|2014-11-26 18:50:00|1.4132775322775095|3|71280824276|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|HIGHLAND BLK MOCHA STOUT 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00712808242765|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|5544fc33d3cf579c40a54cfd385aa256a821e1ac|9.99|2015-02-04 19:09:00|1.4132775322775095|3|71280824276|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|HIGHLAND BLK MOCHA STOUT 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00712808242765|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|d5b45307d12c9b36a471accbe479f751c4a8f223|8.99|2014-11-18 18:09:00|1.4132775322775095|3|71280824276|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|HIGHLAND BLK MOCHA STOUT 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00712808242765|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|5a0cc9e20babe2872352a5c694562998c16dc193|8.99|2014-11-09 13:10:00|1.4132775322775095|3|71280824276|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|HIGHLAND BLK MOCHA STOUT 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00712808242765|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|e28241bac1fd328acdac9f9eb1ff0d1b37bf2b23|8.99|2014-12-08 18:52:00|1.4132775322775095|3|71280824276|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|HIGHLAND BLK MOCHA STOUT 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00712808242765|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|7ce00c60dc7cd0c678ae5e3b088fd999a056b764|9.99|2014-12-30 18:22:00|1.4132775322775095|3|71280824276|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|HIGHLAND BLK MOCHA STOUT 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00712808242765|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|2b84a860e14d50e0ae60f86aab276d3a9eae4c87|9.99|2015-01-11 17:52:00|1.4132775322775095|3|71280824276|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|HIGHLAND BLK MOCHA STOUT 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00712808242765|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|9e6df2fbf79f38f550ccf746e6d506b3d1fb5173|1.47|2014-10-25 15:35:00|1.4132775322775095|3|7203618340|82|0.6114706929155321|0|58|6152|-80.97058|1546|35.03469|BULB-HOUSEHOLD-PRIVATE LABEL|0.0|18|HT 60 WATT SOFT WHITE|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00072036183415|LIGHT BULBS/ELECTRICAL|GM|-80.97058|1.4132032182494703|82|1
35.03469|0d2e3c9f59fabf708d1ce4757b53ebb2bb699e2b|1.47|2014-09-28 19:18:00|1.4132775322775095|3|7203618340|82|0.6114706929155321|0|58|6152|-80.97058|1546|35.03469|BULB-HOUSEHOLD-PRIVATE LABEL|0.47|18|HT 60 WATT SOFT WHITE|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00072036183415|LIGHT BULBS/ELECTRICAL|GM|-80.97058|1.4132032182494703|82|1
35.03469|ac032bf2bc74f0b6cf68a43f49ec27f54d7d3ccc|0.97|2014-11-16 15:28:00|1.4132775322775095|3|7203698758|82|0.6114706929155321|0|58|31|-80.97058|4|35.03469|NON CARBONATED WATER|0.0|1|HT SPRING WATER|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00072036987587|BOTTLED WATER|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|3d920004ea55159ecebd999e4fedf743eeebee66|0.97|2014-11-14 20:38:00|1.4132775322775095|3|7203698758|82|0.6114706929155321|0|58|31|-80.97058|4|35.03469|NON CARBONATED WATER|0.0|1|HT SPRING WATER|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00072036987587|BOTTLED WATER|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|1e5678f881ac3813a335301ff57d2a47d2d7742a|0.97|2014-11-02 16:10:00|1.4132775322775095|3|7203698758|82|0.6114706929155321|0|58|31|-80.97058|4|35.03469|NON CARBONATED WATER|0.0|1|HT SPRING WATER|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00072036987587|BOTTLED WATER|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|b0560008d337685326f56020bc7a358e479bf659|0.97|2014-09-25 19:16:00|1.4132775322775095|3|7203698758|82|0.6114706929155321|0|58|31|-80.97058|4|35.03469|NON CARBONATED WATER|0.0|1|HT SPRING WATER|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00072036987587|BOTTLED WATER|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|400fb88aab27e5df927b78877dbcb8d6cf507cc6|0.97|2014-11-08 08:35:00|1.4132775322775095|3|7203698758|82|0.6114706929155321|0|58|31|-80.97058|4|35.03469|NON CARBONATED WATER|0.0|1|HT SPRING WATER|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00072036987587|BOTTLED WATER|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|d57c1570655d709ea8e58117b4b697369f659109|0.97|2014-12-31 19:19:00|1.4132775322775095|3|7203698758|82|0.6114706929155321|0|58|31|-80.97058|4|35.03469|NON CARBONATED WATER|0.0|1|HT SPRING WATER|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00072036987587|BOTTLED WATER|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|fd815c6e7f548328cd3edc6f707f7f568df23d35|0.97|2015-01-25 11:02:00|1.4132775322775095|3|7203698758|82|0.6114706929155321|0|58|31|-80.97058|4|35.03469|NON CARBONATED WATER|0.0|1|HT SPRING WATER|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00072036987587|BOTTLED WATER|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|ffbf3ce846346812b2951d9b17568ae54a8cd7ff|0.97|2015-02-15 14:07:00|1.4132775322775095|3|7203698758|82|0.6114706929155321|0|58|31|-80.97058|4|35.03469|NON CARBONATED WATER|0.0|1|HT SPRING WATER|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00072036987587|BOTTLED WATER|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|c8ea11cc0403153887146bde19c73cabde82fff8|0.97|2015-02-22 12:45:00|80.970593795509558|3|7203698758|82|35.038078856478108|0|4|31|-80.806073|4|35.106477|NON CARBONATED WATER|0.0|1|HT SPRING WATER|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|35.073829668338668|00072036987587|BOTTLED WATER|G1 GROCERY|-80.97058|80.970586164131277|4|1
35.03469|44965824fb4923010c7ffdabd1ba564640de7a32|0.97|2014-09-10 19:38:00|1.4132775322775095|3|7203698758|82|0.6114706929155321|0|58|31|-80.97058|4|35.03469|NON CARBONATED WATER|0.0|1|HT SPRING WATER|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00072036987587|BOTTLED WATER|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|2d6ecdef951102e5cb6dcb2b1e9ef721e9ed5d9a|0.97|2014-10-19 14:11:00|1.4132775322775095|3|7203698758|82|0.6114706929155321|0|58|31|-80.97058|4|35.03469|NON CARBONATED WATER|0.0|1|HT SPRING WATER|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00072036987587|BOTTLED WATER|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|23d40136e0096f1724800e3c3b2b9794c03928c1|7.99|2014-10-05 15:35:00|1.4132775322775095|3|3061300001|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|BROOKLYN LAGER 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00030613000012|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|663ea9b11b6c8e127c3cd1b86db1aa0c82e9d972|7.99|2014-09-14 18:35:00|1.4132775322775095|3|3061300001|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|BROOKLYN LAGER 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00030613000012|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|ab66bd5c30d17e8e25630eed65c59c097ba621b6|7.99|2014-10-01 19:53:00|1.4132775322775095|3|3061300001|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|BROOKLYN LAGER 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00030613000012|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|2e37548f16c31ad3f6bfa27c0414b97b5d0f349e|8.99|2014-11-06 18:48:00|1.4132775322775095|3|71280823275|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|HIGHLANDS KASHMIR 6PK IPA|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00712808232759|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|c608b63a1eefed963d72b318b026bc888343ac33|8.99|2014-10-31 18:43:00|1.4132775322775095|3|71280823275|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|HIGHLANDS KASHMIR 6PK IPA|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00712808232759|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|07ad63607e4c0a9192731ea33b2b1b8a9145fb20|8.99|2014-11-12 18:20:00|1.4132775322775095|3|3061300004|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|BROOKLYN BROWN 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00030613000043|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|7d87136d4af497e695528e31198b7c5a36f947d3|5.99|2015-01-05 19:49:00|1.4132775322775095|3|9522564910|82|0.6114706929155321|0|58|1288|-80.97058|379|35.03469|LOCAL MUFFINS|0.0|14|MODERN MUFFIN BANANA CHOC CHIP|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00095225649103|MUFFINS|BAKERY|-80.97058|1.4132032182494703|82|1
35.03469|dff06217e0957378221b6246705f5e05332c17d4|5.99|2014-12-28 16:42:00|1.4132775322775095|3|9522564910|82|0.6114706929155321|0|58|1288|-80.97058|379|35.03469|LOCAL MUFFINS|0.0|14|MODERN MUFFIN BANANA CHOC CHIP|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00095225649103|MUFFINS|BAKERY|-80.97058|1.4132032182494703|82|1
35.03469|2b61b35f418667092a32d7ca752247674f31945d|2.99|2014-10-17 19:23:00|1.4132775322775095|3|3680077038|82|0.6114706929155321|0|58|4828|-80.97058|1235|35.03469|ANTISEPTIC/DISINFECTANT|0.0|17|TC HAND SANITIZER ORIGINAL|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00036800174528|FIRST AID|HBC|-80.97058|1.4132032182494703|82|1
35.03469|b9bc75d79b3470c1191eff98e9e43d0abf268325|2.59|2014-09-19 19:54:00|1.4132775322775095|3|3700088179|82|0.6114706929155321|0|58|426|-80.97058|72|35.03469|NFS-PAPER TOWELS|0.0|1|BOUNTY TOWEL 1 RL SAS|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00037000881797|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|6bfe1fac44b0f5043fb82427d7ef427aed0acd1a|2.59|2014-12-20 17:40:00|1.4132775322775095|3|3700088179|82|0.6114706929155321|0|58|426|-80.97058|72|35.03469|NFS-PAPER TOWELS|0.59|1|BOUNTY TOWEL 1 RL SAS|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00037000881797|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|36595ae928d923a6e5ed8c84e6ac36cb3c5fe7d1|2.59|2015-02-28 16:43:00|1.4132775322775095|3|3700088179|82|0.6114706929155321|0|58|426|-80.97058|72|35.03469|NFS-PAPER TOWELS|0.59|1|BOUNTY TOWEL 1 RL SAS|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00037000881797|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.97058|1.4132032182494703|82|1
35.03469|4793f3415926dd32521f6598c7016bb8b2101ff4|9.99|2015-02-17 12:41:00|1.4132775322775095|3|75452700082|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|NEW BELGIUM SEASONAL 6PK NR|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00754527000820|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|2d2031e990cc8adb92ddbdab1fdca4d87b1636e9|9.99|2015-02-20 21:11:00|1.4132775322775095|3|75452700082|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|NEW BELGIUM SEASONAL 6PK NR|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00754527000820|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|2fedfa5a56f97acead8f74f71b9e76cdb5573ae9|9.99|2014-12-23 17:53:00|1.4132775322775095|3|71280812982|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|HIGHLAND GAELIC ALE 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00712808129820|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|26601ad793c690fbd613ec30a7d7324d9eb9b90b|8.99|2014-11-24 19:30:00|1.4132775322775095|3|71280812982|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|HIGHLAND GAELIC ALE 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00712808129820|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|8696330cd4a726342d209025793c8bfd3cf1d87a|8.99|2014-11-21 18:39:00|1.4132775322775095|3|71280812982|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|HIGHLAND GAELIC ALE 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00712808129820|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|6b1aeb231bada1293c7bfece99942af47c1ccd3c|9.99|2015-01-03 16:37:00|1.4132775322775095|3|71280812982|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|HIGHLAND GAELIC ALE 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00712808129820|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|46c8c2b799f1482cbcd8c6f234eeeb3a4a4467df|8.99|2014-12-01 16:49:00|1.4132775322775095|3|71280812982|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|HIGHLAND GAELIC ALE 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00712808129820|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|f9367fdd5abee442e80c12145a64bd22f1e23e6d|8.99|2014-12-12 19:03:00|1.4132775322775095|3|71280812982|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|HIGHLAND GAELIC ALE 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00712808129820|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|68083afff50eda05cc36d02f623aa6ef25e75e73|5.08|2014-12-24 14:59:00|1.4132775322775095|3||82|0.6114706929155321|0|58|523|-80.97058|64|35.03469|FRESH POTATOES|3.15|4|COO SWEET POTATOES, BULK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00204091000004|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|f6628b82bb35b937c3a653657b6a06dadd91659d|2.99|2015-01-17 17:19:00|80.970593795509558|3|7203670325|82|35.038078856478108|0|4|444|-80.806073|76|35.106477|NFS-PLASTIC WRAPS|0.0|1|YH PLASTIC WRAP|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|35.073829668338668|00072036703255|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.97058|80.970586164131277|4|1
35.03469|8a3c7ec548d5320491f3f5496fcb4dfd2ed7741d|7.99|2015-01-04 15:26:00|1.4132775322775095|3|8858640184|82|0.6114706929155321|0|58|9948|-80.97058|886|35.03469|NFS-PREM-CAB SAUVIGNON|0.0|13|COLUMBIA CREST GRAND EST CAB|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00088586401848|PREMIUM ($8-$10.99)|WINE|-80.97058|1.4132032182494703|82|1
35.03469|2f85f50abbcbde1cd619008e5b79be6e02843364|8.99|2014-12-03 18:57:00|1.4132775322775095|3|3410058878|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|LEINENKUGEL HOPPIN HELLES 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00034100588786|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|7cba15ee6d3d6f83c8f993eb5aaab8594fcca4fa|16.98|2014-12-27 15:10:00|1.4132775322775095|3|3410058878|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|LEINENKUGEL HOPPIN HELLES 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00034100588786|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|2
35.03469|8d1d640b292ff842fc44daa160f2b055af8756a3|16.98|2015-01-16 18:16:00|1.4132775322775095|3|3410058878|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|LEINENKUGEL HOPPIN HELLES 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00034100588786|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|2
35.03469|a4543d10b188ac21aa0813cd4997049b1c02dd99|8.99|2014-09-21 16:52:00|1.4132775322775095|3|3410058878|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|LEINENKUGEL HOPPIN HELLES 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00034100588786|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|2684cfc85abf69b61e20b50879c8d0b28a7599d9|8.99|2014-10-10 18:15:00|1.4132775322775095|3|3410058878|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|LEINENKUGEL HOPPIN HELLES 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00034100588786|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|1c1e79ddcd1b032816809cd862e6c8d153b159f2|8.99|2014-09-17 18:22:00|1.4132775322775095|3|3410058878|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|LEINENKUGEL HOPPIN HELLES 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00034100588786|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|abe839d1bb3144c7d0b5bce43aa85b2847348380|9.99|2014-10-22 18:46:00|1.4132775322775095|3|74052210016|82|0.6114706929155321|0|58|458|-80.97058|82|35.03469|CRAFT BEER|0.0|16|BELL'S SEASONAL 6PK|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00740522100160|DOMESTIC BEER|BEER|-80.97058|1.4132032182494703|82|1
35.03469|0874b12bfcef034a055aef0cb03ee945a68410f5|8.99|2015-03-03 19:00:00|1.4132775322775095|3|8858600134|82|0.6114706929155321|0|58|9948|-80.97058|886|35.03469|NFS-PREM-CAB SAUVIGNON|0.0|13|RED DIAMOND CABERNET SAUVIGNON|c77f4c64d2b97b308e2ce8b5df818825d76ac66a|0.23416205853811534|0.61177642288969325|00088586001345|PREMIUM ($8-$10.99)|WINE|-80.97058|1.4132032182494703|82|1
35.603432|4e956b714c39a60c25122f82a258b7908ddb0c35|1.83|2015-01-09 21:37:00|80.891462859624312|4||274|35.644742227944654|0|45|502|-80.85753|64|35.116638|FRESH BANANAS|0.0|4|BANANAS, YELLOW|c9829e5633564fc75a3a8e295c037f7d1af8761d|2.85447103820679|35.636605227883024|00204011000008|FRESH PRODUCE|PRODUCE|-80.895009|80.895257224699805|204|1
35.603432|3c3ba54624eaf57696552cba45ebcaea1ee3ce54|5.5|2014-11-01 16:40:00|80.891462859624312|4|2100065893|274|35.644742327619745|0|45|1441|-80.825175|274|35.152722|MAC AND CHEESE|0.0|1|KRAFT DELUXE DIN SHARP CHEDDAR|c9829e5633564fc75a3a8e295c037f7d1af8761d|2.85447103820679|35.636605227883024|00021000654932|PREP FOODS DINNERS|G1 GROCERY|-80.895009|80.895230702013905|160|2
35.603432|49dd5fc01cac004a67832070590dda0b6690ee99|4.89|2015-01-06 22:46:00|80.891462859624312|4|7313001237|274|35.644742227944654|0|45|1047|-80.85753|167|35.116638|PIZZA CRUST|0.0|7|BOBOLI ORIG PIZZA CRUST PP|c9829e5633564fc75a3a8e295c037f7d1af8761d|2.85447103820679|35.636605227883024|00073130012373|PITA/WRAPS/CRUST|COMMERCIAL BAKERY|-80.895009|80.895257224699805|204|1
35.603432|140ef455ea476e4a52614c6563d80c454e450694|2.49|2014-12-31 13:34:00|80.891462859624312|4|7096900102|274|35.644742327619745|0|45|543|-80.825175|64|35.152722|FRESH GARLIC|0.0|4|GARLIC IN OLIVE OIL, JAR|c9829e5633564fc75a3a8e295c037f7d1af8761d|2.85447103820679|35.636605227883024|00070969001028|FRESH PRODUCE|PRODUCE|-80.895009|80.895230702013905|160|1
35.603432|b111bbed80b02a51f4329984ee411aaf0ab22668|4.79|2015-01-07 17:57:00|80.891462859624312|4|7660656139|274|35.644742227944654|0|45|71|-80.85753|11|35.116638|GROC CONDIMENTS MARINADE|1.2|1|TROPICAL PEP SC MANGO COCONUT|c9829e5633564fc75a3a8e295c037f7d1af8761d|2.85447103820679|35.636605227883024|00076606561399|CONDIMENTS|G1 GROCERY|-80.895009|80.895257224699805|204|1
35.603432|5dcc50a0e6de4c09ee4244d06b8f8150f99c5006|5.69|2015-02-01 22:22:00|80.891462859624312|4|1740010667|274|35.644742227944654|0|45|239|-80.85753|38|35.116638|RICE-PACKAGED & BULK|0.0|1|MAHATMA RICE BASMATI 32OZ|c9829e5633564fc75a3a8e295c037f7d1af8761d|2.85447103820679|35.636605227883024|00017400106676|RICE GRAINS AND BEANS|G1 GROCERY|-80.895009|80.895257224699805|204|1
35.603432|1f8c26069992a7b9c1674c4ae0f799a65e5a71bd|4.19|2015-01-04 22:24:00|80.891462859624312|4|3800031846|274|35.644742227944654|0|45|74|-80.85753|9|35.116638|RTE CEREAL ALL FAMILY|0.0|1|KELL RICE KRISPIES 12|c9829e5633564fc75a3a8e295c037f7d1af8761d|2.85447103820679|35.636605227883024|00038000318467|CEREAL|G1 GROCERY|-80.895009|80.895257224699805|204|1
35.603432|66d63752e683f6ec20504ece884e47d7b687021d|3.99|2014-12-02 21:02:00|80.891462859624312|4|1111101215|274|35.644742324627551|0|45|429|-80.849471|73|35.161696|NFS-BAR SOAP|0.0|1|DOVE MEN EXTRA FRESH 2-BAR|c9829e5633564fc75a3a8e295c037f7d1af8761d|2.85447103820679|35.636605227883024|00011111012158|PERSONAL SOAP/BATH ADDITIVES|G1 GROCERY|-80.895009|80.895231544240062|35|1
35.603432|f3f36b6cf822bdb1f7878f632f61fea1c41e9e22|3.49|2014-12-24 14:46:00|80.891462859624312|4|7146426040|274|35.644742324627551|0|45|577|-80.849471|136|35.161696|OTHER MERCH FR MSC JUICE|0.0|4|BOLTHOUSE AMAZING MANGO|c9829e5633564fc75a3a8e295c037f7d1af8761d|2.85447103820679|35.636605227883024|00071464309503|OTHER MERCHANDISE|PRODUCE|-80.895009|80.895231544240062|35|1
35.603432|dc65ec173cb265860a3fcc1db5a350448485fab8|2.49|2014-11-04 20:36:00|80.891462859624312|4|70537200130|274|35.644742324627551|0|45|6821|-80.849471|1580|35.161696|J HOOK LAMI PROGRAM|0.0|18|SHELL SHINING COMBS|c9829e5633564fc75a3a8e295c037f7d1af8761d|2.85447103820679|35.636605227883024|00705372001302|J-HOOK|GM|-80.895009|80.895231544240062|35|1
35.603432|52ce53330bf35435c4de08f99ecd8e93aaf0b7da|1.57|2015-02-13 16:18:00|80.891462859624312|4||274|35.644742324627551|0|45|502|-80.849471|64|35.161696|FRESH BANANAS|0.0|4|BANANAS, YELLOW|c9829e5633564fc75a3a8e295c037f7d1af8761d|2.85447103820679|35.636605227883024|00204011000008|FRESH PRODUCE|PRODUCE|-80.895009|80.895231544240062|35|1
35.603432|fcfb739ece200664bb1e6c4672cc8a9b4f8222f4|3.99|2015-02-26 20:40:00|80.891462859624312|4|20980000000|274|35.644742227944654|0|45|1677|-80.85753|383|35.116638|INDIVIDUALS (PASTRY CASE)|0.0|14|MASCARPONE CUP/GLASS|c9829e5633564fc75a3a8e295c037f7d1af8761d|2.85447103820679|35.636605227883024|00209811000005|PASTRY CASE|BAKERY|-80.895009|80.895257224699805|204|1
35.603432|257995e1a0e567a0edfd07069a407078a5616285|2.5|2014-11-28 14:03:00|80.891462859624312|4|7203670856|274|35.644742324627551|0|45|427|-80.849471|72|35.161696|NFS-TOILET TISSUE|0.0|1|YH BATH 4 ROLL SS|c9829e5633564fc75a3a8e295c037f7d1af8761d|2.85447103820679|35.636605227883024|00072036708564|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.895009|80.895231544240062|35|1
35.603432|f88a2f078e6851bda183a05820091a7f4ce83331|2.19|2014-12-11 20:13:00|80.891462859624312|4|4900005010|274|35.644742324627551|0|45|55|-80.849471|8|35.161696|REGULAR|0.2|23|SPRITE  2 LITER|c9829e5633564fc75a3a8e295c037f7d1af8761d|2.85447103820679|35.636605227883024|00049000050158|CARBONATED BEVERAGES|BEVERAGE|-80.895009|80.895231544240062|35|1
35.603432|ae0e6fe344e94ca8a19b63ccb8148fdf1619ba79|14.99|2014-10-31 17:22:00|80.891462859624312|4|79837312125|274|35.644742324627551|0|45|458|-80.849471|82|35.161696|CRAFT BEER|0.0|16|MAGIC HAT THIS & THAT 12PK|c9829e5633564fc75a3a8e295c037f7d1af8761d|2.85447103820679|35.636605227883024|00798373121254|DOMESTIC BEER|BEER|-80.895009|80.895231544240062|35|1
35.603432|ca35e51a9fd6bdfc5d380fa4a6cbfdefad4ce559|2.79|2015-01-14 15:14:00|80.891462859624312|4|2740010307|274|35.644742327619745|0|45|313|-80.825175|51|35.152722|MARGARINE|0.0|3|COUNTRY CROCK SPREAD BOWL|c9829e5633564fc75a3a8e295c037f7d1af8761d|2.85447103820679|35.636605227883024|00027400103070|BUTTER & MARGARINE|DAIRY|-80.895009|80.895230702013905|160|1
35.603432|f2411c75feb5c90c9d438d752bbdee6b86e95e17|2.79|2015-01-28 17:25:00|80.891462859624312|4|2740010307|274|35.644742227944654|0|45|313|-80.85753|51|35.116638|MARGARINE|0.0|3|COUNTRY CROCK SPREAD BOWL|c9829e5633564fc75a3a8e295c037f7d1af8761d|2.85447103820679|35.636605227883024|00027400103070|BUTTER & MARGARINE|DAIRY|-80.895009|80.895257224699805|204|1
35.28326|2d1279d65ceb002788fb089651ed9bc3df24f1cd|1.59|2015-01-16 11:58:00|1.4094857484078087|1|20413500000|46|0.6158090578372145|0|26|500|-80.66939|64|35.28326|FRESH APPLES|0.16|4|GALA APPLES|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00891658001354|FRESH PRODUCE|PRODUCE|-80.66939|1.4079464610753885|46|1
35.28326|f630990bc9a73fd4bc3f81628cfec1d11a340c43|1.43|2015-01-04 09:55:00|1.4094857484078087|1|20413500000|46|0.6158090578372145|0|26|500|-80.66939|64|35.28326|FRESH APPLES|0.14|4|GALA APPLES|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00891658001354|FRESH PRODUCE|PRODUCE|-80.66939|1.4079464610753885|46|1
35.28326|6caf754544dcb1309cb7120cdac913a90de5bec2|1.97|2014-09-27 10:44:00|1.4094857484078087|1|7203656065|46|0.6158090578372145|0|26|315|-80.66939|52|35.28326|CHEESE-PROCESSED-SLICED|0.0|3|HT SINGLE WRAP CHEESE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036560650|CHEESE|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|c936d47202438ca1caa3ad71961a4ec412528c44|1.49|2015-01-05 11:10:00|1.4094857484078087|1|7203653022|46|0.6158090578372145|0|26|1273|-80.66939|50|35.28326|BAG VEG NON STEAM|0.5|5|HT WHOLE OKRA|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036537539|VEGETABLES-FROZEN|FROZEN|-80.66939|1.4079464610753885|46|1
35.28326|2374cc872bb20e096f4deab96307d0847c785be7|2.97|2014-12-01 13:32:00|1.4094857484078087|1|7203658035|46|0.6158090578372145|0|26|358|-80.66939|100|35.28326|REGULAR BACON|0.0|19|HT REGULAR SLICED BACON|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036580351|BACON|CASE READY MEATS|-80.66939|1.4079464610753885|46|1
35.28326|6702f4a64bd65ba4fb9175ee5fdda69e4038d257|5.94|2015-03-05 07:16:00|1.4094857484078087|1|7203658035|46|0.6158090578372145|0|26|358|-80.66939|100|35.28326|REGULAR BACON|0.0|19|HT REGULAR SLICED BACON|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036580351|BACON|CASE READY MEATS|-80.66939|1.4079464610753885|46|2
35.28326|c4e1dc125f1531a06761e7d729d26b119c134e15|2.98|2014-12-21 10:14:00|1.4094857484078087|1|7203653022|46|0.6158090578372145|0|26|1273|-80.66939|50|35.28326|BAG VEG NON STEAM|0.0|5|HT CALIFORNIA BLEND|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036535009|VEGETABLES-FROZEN|FROZEN|-80.66939|1.4079464610753885|46|2
35.28326|96b67dd6c3d7ffa844ee4f4b0e02ccca2a09799e|2.97|2015-02-16 12:24:00|1.4094857484078087|1|7203658035|46|0.6158090578372145|0|26|358|-80.66939|100|35.28326|REGULAR BACON|0.0|19|HT REGULAR SLICED BACON|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036580351|BACON|CASE READY MEATS|-80.66939|1.4079464610753885|46|1
35.28326|dbb5305eb7366f941b8c8ff60b64ab8f808107f9|3.49|2014-12-31 11:57:00|1.4094857484078087|1|85281048712|46|0.6158090578372145|0|26|330|-80.66939|55|35.28326|EGGS|0.0|3|LOL ALL NAT XL BROWN EGGS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00852810487126|EGGS FRESH|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|38583eebe718d049117988abd8820c8f2484248b|8.99|2015-02-15 15:20:00|1.4094857484078087|1|71280870122|46|0.6158090578372145|0|26|458|-80.66939|82|35.28326|CRAFT BEER|0.0|16|HIGHLAND SEASONAL 6PK|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00712808701224|DOMESTIC BEER|BEER|-80.66939|1.4079464610753885|46|1
35.28326|562d8f9834e5d66d5ae6c983fdbe366d6210e35a|1.89|2015-02-06 11:14:00|1.4094857484078087|1|64422572783|46|0.6158090578372145|0|26|4778|-80.66939|1230|35.28326|BARS-PROTEIN|0.3|17|POWER CRUNCH COOKIES N CRM BAR|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00644225727221|SPORTS NUTRITIONAL|HBC|-80.66939|1.4079464610753885|46|1
35.28326|9a21b2eed34e64b6a34420f67f948d542c6fc986|1.34|2014-10-07 15:51:00|1.4094857484078087|1|7203641111|46|0.6158090578372145|0|26|242|-80.66939|39|35.28326|CANNED BEANS|0.0|1|HT PEAS BLACKEYE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036411143|VEGETABLES-CAN/JAR|G1 GROCERY|-80.66939|1.4079464610753885|46|2
35.28326|8df1c5502fa80e396b40659e830d8699af635d00|1.34|2015-01-22 16:56:00|1.4094857484078087|1|7203641111|46|0.6158090578372145|0|26|242|-80.66939|39|35.28326|CANNED BEANS|0.0|1|HT PEAS BLACKEYE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036411143|VEGETABLES-CAN/JAR|G1 GROCERY|-80.66939|1.4079464610753885|46|2
35.28326|b467b8791c3329507bc9a4d4967eaf57a32924ae|1.49|2014-12-09 12:35:00|1.4094857484078087|1|7203653022|46|0.6158090578372145|0|26|1273|-80.66939|50|35.28326|BAG VEG NON STEAM|0.0|5|HT BABY BUD BROCCOLI FLORETS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036530790|VEGETABLES-FROZEN|FROZEN|-80.66939|1.4079464610753885|46|1
35.28326|072014b13cf458c382d09bfab15a02e9dc65222b|3.0|2014-09-15 12:20:00|1.4094857484078087|1|7203655029|46|0.6158090578372145|0|26|331|-80.66939|52|35.28326|NATURAL SLICED|1.0|3|HT MOZZARELLA SLICES|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036550293|CHEESE|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|2dd66261bf347d9ef6fafaf068f489920406038d|2.0100000000000002|2014-12-22 18:14:00|1.4094857484078087|1|7203641111|46|0.6158090578372145|0|26|242|-80.66939|39|35.28326|CANNED BEANS|0.24|1|HT PEAS BLACKEYE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036411143|VEGETABLES-CAN/JAR|G1 GROCERY|-80.66939|1.4079464610753885|46|3
35.28326|653dce53a80cb6c34801e69851f5666f41870a04|1.34|2014-12-08 15:56:00|1.4094857484078087|1|7203641111|46|0.6158090578372145|0|26|242|-80.66939|39|35.28326|CANNED BEANS|0.0|1|HT PEAS BLACKEYE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036411143|VEGETABLES-CAN/JAR|G1 GROCERY|-80.66939|1.4079464610753885|46|2
35.28326|e8450dc7e9086c22c4f458934a07a13867948497|1.34|2014-11-21 14:01:00|1.4094857484078087|1|7203641111|46|0.6158090578372145|0|26|242|-80.66939|39|35.28326|CANNED BEANS|0.0|1|HT PEAS BLACKEYE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036411143|VEGETABLES-CAN/JAR|G1 GROCERY|-80.66939|1.4079464610753885|46|2
35.28326|64200a96acfd8376cfdf46fbb294200a12d16969|2.69|2014-09-18 15:09:00|1.4094857484078087|1|7203663996|46|0.6158090578372145|0|26|342|-80.66939|57|35.28326|FRESH MILK|0.0|3|HARRIS TEETER 2%   MILK|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036639998|MILK|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|e603bc4df627ab434671d61570eeeff08e152397|2.69|2015-03-01 12:28:00|1.4094857484078087|1|70935100013|46|0.6158090578372145|0|26|556|-80.66939|64|35.28326|PACKAGED VEGETABLES|0.19|4|APIO BROCCOLI & CAULIFLOWER|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00709351000263|FRESH PRODUCE|PRODUCE|-80.66939|1.4079464610753885|46|1
35.28326|a4ce84b409c0764f01ee6ee01f8db203d21a9d93|2.69|2015-03-03 12:12:00|1.4094857484078087|1|70935100013|46|0.6158090578372145|0|26|556|-80.66939|64|35.28326|PACKAGED VEGETABLES|0.19|4|APIO BROCCOLI & CAULIFLOWER|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00709351000263|FRESH PRODUCE|PRODUCE|-80.66939|1.4079464610753885|46|1
35.28326|8d9c52785c7f481cd67731c8066dc2e2446ff201|1.89|2014-10-18 18:50:00|1.4094857484078087|1|73639310343|46|0.6158090578372145|0|26|247|-80.66939|39|35.28326|VEGETABLES-FLANKER|0.0|1|GLORY TURKEY SND TURNIP GREENS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00736393104239|VEGETABLES-CAN/JAR|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|d3fcf6b7f4ca69dae0aaa6dc36efa9d360ba20a5|5.67|2015-01-01 12:35:00|1.4094857484078087|1|73639310343|46|0.6158090578372145|0|26|247|-80.66939|39|35.28326|VEGETABLES-FLANKER|1.92|1|GLORY TURKEY SND TURNIP GREENS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00736393104239|VEGETABLES-CAN/JAR|G1 GROCERY|-80.66939|1.4079464610753885|46|3
35.28326|91f8cde83c8bf34a3ea5ba98229c7581f19887ec|3.25|2014-11-12 11:59:00|1.4094857484078087|1|7203656080|46|0.6158090578372145|0|26|318|-80.66939|52|35.28326|SHREDDED/GRATED CHEESE|0.0|3|HT FANCY SHRED MEXICAN CHEESE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036590442|CHEESE|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|8433b2633dcd348a19627e83deb50d1cd9e8ab6d|7.94|2015-02-15 18:49:00|80.66957994482128|1|7203658034|46|35.389569600311816|0|38|358|-80.762919|100|35.442529|REGULAR BACON|0.0|19|HT REGULAR SLICED BACON|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00072036580344|BACON|CASE READY MEATS|-80.66939|80.669550336401855|471|2
35.28326|347c54fc5371a89a8519e11f4f8889e22b503fe0|6.38|2014-10-11 13:49:00|1.4094857484078087|1|7271400222|46|0.6158090578372145|0|26|1473|-80.66939|278|35.28326|SWEET POTATOES|1.6|5|MCCAIN SW POT CROSS TRAX FRIES|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072714051210|FROZEN POTATO|FROZEN|-80.66939|1.4079464610753885|46|2
35.28326|815de577f62c2236bcc17990fc10cf8c9ef8f266|5.4|2014-10-09 16:42:00|1.4094857484078087|1|4144311023|46|0.6158090578372145|0|26|247|-80.66939|39|35.28326|VEGETABLES-FLANKER|1.4|1|M HOLMES SND LIMA BEANS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00041443119638|VEGETABLES-CAN/JAR|G1 GROCERY|-80.66939|1.4079464610753885|46|4
35.28326|e41eb485bd018838e92e20a77fbc8e3e13fd727a|3.69|2015-01-07 12:46:00|1.4094857484078087|1|4450034122|46|0.6158090578372145|0|26|357|-80.66939|104|35.28326|SMOKED SAUSAGE ROPES|0.0|19|HILLSHIRE TURKEY SMOKED SAUSAG|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00044500341157|DINNER SAUSAGE|CASE READY MEATS|-80.66939|1.4079464610753885|46|1
35.28326|ba4df808c14f38c9d1d5e3a786d37cef911fc056|2.99|2015-02-14 09:56:00|1.4094857484078087|1|3915310140|46|0.6158090578372145|0|26|214|-80.66939|33|35.28326|BROTH|0.0|1|RACHAEL RAY CHCK LOW SOD STOCK|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00039153101449|SOUP|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|dbf7e40f40a477ec5bdec47b6f1fcb538e32e250|3.39|2014-10-19 12:56:00|1.4094857484078087|1|4610000107|46|0.6158090578372145|0|26|331|-80.66939|52|35.28326|NATURAL SLICED|0.0|3|SARGENTO RF COBY JACK SLICES|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00046100001868|CHEESE|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|80cb9b97a0e605fd8a2640c39979f75f9c150ada|5.29|2015-03-02 07:15:00|1.4094857484078087|1|5150024177|46|0.6158090578372145|0|26|125|-80.66939|19|35.28326|PEANUT BUTTER|0.0|1|JIF CREAMY PEANUT BUTTER|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00051500241776|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|3bcc8b69eb779c32537bdcead4f656a9ce61fa59|5.29|2014-11-02 09:43:00|1.4094857484078087|1|5150024177|46|0.6158090578372145|0|26|125|-80.66939|19|35.28326|PEANUT BUTTER|1.3|1|JIF CREAMY PEANUT BUTTER|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00051500241776|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|40586d5123a3000fe45485766e1a1afd02fec8cd|5.29|2015-01-18 09:26:00|1.4094857484078087|1|5150024177|46|0.6158090578372145|0|26|125|-80.66939|19|35.28326|PEANUT BUTTER|0.0|1|JIF CREAMY PEANUT BUTTER|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00051500241776|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|c42b2bfc5f48f6c6bb62dc4f94210c67324da7b7|7.7|2015-01-18 09:27:00|1.4094857484078087|1|4812127620|46|0.6158090578372145|0|26|1037|-80.66939|164|35.28326|ENGLISH MUFFINS|1.92|7|THOMAS 100% WHEAT ENG MUFN PP|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00048121184070|BREAKFAST|COMMERCIAL BAKERY|-80.66939|1.4079464610753885|46|2
35.28326|77a31361d71205bb41b5567aec99f6bf6ee13ce4|2.99|2014-11-05 17:27:00|1.4094857484078087|1|4760001111|46|0.6158090578372145|0|26|1246|-80.66939|34|35.28326|SPICE BLENDS|0.0|1|WEBER ROASTED GARLIC & HERB|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00047600011074|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|69ed0f14460017c183aae8b92aef00f772c855cd|4.99|2014-09-27 10:43:00|1.4094857484078087|1|5150024177|46|0.6158090578372145|0|26|125|-80.66939|19|35.28326|PEANUT BUTTER|0.0|1|JIF CREAMY PEANUT BUTTER|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00051500241776|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|a86931c45f465ad1005bfad953a2a3f85dfc8050|3.69|2014-12-21 08:47:00|1.4094857484078087|1|2059300015|46|0.6158090578372145|0|26|1459|-80.66939|40|35.28326|FROZEN BISCUITS|0.0|5|MARY B'S BUTTERMILK BISCUIT|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00020593000157|FROZEN DOUGH|FROZEN|-80.66939|1.4079464610753885|46|1
35.28326|d427622071deb5c3320d246f2753997819f790fa|2.99|2015-01-28 09:31:00|80.66957994482128|1|85651300207|46|35.389569509311094|0|38|4778|-80.739|1230|35.141204|BARS-PROTEIN|1.0|17|NOGII HIGH PROTEIN BAR|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00856513002075|SPORTS NUTRITIONAL|HBC|-80.66939|80.669624056046359|171|1
35.28326|8664b1d8f1db2860fbb44e528f997433dc9a1014|2.99|2015-02-06 10:01:00|80.66957994482128|1|85651300207|46|35.389569509311094|0|38|4778|-80.739|1230|35.141204|BARS-PROTEIN|0.6|17|NOGII HIGH PROTEIN BAR|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00856513002075|SPORTS NUTRITIONAL|HBC|-80.66939|80.669624056046359|171|1
35.28326|4a923508659c872c6b08ffc810800f7b347729a5|3.35|2015-01-18 09:25:00|1.4094857484078087|1|1312000286|46|0.6158090578372145|0|26|1469|-80.66939|278|35.28326|REGULAR CUT FRIES|0.0|5|ORE-IDA MINI TATER TOTS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00013120000263|FROZEN POTATO|FROZEN|-80.66939|1.4079464610753885|46|1
35.28326|60666e536f3165d60d5d5221f6c2933d44b632ae|2.99|2015-01-18 10:51:00|80.66957994482128|1|85651300207|46|35.389569509311094|0|38|4778|-80.739|1230|35.141204|BARS-PROTEIN|1.0|17|NOGII HIGH PROTEIN BAR|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00856513002075|SPORTS NUTRITIONAL|HBC|-80.66939|80.669624056046359|171|1
35.28326|9f754787472d24a3d33f78c2955f0c645c3229c9|4.59|2014-11-14 17:24:00|1.4094857484078087|1|1340945132|46|0.6158090578372145|0|26|68|-80.66939|11|35.28326|BARBECUE SAUCES|0.6|1|SWEET BABY RAY 40 BBQ.|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00013409451328|CONDIMENTS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|d9076902df20c8348b81e73ded38b1ab6fb41e30|4.59|2015-02-04 12:37:00|1.4094857484078087|1|1340945132|46|0.6158090578372145|0|26|68|-80.66939|11|35.28326|BARBECUE SAUCES|0.0|1|SWEET BABY RAY 40 BBQ.|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00013409451328|CONDIMENTS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|7da232f1d2769960a73aa4228862b3569c5ba21b|2.99|2015-02-18 11:04:00|80.66957994482128|1|85651300207|46|35.389569509311094|0|38|4778|-80.739|1230|35.141204|BARS-PROTEIN|0.6|17|NOGII HIGH PROTEIN BAR|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00856513002075|SPORTS NUTRITIONAL|HBC|-80.66939|80.669624056046359|171|1
35.28326|26b747d51018ea54104d9a067395ac6d8cea5030|2.49|2014-09-29 17:03:00|1.4094857484078087|1|1410008550|46|0.6158090578372145|0|26|87|-80.66939|13|35.28326|CHEESE CRACKERS|0.0|1|PF GF FLAVOR BLAST PIZZA|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00014100085539|CRACKERS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|160c249620d81876a73fcbc97e89307f62c5486e|2.99|2015-01-16 10:42:00|80.66957994482128|1|85651300207|46|35.389569509311094|0|38|4778|-80.739|1230|35.141204|BARS-PROTEIN|1.0|17|NOGII HIGH PROTEIN BAR|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00856513002075|SPORTS NUTRITIONAL|HBC|-80.66939|80.669624056046359|171|1
35.28326|09d35e48650c4c2be9632b206294f194235b4991|2.99|2015-02-23 10:38:00|80.66957994482128|1|85651300207|46|35.389569509311094|0|38|4778|-80.739|1230|35.141204|BARS-PROTEIN|0.6|17|NOGII HIGH PROTEIN BAR|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00856513002075|SPORTS NUTRITIONAL|HBC|-80.66939|80.669624056046359|171|1
35.28326|3fb01b55316e9cdc8a1521b3c9d1c34684a8fa0c|1.78|2015-01-14 11:38:00|1.4094857484078087|1||46|0.6158090578372145|0|26|532|-80.66939|64|35.28326|FRESH CUCUMBERS|0.0|4|COO CUCUMBERS S/S|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00204062000002|FRESH PRODUCE|PRODUCE|-80.66939|1.4079464610753885|46|2
35.28326|0bdc62c9e2221e9cdd7e5a4545854b740ead108f|5.88|2014-11-24 12:36:00|1.4094857484078087|1|20543300000|46|0.6158090578372145|0|26|1832|-80.66939|415|35.28326|BH SLICING CHEESE|0.0|6|BOARS HEAD HAVARTI - JALAPENO|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00205433000003|SLICING CHEESE|DELI|-80.66939|1.4079464610753885|46|1
35.28326|91e87f36c0cfaef79fadd3dc0a6dc8cdb6ed7cea|4.75|2014-09-15 12:17:00|1.4094857484078087|1|20543300000|46|0.6158090578372145|0|26|1832|-80.66939|415|35.28326|BH SLICING CHEESE|0.0|6|BOARS HEAD HAVARTI - JALAPENO|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00205433000003|SLICING CHEESE|DELI|-80.66939|1.4079464610753885|46|1
35.28326|65b6a91d578be7cd3b7f665f1208895c2a45fc79|6.35|2014-11-17 11:36:00|80.66957994482128|1||46|35.389569509311094|0|38|503|-80.739|64|35.141204|FRESH GRAPES|0.91|4|GREEN GRAPES, SEEDLESS 12/16|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00204022000004|FRESH PRODUCE|PRODUCE|-80.66939|80.669624056046359|171|1
35.28326|eb3c9c88f159de46a6fefaf8faed76ff612ab9e4|4.39|2015-01-15 14:54:00|1.4094857484078087|1||46|0.6158090578372145|0|26|503|-80.66939|64|35.28326|FRESH GRAPES|0.22|4|GREEN GRAPES, SEEDLESS 12/16|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00204022000004|FRESH PRODUCE|PRODUCE|-80.66939|1.4079464610753885|46|1
35.28326|3978da13634f05d0714e8e266562c25b970418d1|10.38|2015-01-09 12:54:00|1.4094857484078087|1|80276308590|46|0.6158090578372145|0|26|118|-80.66939|17|35.28326|PRUNES|5.38|1|SUNSWEET PLUMS SNK 8PK|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00802763085900|FRUIT-DRIED|G1 GROCERY|-80.66939|1.4079464610753885|46|2
35.28326|23af9867cc890a426b12c798ee16135f3e9f6cba|1.99|2014-12-29 10:52:00|1.4094857484078087|1|2400016717|46|0.6158090578372145|0|26|115|-80.66939|16|35.28326|REMAINING FRUIT|0.32|1|DEL MONTE RED GRAPEFRUIT LS 15|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00733803103578|FRUIT-CAN/JAR|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|93c548f7abf3589aac820fbb813da1b75a24d040|2.49|2015-01-25 12:14:00|1.4094857484078087|1|61126999100|46|0.6158090578372145|0|26|97|-80.66939|8|35.28326|ENERGY DRINKS|0.49|23|CB RED BULL SUGAR FREE SINGLE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00611269101713|CARBONATED BEVERAGES|BEVERAGE|-80.66939|1.4079464610753885|46|1
35.28326|b33e1356278c4f00434e83440ab1f9dc090cec11|1.99|2015-02-12 16:37:00|1.4094857484078087|1|75606305414|46|0.6158090578372145|0|26|4926|-80.66939|1245|35.28326|EAR-EAR PLUGS|0.0|17|HEAROS ULT SOFTNESS EAR PLUGS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00756063054145|EYE & EAR CARE|HBC|-80.66939|1.4079464610753885|46|1
35.28326|aa1a0107eb0d15045685ed735a0366d60aee8bca|1.29|2015-02-09 11:58:00|1.4094857484078087|1|8379152001|46|0.6158090578372145|0|26|1981|-80.66939|480|35.28326|CHIPS|0.0|6|DIRTY POTATO CHIP SOUR CRM|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00083791520094|DRY GOODS|DELI|-80.66939|1.4079464610753885|46|1
35.28326|de3b8eef945b37384d36c43c24f3e8c5cfff9083|4.65|2015-03-05 12:10:00|1.4094857484078087|1|8000051306|46|0.6158090578372145|0|26|189|-80.66939|29|35.28326|TUNA-POUCH|0.8999999999999999|1|STARKIST TUNA PCH HICKORY SMKD|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00080000513069|SEAFOOD-CANNED|G1 GROCERY|-80.66939|1.4079464610753885|46|3
35.28326|e3b2a1d48fa66dea946f701c0317119a6eac2db4|1.79|2015-02-24 12:13:00|1.4094857484078087|1|1200000157|46|0.6158090578372145|0|26|31|-80.66939|4|35.28326|NON CARBONATED WATER|1.04|1|AQUAFINA WATER  1 LITER|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00012000001574|BOTTLED WATER|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|63c6959385e70d3393882fc89a749f4a2e786275|1.79|2015-01-13 12:58:00|1.4094857484078087|1|1200000157|46|0.6158090578372145|0|26|31|-80.66939|4|35.28326|NON CARBONATED WATER|1.04|1|AQUAFINA WATER  1 LITER|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00012000001574|BOTTLED WATER|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|5d3ea8120cbd868c5c1080f4fb04cd0e56300416|3.69|2014-12-29 10:54:00|1.4094857484078087|1|7203688073|46|0.6158090578372145|0|26|523|-80.66939|64|35.28326|FRESH POTATOES|0.0|4|HT BAKER POTATO 4 CT PKG|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036880734|FRESH PRODUCE|PRODUCE|-80.66939|1.4079464610753885|46|1
35.28326|99d55b7b29cea6185475d887024715723f205017|7.98|2014-09-25 17:43:00|1.4094857484078087|1|3760039885|46|0.6158090578372145|0|26|362|-80.66939|102|35.28326|PEPPERONIS|0.0|19|HORMEL PEPPERONI MINIS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00037600591829|LUNCHMEATS|CASE READY MEATS|-80.66939|1.4079464610753885|46|2
35.28326|efc1d98e76c94538bbd796d39557c47e4dcc96aa|2.89|2014-09-26 17:21:00|1.4094857484078087|1|3800040260|46|0.6158090578372145|0|26|1269|-80.66939|41|35.28326|BREAKFAST SYRUP CARRIER|0.0|5|EGGO BUTTERMILK WAFFLES|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00038000402906|BREAKFAST FOODS FROZEN|FROZEN|-80.66939|1.4079464610753885|46|1
35.28326|3edcdc846fa49dd5638af3e95eac057f1e143f31|3.99|2014-09-25 17:43:00|1.4094857484078087|1|3760039885|46|0.6158090578372145|0|26|362|-80.66939|102|35.28326|PEPPERONIS|0.0|19|HORMEL PEPPERONI MINIS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00037600591829|LUNCHMEATS|CASE READY MEATS|-80.66939|1.4079464610753885|46|1
35.28326|f9fa513a49af311acd0fcd10dfd9433745c9d215|3.35|2014-11-19 15:41:00|1.4094857484078087|1|1600042040|46|0.6158090578372145|0|26|13|-80.66939|2|35.28326|ROLLS/BISCUIT MIXES|0.0|1|BC BISQUICK|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00016000420403|BAKING MIXES|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|de8b4bedb3c9f7ae931ea11199f15ae5310c8fce|3.49|2014-11-17 12:07:00|1.4094857484078087|1|2840024053|46|0.6158090578372145|0|26|198|-80.66939|31|35.28326|CORN CHIPS|0.99|1|FRITOS BBQ|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00028400240543|SNACKS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|22b9e8daed43b42de07ce37ceef3fdca12573aaa|1.0|2014-11-18 17:14:00|1.4094857484078087|1|4000000435|46|0.6158090578372145|0|26|47|-80.66939|7|35.28326|REGISTER BARS|0.2|1|(FE)TWIX CARAMEL COOKIE BAR|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00040000004356|CANDY|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|341674fd519b0ae944728ac924e069a5c0043e22|15.49|2014-10-02 10:42:00|80.66957994482128|1|84105801560|46|35.389569509311094|0|38|3925|-80.739|1075|35.141204|RAZOR BLADES-MEN|0.0|17|HYDRO 5 SENS REFILL CARTRDG|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00841058015604|SHAVING NEEDS/MEN HAIR|HBC|-80.66939|80.669624056046359|171|1
35.28326|e080b4ba97d973548228f69eb34cb9408fc0372a|2.39|2014-12-21 10:13:00|1.4094857484078087|1|1480058223|46|0.6158090578372145|0|26|139|-80.66939|20|35.28326|REMAINING SHELF STABLE JUICES|0.0|1|REALEMON LEMON JUICE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00014800582239|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|09e4a35e7f8620f4fdd516b7a181cb1fc53795b4|5.19|2015-01-23 11:42:00|80.66957994482128|1|3700006222|46|35.389569590654133|0|38|4080|-80.810056|1080|35.219587|TOOTHPASTE-MULTI BENEFIT|1.7|17|CREST CMPLT+SCOPE X WH MNT BL|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00037000496311|ORAL HYGIENE|HBC|-80.66939|80.669559686082437|401|1
35.28326|70f4b149946a359acb638e214f13d9dea9c726f1|3.99|2014-11-15 09:57:00|1.4094857484078087|1|4163600020|46|0.6158090578372145|0|26|175|-80.66939|27|35.28326|CANNED MEATS|0.0|1|MRS FEARNOWS BRUNSWICK STEW|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00041636000200|PREPARED FOODS-RTS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|c73bb8d814a7c7cdc852090829c703eac236c2ca|11.45|2015-02-16 12:26:00|1.4094857484078087|1|4112907700|46|0.6158090578372145|0|26|1219|-80.66939|275|35.28326|PASTA SC CORE|0.0|1|CLASSICO SC ALFREDO 4 CHS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00041129274637|PASTA SAUCES|G1 GROCERY|-80.66939|1.4079464610753885|46|5
35.28326|542f4932f77a582698e103c9eb9687486d384944|4.99|2015-02-16 12:24:00|1.4094857484078087|1|4116701704|46|0.6158090578372145|0|26|4895|-80.66939|1240|35.28326|FOOT ODOR/WETNESS|0.0|17|GOLD BOND FOOT POWDER -01704|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00041167017043|FOOT CARE|HBC|-80.66939|1.4079464610753885|46|1
35.28326|4f99e8f06420bf5e0b573a8d7ed10c26c3d52096|3.75|2015-01-05 09:54:00|1.4094857484078087|1|4610000012|46|0.6158090578372145|0|26|318|-80.66939|52|35.28326|SHREDDED/GRATED CHEESE|1.25|3|SARGENTO OTB MONT JK FINE CUT|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00046100000182|CHEESE|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|859177019ea60e4ad7b79f50a1d0b789538f4f48|1.69|2015-01-13 12:58:00|1.4094857484078087|1|2840005509|46|0.6158090578372145|0|26|201|-80.66939|31|35.28326|POTATO CHIPS|0.0|1|LAYS STAX SALT&VINEGAR|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00028400055147|SNACKS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|62fee107d59ec7bd994359a85716a241c49fccc9|3.99|2014-10-21 11:06:00|80.66957994482128|1|7339001404|46|35.389569509311094|0|38|45|-80.739|7|35.141204|PEG GUM|2.0|1|MENTOS BUBBL FRSH COTTON CANDY|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00073390013684|CANDY|G1 GROCERY|-80.66939|80.669624056046359|171|1
35.28326|1f1ec698991276f8a0064d98c644e47e0c98d8ae|4.78|2014-11-03 12:13:00|1.4094857484078087|1|7084781116|46|0.6158090578372145|0|26|97|-80.66939|8|35.28326|ENERGY DRINKS|0.89|23|MONSTER ABSOLUTELY ZERO CAN|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00070847000037|CARBONATED BEVERAGES|BEVERAGE|-80.66939|1.4079464610753885|46|2
35.28326|24bdbef44560bb8821718c175e1b0182e46b5900|2.39|2015-01-22 16:50:00|1.4094857484078087|1|7084781116|46|0.6158090578372145|0|26|97|-80.66939|8|35.28326|ENERGY DRINKS|0.0|23|MONSTER ABSOLUTELY ZERO CAN|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00070847000037|CARBONATED BEVERAGES|BEVERAGE|-80.66939|1.4079464610753885|46|1
35.28326|d6887924c49ba2a2841c9ab4641f0cb2d72c22ab|3.99|2014-11-07 10:32:00|80.66957994482128|1|7339001404|46|35.389569509311094|0|38|45|-80.739|7|35.141204|PEG GUM|2.0|1|MENTOS BUBBL FRSH COTTON CANDY|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00073390013684|CANDY|G1 GROCERY|-80.66939|80.669624056046359|171|1
35.28326|ac0dcb2595b0a3c13fc45fc51186d420d6bc0c59|1.29|2014-11-13 11:57:00|1.4094857484078087|1|8379152001|46|0.6158090578372145|0|26|1981|-80.66939|480|35.28326|CHIPS|0.0|6|DIRTY POTATO CHIP BBQ|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00083791520049|DRY GOODS|DELI|-80.66939|1.4079464610753885|46|1
35.28326|40fdb8969905abfe3dbf8e9657ad2cb6fa04ce42|1.29|2015-02-10 12:20:00|1.4094857484078087|1|8379152001|46|0.6158090578372145|0|26|1981|-80.66939|480|35.28326|CHIPS|0.18|6|DIRTY POTATO CHIP BBQ|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00083791520049|DRY GOODS|DELI|-80.66939|1.4079464610753885|46|1
35.28326|be4de739d8b1388507ce06226d381a3209bda2cd|2.47|2014-10-13 17:44:00|1.4094857484078087|1|7203648998|46|0.6158090578372145|0|26|1460|-80.66939|40|35.28326|FROZEN BREAD AND ROLLS|0.0|5|HT  YEAST DINNER ROLLS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036489982|FROZEN DOUGH|FROZEN|-80.66939|1.4079464610753885|46|1
35.28326|0c81e35b656396ca5e71961ca9b6998817d6ee38|1.0|2015-02-13 15:52:00|1.4094857484078087|1||46|0.6158090578372145|0|26|565|-80.66939|64|35.28326|REDUCED PRODUCE|0.0|4|PRODUCE REWRAP BY CT|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00204845000007|FRESH PRODUCE|PRODUCE|-80.66939|1.4079464610753885|46|1
35.28326|81e9151f3a9c7662e2f0c50f554490b2cf43784f|2.0|2015-01-21 12:30:00|1.4094857484078087|1||46|0.6158090578372145|0|26|565|-80.66939|64|35.28326|REDUCED PRODUCE|0.0|4|PRODUCE REWRAP BY CT|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00204845000007|FRESH PRODUCE|PRODUCE|-80.66939|1.4079464610753885|46|2
35.28326|544a6f7c0367f6dbbbb0ce1981ff165e9ebfe85c|3.99|2015-01-05 09:53:00|1.4094857484078087|1|4157005982|46|0.6158090578372145|0|26|1148|-80.66939|21|35.28326|ALMONDS|0.5|1|BLUE DIAM HNY RST CHIPOTLE ALM|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00041570109847|NUTS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|7b3aefdeb0eb8c454c0a8e6d200f1f89292bf929|12.79|2015-01-31 10:11:00|1.4094857484078087|1|3700050963|46|0.6158090578372145|0|26|1513|-80.66939|66|35.28326|NFS-LAUNDRY DETERGENT PODS|0.0|1|TIDE PODS SPRING MEADOW 35CT|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00037000509639|DETERGENTS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|e8dae311f0aae55f3ebdc1c326dfa62f5c1f1ffa|1.49|2015-01-04 09:54:00|1.4094857484078087|1|3890000473|46|0.6158090578372145|0|26|115|-80.66939|16|35.28326|REMAINING FRUIT|0.0|1|DOLE PINEAPPLE 20 CHUNKS JC.|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00038900004736|FRUIT-CAN/JAR|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|695aad6e5b9ed77222cca4f211e01cfb8501d86c|2.99|2015-01-19 11:20:00|1.4094857484078087|1||46|0.6158090578372145|0|26|561|-80.66939|64|35.28326|FR PROD ORGANIC PRODUCE|0.0|4|ORG BUNCHED RED BEETS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00294539000000|FRESH PRODUCE|PRODUCE|-80.66939|1.4079464610753885|46|1
35.28326|63337ade1e0dca34443cfd1e706d3b6a4a51ee22|11.98|2015-02-14 16:43:00|80.66957994482128|1|20932700000|46|35.389569499749136|0|38|676|-80.605588|148|35.43259|TAILS|0.0|12|2PK LOBSTER TAILS 4.2 OZ MIN|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00209327000001|LOBSTERS|SEAFOOD|-80.66939|80.669630493766562|202|1
35.28326|7609c188805fcac2650f02db39120f1b3adae9c6|2.45|2015-03-02 16:12:00|80.66957994482128|1||46|35.389569509311094|0|38|500|-80.739|64|35.141204|FRESH APPLES|0.29|4|RED DEL APPLE, WA  48|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00233284000002|FRESH PRODUCE|PRODUCE|-80.66939|80.669624056046359|171|1
35.28326|c2b56734365a8b3184089db3cc1a6427dd2f5691|2.99|2015-02-04 12:38:00|1.4094857484078087|1|7680800149|46|0.6158090578372145|0|26|714|-80.66939|274|35.28326|MICROWAVE MEALS|0.0|1|BARILLA RTS SAUSAGE TOM ROTINI|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00076808004564|PREP FOODS DINNERS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|20ce8f3f7e3a7edcb65db5cd19d645f501368179|1.79|2014-10-12 09:22:00|1.4094857484078087|1|8079380770|46|0.6158090578372145|0|26|99|-80.66939|32|35.28326|LIQUID TEA|0.12|1|D FUZE SLENDER TROPICAL PUNCH|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00080793807765|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|227db9aa37f0c72faaea9dde2ff6177719492b20|2.59|2015-02-13 19:27:00|80.66957994482128|1|7080004600|46|35.389569600311816|0|38|361|-80.762919|105|35.442529|BREAKFAST SAUSAGE|0.6|19|JAMESTOWN MILD PORK SAUSAGE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00070800046003|BREAKFAST SAUSAGE|CASE READY MEATS|-80.66939|80.669550336401855|471|1
35.28326|81598fac5b17b2f837a845174d4c22267721ce28|6.98|2015-02-19 12:18:00|1.4094857484078087|1|2733100023|46|0.6158090578372145|0|26|495|-80.66939|108|35.28326|NON REFRIGERATED|1.98|19|LA BANDERITA L/CARB TORTILLAS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00027331000233|TORTILLAS|CASE READY MEATS|-80.66939|1.4079464610753885|46|2
35.28326|19debe484d399c05ecb63e25ec4637011389eef0|3.49|2015-02-07 12:50:00|1.4094857484078087|1|2733100023|46|0.6158090578372145|0|26|495|-80.66939|108|35.28326|NON REFRIGERATED|0.0|19|LA BANDERITA L/CARB TORTILLAS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00027331000233|TORTILLAS|CASE READY MEATS|-80.66939|1.4079464610753885|46|1
35.28326|167588d13cf24af01ff2e4a3c969f00cf7a0cf14|3.49|2015-02-26 12:18:00|1.4094857484078087|1|2733100023|46|0.6158090578372145|0|26|495|-80.66939|108|35.28326|NON REFRIGERATED|0.0|19|LA BANDERITA L/CARB TORTILLAS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00027331000233|TORTILLAS|CASE READY MEATS|-80.66939|1.4079464610753885|46|1
35.28326|c5120def1bca4f5ae4e007c9b582a275896062c0|3.49|2015-03-01 12:17:00|1.4094857484078087|1|2733100023|46|0.6158090578372145|0|26|495|-80.66939|108|35.28326|NON REFRIGERATED|0.0|19|LA BANDERITA L/CARB TORTILLAS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00027331000233|TORTILLAS|CASE READY MEATS|-80.66939|1.4079464610753885|46|1
35.28326|d1e33acdce670afac7a96c7f0bf92120b00bbb8a|3.49|2015-02-14 09:55:00|1.4094857484078087|1|2733100023|46|0.6158090578372145|0|26|495|-80.66939|108|35.28326|NON REFRIGERATED|0.0|19|LA BANDERITA L/CARB TORTILLAS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00027331000233|TORTILLAS|CASE READY MEATS|-80.66939|1.4079464610753885|46|1
35.28326|4571649d81bc7d6848cd9d7675586a2b8a5a786d|2.79|2015-02-02 11:33:00|1.4094857484078087|1|2100064353|46|0.6158090578372145|0|26|184|-80.66939|28|35.28326|SALAD DRESSINGS-LIQUID|0.79|1|KRAFT DRS RANCH 16|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00021000643615|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|ccd37c0099b36ff0c7adb40c007600bab0f7fd40|12.530000000000001|2014-10-17 14:27:00|1.4094857484078087|1|20328700000|46|0.6158090578372145|0|26|641|-80.66939|137|35.28326|PREMIUM PORK|0.0|2|PORK LOIN RIB END CHOPS BNLS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00203287000002|PORK|MEAT|-80.66939|1.4079464610753885|46|2
35.28326|d09048b8db20c1d3ab617511890b9f14aadd3681|8.15|2014-10-09 16:20:00|1.4094857484078087|1|20328700000|46|0.6158090578372145|0|26|641|-80.66939|137|35.28326|PREMIUM PORK|0.0|2|PORK LOIN RIB END CHOPS BNLS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00203287000002|PORK|MEAT|-80.66939|1.4079464610753885|46|1
35.28326|441dc4e750ad2c595c18caeac885cd996db3a4e9|1.49|2014-12-22 18:16:00|1.4094857484078087|1|7618316363|46|0.6158090578372145|0|26|99|-80.66939|32|35.28326|LIQUID TEA|0.5|1|SNAPPLE KIWI STRAWBERRY|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00076183163634|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|79afc16916a72626920d73420271972859dc22d2|4.39|2015-02-10 12:26:00|1.4094857484078087|1|1600027533|46|0.6158090578372145|0|26|81|-80.66939|9|35.28326|RTE CEREAL KIDS|1.89|1|GM GOLDEN GRAHAMS 16|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00016000275331|CEREAL|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|2c81334b038317deda40e2259ea83f58c9bb1ae1|7.99|2014-11-08 09:43:00|1.4094857484078087|1|79285056999|46|0.6158090578372145|0|26|3939|-80.66939|1075|35.28326|SHAVING CREAM MEN-CREAM|0.0|17|BURTS B SHAVE CREAM|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00792850569997|SHAVING NEEDS/MEN HAIR|HBC|-80.66939|1.4079464610753885|46|1
35.28326|41063e8165c3c7785c5334dd354765c60aafa229|6.99|2014-11-05 17:28:00|1.4094857484078087|1|7203698109|46|0.6158090578372145|0|26|252|-80.66939|45|35.28326|PREMIUM ICE CREAM|0.0|5|HT VANILLA 4QT PAIL IC|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036981097|ICE CREAM|FROZEN|-80.66939|1.4079464610753885|46|1
35.28326|dca956ced0b4fdb7501141a0a2f257aa0de008bc|2.29|2015-01-16 11:57:00|1.4094857484078087|1|85290900355|46|0.6158090578372145|0|26|1265|-80.66939|57|35.28326|ALMOND MILK|0.3|3|CALIFIA FRM CHOC ALM MLK W/PRO|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00852909003619|MILK|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|5ded83b6104d50bd20642c9e6e6be8360c5ab578|1.79|2014-12-08 15:57:00|1.4094857484078087|1|7339000393|46|0.6158090578372145|0|26|48|-80.66939|7|35.28326|REGISTER GUM|0.0|1|MENTOS FRSH SPEARMNT GUM 15CT|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00073390013875|CANDY|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|97e4180642c5bd07ea246f62b1791c2ff2635d50|4.99|2015-02-22 12:57:00|80.66957994482128|1|7203695649|46|35.389569600311816|0|38|1699|-80.762919|387|35.442529|EVERYDAY (COOKIES)|1.5|14|HT PINK SOFT SUGAR COOKIES|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00072036956491|COOKIES|BAKERY|-80.66939|80.669550336401855|471|1
35.28326|c19742c7cda21e1c50bf6d6bc630095c319d86db|1.79|2015-02-04 12:39:00|1.4094857484078087|1|7339000393|46|0.6158090578372145|0|26|48|-80.66939|7|35.28326|REGISTER GUM|0.0|1|MENTOS FRSH SPEARMNT GUM 15CT|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00073390013875|CANDY|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|3f3f8728a97cd2de785642b7cb13bb1307fef7a1|2.0|2015-01-26 11:49:00|80.66957994482128|1|4000000435|46|35.389569621679748|0|38|47|-80.746334|7|35.41832|REGISTER BARS|0.5|1|(FE)M&M PEANUT CANDY|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00040000000327|CANDY|G1 GROCERY|-80.66939|80.669527407304514|190|2
35.28326|db23016cdf36d4cedc9901f2ccf3f55630775d60|1.89|2014-11-12 12:00:00|1.4094857484078087|1|3800084496|46|0.6158090578372145|0|26|201|-80.66939|31|35.28326|POTATO CHIPS|0.0|1|PRINGLES CHEDDAR CHEESE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00038000844980|SNACKS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|ffc526043d5e3f6c669f701865748391d0b1db5c|3.99|2015-02-06 11:14:00|1.4094857484078087|1|9451441965|46|0.6158090578372145|0|26|389|-80.66939|66|35.28326|NFS-LAUNDRY DETERGENTS|0.0|1|XTRA DETERGENT MOUNTAIN RAIN|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00094514419656|DETERGENTS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|b6aff92c628c54d285bab459f74e489f389aa783|10.31|2014-12-09 12:40:00|1.4094857484078087|1|20598600000|46|0.6158090578372145|0|26|1800|-80.66939|400|35.28326|FFM BEEF|0.0|6|HT ROAST  BEEF|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00205986000000|FFM MEAT|DELI|-80.66939|1.4079464610753885|46|1
35.28326|c6733a324941bd046b4e52a97337b6487a7a2ee7|1.69|2014-11-26 19:40:00|1.4094857484078087|1|4900000044|46|0.6158090578372145|0|26|54|-80.66939|8|35.28326|DIET|0.0|23|CB COKE ZERO 20 OZ|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00049000040869|CARBONATED BEVERAGES|BEVERAGE|-80.66939|1.4079464610753885|46|1
35.28326|e510a39fa5b5fa8eb01db4242279ee9280bbf762|0.61|2014-11-13 12:09:00|1.4094857484078087|1||46|0.6158090578372145|0|26|502|-80.66939|64|35.28326|FRESH BANANAS|0.0|4|BANANAS, YELLOW|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00204011000008|FRESH PRODUCE|PRODUCE|-80.66939|1.4079464610753885|46|1
35.28326|7d5972bcecc45fd2790e1f843c1c44946d9d642b|5.55|2015-02-06 11:15:00|1.4094857484078087|1|3700006194|46|0.6158090578372145|0|26|3527|-80.66939|1045|35.28326|HAIR CARE SHPOO-MED|0.0|17|H&S REFRESH SHAMPOO NB|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00037000061984|HAIR & SCALP CARE|HBC|-80.66939|1.4079464610753885|46|1
35.28326|716c9c1490e08f5a175df87944a8e003a63e37d7|3.58|2014-11-03 12:14:00|1.4094857484078087|1|3940001614|46|0.6158090578372145|0|26|243|-80.66939|39|35.28326|BAKED BEANS|0.0|1|BUSH BKD BEAN HONEY 28|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00039400019855|VEGETABLES-CAN/JAR|G1 GROCERY|-80.66939|1.4079464610753885|46|2
35.28326|6db90c4908b5067ef73cbb6ab478e32b1f1cd542|3.58|2014-12-15 17:42:00|1.4094857484078087|1|3940001614|46|0.6158090578372145|0|26|243|-80.66939|39|35.28326|BAKED BEANS|0.0|1|BUSH GRL BEAN BOURBON|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00039400019107|VEGETABLES-CAN/JAR|G1 GROCERY|-80.66939|1.4079464610753885|46|2
35.28326|e0aa85f217687c22dfec0f7820c751944edd3473|1.38|2015-02-07 12:49:00|1.4094857484078087|1|71070842249|46|0.6158090578372145|0|26|580|-80.66939|136|35.28326|OTHER MERCH DRESSINGS|0.0|4|ORGANIC FF ITALIAN DRESSING|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00710708422492|OTHER MERCHANDISE|PRODUCE|-80.66939|1.4079464610753885|46|2
35.28326|75ec0f646bcc19b2e5671ce98f9a32b5304ecc71|4.99|2014-11-17 12:03:00|1.4094857484078087|1|4400004552|46|0.6158090578372145|0|26|92|-80.66939|13|35.28326|REMAINING CRACKERS|0.5|1|NABISCO EASY CHEESE SHARP|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00044000045531|CRACKERS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|671d970722eb629878529c0cd209db9a29d6b291|3.59|2014-12-11 09:34:00|1.4094857484078087|1|7353000003|46|0.6158090578372145|0|26|68|-80.66939|11|35.28326|BARBECUE SAUCES|0.0|1|CAROLINA TREET BBQ SAUCE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00073530000031|CONDIMENTS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|c45def3ba501aa0ee80ded84527714bfeed6dc53|2.58|2015-01-19 11:19:00|1.4094857484078087|1|4144311023|46|0.6158090578372145|0|26|247|-80.66939|39|35.28326|VEGETABLES-FLANKER|0.29|1|M HOLMES HOPPIN' JOHN|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00041443116330|VEGETABLES-CAN/JAR|G1 GROCERY|-80.66939|1.4079464610753885|46|2
35.28326|6991e364cdb04d7ea9c34167c9557c6a1767864b|6.99|2014-12-07 19:36:00|1.4094857484078087|1|4242122579|46|0.6158090578372145|0|26|358|-80.66939|100|35.28326|REGULAR BACON|1.5|19|BOARS HEAD SMOKED BACON 16 OZ|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00042421225792|BACON|CASE READY MEATS|-80.66939|1.4079464610753885|46|1
35.28326|a1e2a0a139825003c81eba6544277ce934cc4ffc|4.39|2015-03-07 12:58:00|80.66957994482128|1|3500068818|46|35.389569509311094|0|38|4056|-80.739|1080|35.141204|TOOTH BRUSH-PREMIUM|1.39|17|COLGATE 360 FULL MED TBRUSH|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00035000688187|ORAL HYGIENE|HBC|-80.66939|80.669624056046359|171|1
35.28326|ea78288e9ab02de742a1d29e42bb1b1cc2ed741f|6.99|2015-02-12 16:36:00|1.4094857484078087|1|4242122579|46|0.6158090578372145|0|26|358|-80.66939|100|35.28326|REGULAR BACON|1.0|19|BOARS HEAD SMOKED BACON 16 OZ|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00042421225792|BACON|CASE READY MEATS|-80.66939|1.4079464610753885|46|1
35.28326|ade63b5a5498c3f6059b2f3944bd81f3289e0270|6.99|2015-02-24 07:33:00|1.4094857484078087|1|4242122579|46|0.6158090578372145|0|26|358|-80.66939|100|35.28326|REGULAR BACON|1.0|19|BOARS HEAD SMOKED BACON 16 OZ|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00042421225792|BACON|CASE READY MEATS|-80.66939|1.4079464610753885|46|1
35.28326|338b158c8d249cf2f8502a1401372b169212b4d7|9.98|2014-12-10 17:11:00|1.4094857484078087|1|3500026859|46|0.6158090578372145|0|26|726|-80.66939|73|35.28326|NFS-BODY WASHES|2.49|1|GEAR 3 N 1 BODYWASH|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00035000268570|PERSONAL SOAP/BATH ADDITIVES|G1 GROCERY|-80.66939|1.4079464610753885|46|2
35.28326|5cb1a62a3ed25294f0e912eac26b06363b34f9c6|3.99|2014-11-21 14:00:00|1.4094857484078087|1|3010004911|46|0.6158090578372145|0|26|90|-80.66939|13|35.28326|SNACK CRACKERS|0.99|1|KEEBLER TOASTED WHEAT CRACKER|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00030100049111|CRACKERS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|bc4484f891302ece274dc3aa42e07ed680587d18|2.79|2015-02-02 17:27:00|1.4094857484078087|1|2740010307|46|0.6158090578372145|0|26|313|-80.66939|51|35.28326|MARGARINE|0.0|3|COUNTRY CROCK LIGHT|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00027400224027|BUTTER & MARGARINE|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|d998d20ea658e6081f97c16979fe370b7275fae7|3.99|2015-01-10 17:09:00|1.4094857484078087|1|3010004911|46|0.6158090578372145|0|26|90|-80.66939|13|35.28326|SNACK CRACKERS|0.0|1|KEEBLER TOASTED WHEAT CRACKER|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00030100049111|CRACKERS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|b2a2b353aa8e23f13981e519ff590869bd20e138|2.97|2014-11-02 09:42:00|1.4094857484078087|1|7203619046|46|0.6158090578372145|0|26|122|-80.66939|19|35.28326|HONEY|0.0|1|E  HT PURE HONEY BEAR|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036190468|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|ecff9414b2c45e8bad4992e8ac1dc60b51d53332|3.58|2014-12-01 10:08:00|80.66957994482128|1|5200033875|46|35.389569509311094|0|38|171|-80.739|20|35.141204|ISOTONIC DRINKS|0.82|1|GATORADE LEMON LIME|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00052000338775|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.66939|80.669624056046359|171|2
35.28326|19617c757c6a830408ff4684f764e5fcc1c20c8f|5.98|2014-11-29 15:08:00|1.4094857484078087|1|5100021232|46|0.6158090578372145|0|26|212|-80.66939|33|35.28326|CONDENSED SOUP|0.0|1|CAMP COND CREAM CHICKEN FAMILY|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00051000212436|SOUP|G1 GROCERY|-80.66939|1.4079464610753885|46|2
35.28326|34bea2bf61f0037f5950d50fc7f0fdfad5efda0b|3.38|2014-10-10 13:02:00|1.4094857484078087|1|5200033875|46|0.6158090578372145|0|26|171|-80.66939|20|35.28326|ISOTONIC DRINKS|0.62|1|GATORADE LEMON LIME|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00052000338775|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.66939|1.4079464610753885|46|2
35.28326|2acfbdd132037b64460aa4ebb1f118fa74624aba|1.89|2015-02-09 11:59:00|1.4094857484078087|1|3800084496|46|0.6158090578372145|0|26|201|-80.66939|31|35.28326|POTATO CHIPS|0.39|1|PRINGLES ORIGINAL|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00038000844966|SNACKS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|2520a41a75345fad02959ebb8fdbb080fd23fc69|1.89|2014-09-15 12:22:00|1.4094857484078087|1|3800084496|46|0.6158090578372145|0|26|201|-80.66939|31|35.28326|POTATO CHIPS|0.0|1|PRINGLES ORIGINAL|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00038000844966|SNACKS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|3467d58f957c8d0bffa1a0c6bc2adf2c9e7b8a66|1.69|2015-01-25 12:12:00|1.4094857484078087|1|4900000977|46|0.6158090578372145|0|26|31|-80.66939|4|35.28326|NON CARBONATED WATER|0.0|1|CB DASANI WATER 20 OZ SINGLES|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00049000009774|BOTTLED WATER|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|a2cfb17a2e2424ebb4b9075ac294f27be2c69e3e|1.69|2015-01-26 11:52:00|1.4094857484078087|1|4900000044|46|0.6158090578372145|0|26|55|-80.66939|8|35.28326|REGULAR|0.0|23|CB SPRITE PROPRIETARY 20 OZ|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00049000007640|CARBONATED BEVERAGES|BEVERAGE|-80.66939|1.4079464610753885|46|1
35.28326|7834457caf6a8a70699217a8403374e3d1b00c63|3.15|2014-10-12 09:23:00|1.4094857484078087|1|4300094511|46|0.6158090578372145|0|26|209|-80.66939|20|35.28326|POWDERED SOFT DRINKS|1.16|1|CRYSTAL LT OTG CHRY POMEGRANTE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00043000017289|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|5925b5867c04fe78fb6691eef947f5342f4a5cb8|1.69|2014-11-05 17:26:00|1.4094857484078087|1|4900000977|46|0.6158090578372145|0|26|31|-80.66939|4|35.28326|NON CARBONATED WATER|0.0|1|CB DASANI WATER 20 OZ SINGLES|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00049000009774|BOTTLED WATER|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|26c9595cea9e1d683cabce21d1a6e8dfa01245b2|1.69|2014-11-19 15:43:00|1.4094857484078087|1|4900000977|46|0.6158090578372145|0|26|31|-80.66939|4|35.28326|NON CARBONATED WATER|0.0|1|CB DASANI WATER 20 OZ SINGLES|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00049000009774|BOTTLED WATER|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|6fce0d3eb3c3c0dbc8d57a9331e9e71b3a6eebca|1.69|2015-02-02 11:19:00|1.4094857484078087|1|1200000129|46|0.6158090578372145|0|26|55|-80.66939|8|35.28326|REGULAR|0.0|23|CB DR PEPPER 20 OZ NR SINGLE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00078000082401|CARBONATED BEVERAGES|BEVERAGE|-80.66939|1.4079464610753885|46|1
35.28326|d7a7a5d392dd4e8551f20bfee06855e17329a749|5.69|2015-02-05 13:18:00|1.4094857484078087|1|5190001602|46|0.6158090578372145|0|26|839|-80.66939|102|35.28326|STACK PACKS|1.7|19|LOF PREMIUM HONEY TURKEY|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00051900016059|LUNCHMEATS|CASE READY MEATS|-80.66939|1.4079464610753885|46|1
35.28326|bd33cd139f66bc267c2032024afc60672cd625a1|2.75|2015-01-21 12:23:00|80.66957994482128|1|5150025537|46|35.389569600311816|0|38|125|-80.762919|19|35.442529|PEANUT BUTTER|0.75|1|JIF CREAMY PEANUT BUTTER|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00051500255162|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.66939|80.669550336401855|471|1
35.28326|f4534d0f90f276fd492abeda3933e203362f4473|6.29|2015-01-05 11:53:00|80.66957994482128|1|5150072001|46|35.389569600311816|0|38|125|-80.762919|19|35.442529|PEANUT BUTTER|0.0|1|JIF CREAMY PEANUT BUTTER|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00051500720011|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.66939|80.669550336401855|471|1
35.28326|90dc2ff2143f0994ed57c7d4657365868b5bef06|2.75|2015-02-13 15:49:00|1.4094857484078087|1|5150025537|46|0.6158090578372145|0|26|125|-80.66939|19|35.28326|PEANUT BUTTER|0.0|1|JIF CREAMY PEANUT BUTTER|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00051500255162|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|62ab3b4ea77c8ba742505eb2c96c6e2e08ddc1b2|3.99|2014-11-21 13:56:00|1.4094857484078087|1|7006601706|46|0.6158090578372145|0|26|3963|-80.66939|1075|35.28326|SHAVING NEEDS-OTHER|0.0|17|CLUBMAN MOUSTACHE WAX NEUTRAL|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00070066017069|SHAVING NEEDS/MEN HAIR|HBC|-80.66939|1.4079464610753885|46|1
35.28326|586da5456c5c4c2081f3c878ef30c34a3831bd20|0.69|2014-09-27 10:53:00|80.66957994482128|1|7203670022|46|35.389569509311094|0|38|4854|-80.739|1235|35.141204|HYDROGEN PEROXIDE|0.0|17|HT HYDROGEN PEROXIDE -70022|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00072036700223|FIRST AID|HBC|-80.66939|80.669624056046359|171|1
35.28326|6db8b8caf660ba76ebf0448fcdcf170676ba9a6a|1.47|2014-11-28 08:07:00|1.4094857484078087|1||46|0.6158090578372145|0|26|524|-80.66939|64|35.28326|FRESH PROD FRESH ONIONS|0.43|4|COO HONEY SWEET ONIONS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00204166000007|FRESH PRODUCE|PRODUCE|-80.66939|1.4079464610753885|46|1
35.28326|c42d30526470895eb0edbb008cf9adce14230f3d|3.98|2015-03-08 09:42:00|1.4094857484078087|1|4900004574|46|0.6158090578372145|0|26|171|-80.66939|20|35.28326|ISOTONIC DRINKS|2.4|1|POWERADE ZERO FRUIT PUNCH|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00049000056143|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.66939|1.4079464610753885|46|2
35.28326|c3d6f566e4b618615a091765fdf6f467c56a4b10|1.99|2015-02-24 12:13:00|1.4094857484078087|1|4900004574|46|0.6158090578372145|0|26|171|-80.66939|20|35.28326|ISOTONIC DRINKS|1.19|1|POWERADE ZERO FRUIT PUNCH|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00049000056143|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|a4ac154ec95e89915f6d2da87b8154aca7173ea5|3.98|2015-01-14 11:34:00|1.4094857484078087|1|4900004574|46|0.6158090578372145|0|26|171|-80.66939|20|35.28326|ISOTONIC DRINKS|0.74|1|POWERADE ZERO ORANGE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00049000054361|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.66939|1.4079464610753885|46|2
35.28326|3d827c37c908d3c01be70dbcf539c58e29cd8851|2.79|2015-01-31 10:14:00|1.4094857484078087|1|5210000245|46|0.6158090578372145|0|26|1246|-80.66939|34|35.28326|SPICE BLENDS|0.79|1|MC GRILL MATE SMOKEHOUSE MAPLE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00052100574110|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|3d77dc7fb4b68c404d155bf1d54796066dc35e78|4.29|2014-11-17 12:04:00|1.4094857484078087|1|4400002747|46|0.6158090578372145|0|26|91|-80.66939|13|35.28326|SPRAYED BUTTER CRACKERS|1.29|1|RTIZ HINT OF SALT|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00044000031190|CRACKERS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|4ea321a39c9808373d7041358548454dc35f3987|1.65|2015-01-04 09:55:00|1.4094857484078087|1||46|0.6158090578372145|0|26|500|-80.66939|64|35.28326|FRESH APPLES|0.0|4|GRANNY SMITH APPLES 72|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00204017000002|FRESH PRODUCE|PRODUCE|-80.66939|1.4079464610753885|46|1
35.28326|6ae87e12a8279e364dc26bc3c32da123f2a9ab96|8.49|2015-03-03 12:00:00|1.4094857484078087|1|2301200013|46|0.6158090578372145|0|26|1477|-80.66939|485|35.28326|SUSHI HYBRID|0.0|6|PLUS ROLL|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00023012000134|SUSHI|DELI|-80.66939|1.4079464610753885|46|1
35.28326|68e1ea3ca2ed76042adae3197a15ea1d974bfbab|8.49|2014-09-11 12:42:00|1.4094857484078087|1|2301200013|46|0.6158090578372145|0|26|1477|-80.66939|485|35.28326|SUSHI HYBRID|0.0|6|PLUS ROLL|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00023012000134|SUSHI|DELI|-80.66939|1.4079464610753885|46|1
35.28326|053c899b9e8388780889e3b949985b9878e72c97|8.49|2014-10-04 12:08:00|1.4094857484078087|1|2301200013|46|0.6158090578372145|0|26|1477|-80.66939|485|35.28326|SUSHI HYBRID|0.0|6|PLUS ROLL|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00023012000134|SUSHI|DELI|-80.66939|1.4079464610753885|46|1
35.28326|e3f2f9e651cec1610d3a7e834dedbe69f0440eb2|2.69|2014-12-29 10:51:00|1.4094857484078087|1|5000032822|46|0.6158090578372145|0|26|341|-80.66939|57|35.28326|CREAMERS|0.0|3|COFFEE-MATE SNICKERDOODLE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00050000904976|MILK|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|24e63285a07ace48e74a7d872c75762189c948f3|2.69|2014-12-10 17:09:00|1.4094857484078087|1|5000032822|46|0.6158090578372145|0|26|341|-80.66939|57|35.28326|CREAMERS|0.69|3|COFFEE-MATE SNICKERDOODLE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00050000904976|MILK|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|2e5b634b5dce7dae0d6a527d4adc508e693c4a17|4.99|2015-01-10 17:08:00|1.4094857484078087|1|2410044068|46|0.6158090578372145|0|26|87|-80.66939|13|35.28326|CHEESE CRACKERS|2.5|1|CHEEZ-IT PEPPERJACK|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00024100789252|CRACKERS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|08c4fd118e2fc8be69332589243796af669d00dd|4.29|2015-02-07 12:18:00|80.66957994482128|1|2840016014|46|35.389569600311816|0|38|201|-80.762919|31|35.442529|POTATO CHIPS|0.29|1|LAYS WAVY REGULAR|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00028400160209|SNACKS|G1 GROCERY|-80.66939|80.669550336401855|471|1
35.28326|f29eab10c8a8b19530e90b060f21e1bbe3a8f339|5.17|2015-01-25 12:13:00|1.4094857484078087|1||46|0.6158090578372145|0|26|561|-80.66939|64|35.28326|FR PROD ORGANIC PRODUCE|0.0|4|ORG GALA APPLES|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00294133000000|FRESH PRODUCE|PRODUCE|-80.66939|1.4079464610753885|46|1
35.28326|8567a431d7a7ae0b14d113d82cca7a8d21aec019|2.39|2014-09-18 15:11:00|1.4094857484078087|1|7084781116|46|0.6158090578372145|0|26|97|-80.66939|8|35.28326|ENERGY DRINKS|0.0|23|MONSTER LOW CARB ENRGY CAN|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00070847811268|CARBONATED BEVERAGES|BEVERAGE|-80.66939|1.4079464610753885|46|1
35.28326|7625af6d005076916b705345527a393d24ae5cf3|7.38|2015-03-05 12:10:00|1.4094857484078087|1|1340935231|46|0.6158090578372145|0|26|68|-80.66939|11|35.28326|BARBECUE SAUCES|1.85|1|SWEET BABY RAY 28 BBQ SC|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00013409352311|CONDIMENTS|G1 GROCERY|-80.66939|1.4079464610753885|46|2
35.28326|e6751321bdd4c9ff13868696f4ba6b346c7075e7|1.29|2014-12-08 15:56:00|1.4094857484078087|1|980000761|46|0.6158090578372145|0|26|48|-80.66939|7|35.28326|REGISTER GUM|0.0|1|(FE)TIC TAC FRUIT ADVENTURE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00009800007608|CANDY|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|75d03f5561a9d41b008b1b95af30d64c5a4a010d|4.99|2015-01-04 09:52:00|1.4094857484078087|1|1030054325|46|0.6158090578372145|0|26|1148|-80.66939|21|35.28326|ALMONDS|2.5|1|EMERALD 100 CAL WALNUT&ALMONDS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00010300543251|NUTS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|36f465ee5b590a09ad2dcd53ed5cfb199054cd8a|6.99|2015-03-06 12:35:00|80.66957994482128|1|1650053761|46|35.389569600311816|0|38|4236|-80.762919|1200|35.442529|DEX ADULT/CHILDREN|1.5|17|ALKA SELTZER COLD/COUGH 50592|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00016500537601|COUGH/COLD/SINUS|HBC|-80.66939|80.669550336401855|471|1
35.28326|ac91af02d5dd8d6dcd81452586f6eb577d13dc8b|4.29|2014-10-10 12:58:00|1.4094857484078087|1|3940001617|46|0.6158090578372145|0|26|243|-80.66939|39|35.28326|BAKED BEANS|0.0|1|BUSH BKD BEAN HOMESTYLE 55|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00039400016298|VEGETABLES-CAN/JAR|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|b193aec4792d5978ce4c791bac5aa6c2376b0708|2.85|2014-12-04 12:28:00|1.4094857484078087|1|4133500053|46|0.6158090578372145|0|26|184|-80.66939|28|35.28326|SALAD DRESSINGS-LIQUID|0.0|1|KENS DRS RANCH|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00041335332183|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|39cbd77422890c7da10258f7cc0473eb3934fb88|2.49|2014-09-27 19:37:00|1.4094857484078087|1|4410010755|46|0.6158090578372145|0|26|341|-80.66939|57|35.28326|CREAMERS|0.82|3|BAILEYS IRISH CREAM|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00044100107559|MILK|DAIRY|-80.66939|1.4079464610753885|46|1
35.28326|910a4d6957e499b9c68af0807d280e607f71a2d6|5.99|2014-09-18 15:10:00|1.4094857484078087|1|7164180174|46|0.6158090578372145|0|26|6604|-80.66939|1564|35.28326|DRY ERASE MARKER|0.0|18|EXPO LOW ODOR CHISEL 4CT|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00071641801745|SCHOOL & OFFICE SUPPLY|GM|-80.66939|1.4079464610753885|46|1
35.28326|49d55fba95e91d525658eda2c28a73ff3ce4855d|1.5|2015-01-29 11:50:00|80.66957994482128|1|7203641160|46|35.389569600311816|0|38|247|-80.762919|39|35.442529|VEGETABLES-FLANKER|0.0|1|HT GREEN BEANS ITALIAN CUT|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00072036411969|VEGETABLES-CAN/JAR|G1 GROCERY|-80.66939|80.669550336401855|471|2
35.28326|ba6f89ed40796fe3046372a73978af7bce10ddce|1.39|2014-11-24 12:38:00|1.4094857484078087|1|1254661959|46|0.6158090578372145|0|26|48|-80.66939|7|35.28326|REGISTER GUM|0.0|1|TRIDENT WATERMELON TWIST|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00012546615952|CANDY|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|e1c26c8b5b7fa4630ac9b629c43d24b759fd8abd|9.98|2014-12-31 11:56:00|1.4094857484078087|1|7203660022|46|0.6158090578372145|0|26|355|-80.66939|104|35.28326|FRESH GRILLING SAUSAGE|1.49|19|HT BRATWURST SAUSAGE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036600240|DINNER SAUSAGE|CASE READY MEATS|-80.66939|1.4079464610753885|46|2
35.28326|ac490887f9494b9ef10b1c9dcda6116fc990af09|2.69|2015-02-22 08:56:00|80.66957994482128|1|7203663217|46|35.389569509311094|0|38|330|-80.739|55|35.141204|EGGS|0.0|3|HT GRADE A LARGE EGGS 18 CT|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00072036632173|EGGS FRESH|DAIRY|-80.66939|80.669624056046359|171|1
35.28326|34f780805030eb304e6e7b607d26858fa200982e|2.38|2015-02-24 12:13:00|1.4094857484078087|1|7203653022|46|0.6158090578372145|0|26|1273|-80.66939|50|35.28326|BAG VEG NON STEAM|0.0|5|HT BRUSSEL SPROUTS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036531018|VEGETABLES-FROZEN|FROZEN|-80.66939|1.4079464610753885|46|2
35.28326|4d6602ce979015b4d89901e7cdc29fde98db2006|1.37|2014-10-11 13:49:00|1.4094857484078087|1|7203626061|46|0.6158090578372145|0|26|719|-80.66939|10|35.28326|NFS-COFFEE FILTERS|0.0|1|HT 12 CUP BASKET FILTERS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036260611|COFFEE|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|f3a52d6f5d807cfc7ce33981be1cc329e47e7c74|5.25|2014-12-11 11:09:00|80.66957994482128|1|7203633086|46|35.389569509311094|0|38|1148|-80.739|21|35.141204|ALMONDS|1.75|1|HT SMOKED ALMONDS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00072036330857|NUTS|G1 GROCERY|-80.66939|80.669624056046359|171|1
35.28326|518d3f0c4220e2b4fa1c767d0f3bbb6035cbfcb7|5.38|2015-02-07 06:29:00|1.4094857484078087|1|1450000253|46|0.6158090578372145|0|26|1272|-80.66939|50|35.28326|BAG VEG STEAM|1.34|5|BE STFRSH BROCC & CAULIF|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00014500011329|VEGETABLES-FROZEN|FROZEN|-80.66939|1.4079464610753885|46|2
35.28326|d1ffa020bad1ed5594fee25d7e41e3ed2f7a54d8|3.19|2015-03-08 09:42:00|1.4094857484078087|1|5100015339|46|0.6158090578372145|0|26|137|-80.66939|20|35.28326|TOMATO & VEGETABLE JUICE|0.0|1|V8 VEGGIE BLNDS-PURPLE POWER|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00051000217363|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|61544a6a184eb81b73fefd794d4dc65ae223b856|6.99|2015-03-05 12:08:00|1.4094857484078087|1|1200080994|46|0.6158090578372145|0|26|55|-80.66939|8|35.28326|REGULAR|3.5|23|DR. PEPPER FRIDGEMATE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00078000082166|CARBONATED BEVERAGES|BEVERAGE|-80.66939|1.4079464610753885|46|1
35.28326|9034e4fba4d33ac1608ea2d6339919e51016f941|1.79|2014-12-04 10:56:00|80.66957994482128|1|2830000089|46|35.389569453763507|0|38|1134|-80.825175|57|35.152722|CARTON MILK|0.0|3|SHAMROCK FARMS 2% CHOC MILK|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00028300003224|MILK|DAIRY|-80.66939|80.669659313048911|160|1
35.28326|fd6a7f7c473b47aa693532f6f5a57e2a248891b2|3.19|2014-11-15 09:57:00|1.4094857484078087|1|7203670212|46|0.6158090578372145|0|26|400|-80.66939|69|35.28326|NFS-LIQUID CLEANERS|0.0|1|YH PINE CLEANER|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036702128|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|10442cafdac720f36057ae317c58cfdb98f0c6c6|7.7|2015-01-02 12:02:00|1.4094857484078087|1|4812127620|46|0.6158090578372145|0|26|1037|-80.66939|164|35.28326|ENGLISH MUFFINS|1.93|7|THOMAS DBL PROTEINOATML EM PP|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00048121184032|BREAKFAST|COMMERCIAL BAKERY|-80.66939|1.4079464610753885|46|2
35.28326|bdc218a84fe9493b58b166158ab6570b727f4bd9|7.7|2015-01-02 12:01:00|1.4094857484078087|1|4812127620|46|0.6158090578372145|0|26|1037|-80.66939|164|35.28326|ENGLISH MUFFINS|1.93|7|THOMAS DBL PROTEINOATML EM PP|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00048121184032|BREAKFAST|COMMERCIAL BAKERY|-80.66939|1.4079464610753885|46|2
35.28326|47d040360085b556aa7900e8e149d8ddd2c4cb7b|4.99|2014-11-16 21:11:00|1.4094857484078087|1|5000031474|46|0.6158090578372145|0|26|144|-80.66939|229|35.28326|CEAMERS-POWDERED|0.0|1|COFFEE MATE CREAMY CHOCOLATE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00050000045952|COCOAS CREAMERS SYRUPS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|5f994f415e883a685e9b46c3a52dcacf2196b3ee|7.38|2014-09-27 19:36:00|1.4094857484078087|1|5000012734|46|0.6158090578372145|0|26|341|-80.66939|57|35.28326|CREAMERS|2.38|3|COFFEEMATE FRENCH VANILLA|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00050000322756|MILK|DAIRY|-80.66939|1.4079464610753885|46|2
35.28326|9f74f0ddeb75921c3aa94a0c4ac18c0304aef254|2.99|2015-01-21 18:05:00|1.4094857484078087|1|7084781310|46|0.6158090578372145|0|26|97|-80.66939|8|35.28326|ENERGY DRINKS|0.0|23|MONSTER VANILLA LIGHT CAN|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00070847813101|CARBONATED BEVERAGES|BEVERAGE|-80.66939|1.4079464610753885|46|1
35.28326|239539c98106bdf2acb0a6e7e28ad57fc0b88433|4.99|2015-01-12 11:52:00|1.4094857484078087|1|7885852039|46|0.6158090578372145|0|26|495|-80.66939|108|35.28326|NON REFRIGERATED|2.5|19|LA TORTILLA LOW CARB LARGE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00078858520391|TORTILLAS|CASE READY MEATS|-80.66939|1.4079464610753885|46|1
35.28326|cf1828333e746213dfafbb7e73fa898c099166c7|5.58|2015-02-15 17:08:00|1.4094857484078087|1|7110021162|46|0.6158090578372145|0|26|1439|-80.66939|274|35.28326|DRY DINNERS|0.0|1|HVR SOUTHWEST RANCH PAST SALAD|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00071100211627|PREP FOODS DINNERS|G1 GROCERY|-80.66939|1.4079464610753885|46|2
35.28326|6d1dbcd7321dcde31743e39fec69c5fbe46724c4|3.99|2015-02-11 13:21:00|80.66957994482128|1|7339001404|46|35.389569509311094|0|38|48|-80.739|7|35.141204|REGISTER GUM|1.99|1|MENTOS GUM MINT BOTTLE 50CT|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00073390014049|CANDY|G1 GROCERY|-80.66939|80.669624056046359|171|1
35.28326|9de5d2095e38e0667217ec840029f1997cb1e776|10.99|2014-11-08 09:43:00|1.4094857484078087|1|32586610506|46|0.6158090578372145|0|26|4335|-80.66939|1205|35.28326|NAPROXEN SODIUM|0.0|17|ALEVE ARTHRITIS CAPLET|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00325866536471|PAIN RELIEF|HBC|-80.66939|1.4079464610753885|46|1
35.28326|e14c4696da73584074995ed056ae780f91a94f8b|3.99|2014-12-14 18:32:00|1.4094857484078087|1|7778202983|46|0.6158090578372145|0|26|488|-80.66939|104|35.28326|SMOKED SAUSAGE LINKS|0.0|19|JOHNSONVILLE BETTER W/ CHEDDAR|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00077782023930|DINNER SAUSAGE|CASE READY MEATS|-80.66939|1.4079464610753885|46|1
35.28326|2027a9e08dd67a854129f782ffb8c098e238c262|5.69|2015-03-05 12:08:00|1.4094857484078087|1|7203633086|46|0.6158090578372145|0|26|1148|-80.66939|21|35.28326|ALMONDS|1.69|1|HT ROASTED & SALTED ALMONDS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036330864|NUTS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|b9126e50bed0e0ae199ea0b11bd8e1083c3a000c|5.0|2014-12-06 11:32:00|1.4094857484078087|1|7203670539|46|0.6158090578372145|0|26|164|-80.66939|39|35.28326|VEGETABLES-SPECIALTY|0.0|1|HT ASPARAGUS CUTS & TIPS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036705396|VEGETABLES-CAN/JAR|G1 GROCERY|-80.66939|1.4079464610753885|46|3
35.28326|50392f660cc11a1a9ff2af7e515b2f980f0872b8|4.29|2014-09-15 12:19:00|1.4094857484078087|1|4400003037|46|0.6158090578372145|0|26|90|-80.66939|13|35.28326|SNACK CRACKERS|1.29|1|WHEAT THINS RANCH|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00044000030421|CRACKERS|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|cbed3f06f5829a3515128e678b3ae46028a16793|7.99|2014-12-21 09:14:00|80.66957994482128|1|64786510001|46|35.389569509311094|0|38|4195|-80.739|1200|35.141204|COUGH & COLD REMEDY-ADULT|0.0|17|AIRBORNE CHEWABLE TABS BERRY|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00647865202219|COUGH/COLD/SINUS|HBC|-80.66939|80.669624056046359|171|1
35.28326|89aeeaebd1e81750f201831ed3ac9580edcab5b0|3.95|2014-12-10 17:11:00|1.4094857484078087|1|74816261452|46|0.6158090578372145|0|26|1460|-80.66939|40|35.28326|FROZEN BREAD AND ROLLS|1.45|5|SCHUBERTS PARKERHOUSE ROLLS|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00748162614528|FROZEN DOUGH|FROZEN|-80.66939|1.4079464610753885|46|1
35.28326|696196095291cd3165b438969a957e9d14d8a33e|1.89|2014-11-14 14:56:00|80.66957994482128|1||46|35.389569526736679|0|38|500|-80.80146|64|35.17739|FRESH APPLES|0.19|4|FUJI APPLES|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00204131000001|FRESH PRODUCE|PRODUCE|-80.66939|80.669611844116787|208|1
35.28326|9dadcf5eb6868e9c84bf010cf1a870ca82ca5595|13.69|2015-01-29 09:29:00|1.4094857484078087|1|20897500000|46|0.6158090578372145|0|26|977|-80.66939|201|35.28326|FRESH HT CHICKEN|6.86|2|FRESH BONELESS CHICKEN BREAST|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00208975000005|POULTRY|MEAT|-80.66939|1.4079464610753885|46|1
35.28326|1efca2623479be129a5633e15726743aed214fc6|1.69|2014-11-11 17:49:00|1.4094857484078087|1|1200000129|46|0.6158090578372145|0|26|55|-80.66939|8|35.28326|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.66939|1.4079464610753885|46|1
35.28326|3a920c89169c0e792a16a6a84fea71abf25f4510|1.69|2014-11-18 17:13:00|1.4094857484078087|1|1200000129|46|0.6158090578372145|0|26|55|-80.66939|8|35.28326|REGULAR|0.0|23|CB MTN DEW 20 OZ SINGLES|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00012000001314|CARBONATED BEVERAGES|BEVERAGE|-80.66939|1.4079464610753885|46|1
35.28326|1a60a738a85e17a79270864011d7a5c0d72f91e0|4.99|2014-10-26 10:23:00|80.66957994482128|1|2120097962|46|35.389569509311094|0|38|5607|-80.739|1512|35.141204|BRUSH-LINT|2.0|18|SCOTCH LINT ROLLER|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00021200979620|BROOMS/MOPS & BRUSHES|GM|-80.66939|80.669624056046359|171|1
35.28326|e8ed228ca805a0e5a051190e7036e666b51836d7|2.79|2015-02-02 11:33:00|1.4094857484078087|1|2100064353|46|0.6158090578372145|0|26|184|-80.66939|28|35.28326|SALAD DRESSINGS-LIQUID|0.79|1|KRAFT DRS ZESTY CATALINA|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00021000028276|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.66939|1.4079464610753885|46|1
35.28326|373aa675ecd95494a553603ce34c2ce30bd905f5|3.99|2015-01-07 12:46:00|1.4094857484078087|1|7778202983|46|0.6158090578372145|0|26|488|-80.66939|104|35.28326|SMOKED SAUSAGE LINKS|0.0|19|JOHNSONVILLE NO. ANDOUILLE|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00077782023954|DINNER SAUSAGE|CASE READY MEATS|-80.66939|1.4079464610753885|46|1
35.28326|8795ac37a5f09f8494f50525219ed113b6287990|2.29|2015-02-07 18:19:00|80.66957994482128|1|31254662920|46|35.389569600311816|0|38|4207|-80.762919|1200|35.442529|COUGH DROP-ADULT|0.0|17|HALLS PLUS CHERRY 62920|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00312546629202|COUGH/COLD/SINUS|HBC|-80.66939|80.669550336401855|471|1
35.28326|00882215204fe4b7c2a3fa083052a3f0cdcf90d9|3.29|2014-12-14 18:35:00|1.4094857484078087|1|7203644036|46|0.6158090578372145|0|26|273|-80.66939|43|35.28326|PREMIUM NOVELTIES|0.29|5|HT ICE CREAM SANDWICH-12PK|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|0.61471665291522548|00072036440365|FROZEN NOVELTIES|FROZEN|-80.66939|1.4079464610753885|46|1
35.28326|a1327b31cb0ba8582008eaeadea5b9ab57103dcd|3.99|2015-02-15 09:34:00|80.66957994482128|1|7203698196|46|35.389569587456172|0|38|276|-80.70901|45|35.17335|ICE MILK/SHERBET/YOGURT-FROZEN|0.99|5|HTT KEY LIME GRAHAM CRKR GEL|caeed762f127fd7d30f70fcf73f0b225cdc679f3|7.345742212861099|35.385064306269825|00072036981981|ICE CREAM|FROZEN|-80.66939|80.669562670511482|174|1
35.037115|7ad8352f2121218f94f90b41689b6fc62eb9d367|5.99|2014-10-19 12:53:00|80.805842308733688|1|4600029549|27|35.05573692327409|0|49|1213|-80.848528|272|35.053394|HISP DINNERS/SHELLS|0.0|1|OEP VAL PK KIT HARD SOFT|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00046000295497|HISPANIC PREP. FOODS|G1 GROCERY|-80.8062|80.806200491266651|11|1
35.037115|c57d3789d69f077fcbc3bfbe1c51be51040a3eec|1.69|2014-11-08 15:54:00|80.805842308733688|1|4600083251|27|35.055736922291381|0|49|1212|-80.770346|272|35.052812|HISP BEANS/PEPPERS|0.0|1|OEP CHILIES GREEN CHOPPED|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00046000832517|HISPANIC PREP. FOODS|G1 GROCERY|-80.8062|80.806207405918826|40|1
35.037115|ba38d979754c238e7d30584ee393be8506ae42d0|3.19|2015-01-04 18:32:00|80.805842308733688|1|4667501350|27|35.055736922602016|0|49|682|-80.850065|61|35.030252|KIDS|0.0|3|YOCRUNCH VAN/SNICKERS 4PK|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00046675013266|YOGURT|DAIRY|-80.8062|80.80620613079445|470|1
35.037115|0b3805263e14009284a0278701cea2710f6d044e|3.89|2014-09-17 14:22:00|80.805842308733688|1|4300095051|27|35.055736922291381|0|49|209|-80.770346|20|35.052812|POWDERED SOFT DRINKS|0.9|1|CRYSTAL LIGHT LEMONADE   12 QT|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00043000950654|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.8062|80.806207405918826|40|1
35.037115|39084dc82767901062b4cf4e0b2850920ee95497|3.89|2014-10-10 18:40:00|1.4091206135396188|1|4300095051|27|0.611513017149893|0|47|209|-80.8062|20|35.037115|POWDERED SOFT DRINKS|0.9|1|CRYSTAL LIGHT LEMONADE   12 QT|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|0.61242566243833529|00043000950654|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.8062|1.4103342460250419|27|1
35.037115|82459077b0e38b0c3207c66a57acf502377c1679|3.19|2015-01-02 19:57:00|80.805842308733688|1|4667501350|27|35.055736922602016|0|49|682|-80.850065|61|35.030252|KIDS|0.0|3|YOCRUNCH VAN/SNICKERS 4PK|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00046675013266|YOGURT|DAIRY|-80.8062|80.80620613079445|470|1
35.037115|9d01c28ce1b910e251300c6759ac6d7679907128|7.5|2015-01-05 15:56:00|80.805842308733688|1|4610000012|27|35.055736922338575|0|49|318|-80.847383|52|35.024464|SHREDDED/GRATED CHEESE|2.5|3|SARGENTO OTB TRAD 4 CHS MEX|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00046100011072|CHEESE|DAIRY|-80.8062|80.806207226728617|317|2
35.037115|f2aadba55d8c4a29c2aa50afb46149e47180f9dd|3.59|2014-10-13 15:47:00|80.805842308733688|1|4127100970|27|35.055736922602016|0|49|341|-80.850065|57|35.030252|CREAMERS|0.59|3|I/O ITNAT'L PUMPKIN PIE SPICE|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00041271009705|MILK|DAIRY|-80.8062|80.80620613079445|470|1
35.037115|87591e828b728a6727a5103a662741f67d88ca68|2.95|2015-03-02 15:32:00|80.805842308733688|1|3800012158|27|35.055736922937022|0|49|42|-80.816172|6|35.059823|GRANOLA/YOGURT BARS|0.45|1|SPECIAL K PASTRY STRAWBRY|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00038000490651|BREAKFAST FOODS|G1 GROCERY|-80.8062|80.806204355605288|66|1
35.037115|1539d160ac4331a57aa66dedd1fc004a8748ec1c|3.55|2015-02-22 13:44:00|80.805842308733688|1|3800039125|27|35.055736922937022|0|49|81|-80.816172|9|35.059823|RTE CEREAL KIDS|1.05|1|KELLOGG FROOT LOOPS 8.7|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00038000391255|CEREAL|G1 GROCERY|-80.8062|80.806204355605288|66|1
35.037115|c93048a29d39516ce3be75ac988748ed122443d8|5.79|2015-02-23 16:37:00|1.4091206135396188|1|1780015014|27|0.611513017149893|0|47|152|-80.8062|24|35.037115|NFS-CAT FOOD DRY|2.9|1|CAT CHOW INDOOR FORMULA|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|0.61242566243833529|00017800150187|PET FOOD/SUPPLIES|G1 GROCERY|-80.8062|1.4103342460250419|27|1
35.037115|9106ebb58cff0c346c9d81e274a9345f8bdc5a4b|3.99|2015-01-10 15:41:00|80.805842308733688|1|1906301228|27|35.055736922602016|0|49|31|-80.850065|4|35.030252|NON CARBONATED WATER|0.0|1|VYFINE FRUIT 2 O NAT GRAPE 6PK|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00019063012288|BOTTLED WATER|G1 GROCERY|-80.8062|80.80620613079445|470|1
35.037115|8c1948895eedd4a647080a96cbeed1c5d67fc19b|6.57|2014-10-05 10:37:00|80.805842308733688|1|2400016717|27|35.05573692327409|0|49|110|-80.848528|16|35.053394|FRUIT-CORE|1.57|1|DEL MONTE CHERRY MXD FRT LS.|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00024000019091|FRUIT-CAN/JAR|G1 GROCERY|-80.8062|80.806200491266651|11|3
35.037115|730b0bf325603b99fbdbd4746e2ab60cbdb45df7|1.29|2014-11-16 10:59:00|80.805842308733688|1|2200000899|27|35.05573692327409|0|49|48|-80.848528|7|35.053394|REGISTER GUM|0.0|1|EXTRA POLAR ICE 15 PC|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00022000008985|CANDY|G1 GROCERY|-80.8062|80.806200491266651|11|1
35.037115|ee367bfc457a377c8f7b5de69fa946498046d747|4.9|2014-09-10 18:30:00|80.805842308733688|1|1450000253|27|35.055736922291381|0|49|1272|-80.770346|50|35.052812|BAG VEG STEAM|1.23|5|BE STEAMFRESH GOLD/WHT CORN|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00014500012838|VEGETABLES-FROZEN|FROZEN|-80.8062|80.806207405918826|40|2
35.037115|7171f82bdb09721fa74ceb95295e80d339897d08|6.3|2015-01-24 15:52:00|80.805842308733688|1|2580002320|27|35.055736917200093|0|49|1271|-80.732725|41|35.082768|PROTEIN BREAKFAST|1.3|5|WW SMART ONES TRKY SAUS MUFFIN|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00025800026500|BREAKFAST FOODS FROZEN|FROZEN|-80.8062|80.806218378140883|147|2
35.037115|f3d05295a6b04fc689494fa0f8334f874e180d52|3.35|2015-01-26 15:48:00|80.805842308733688|1|2840005597|27|35.055736922602016|0|49|199|-80.850065|31|35.030252|DIPS & SALSAS|0.35|1|TOSTITOS RESTRNT  STYLE SALSA|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00028400089364|SNACKS|G1 GROCERY|-80.8062|80.80620613079445|470|1
35.037115|598c109dd34427431ad32a1fc53eb91c11728221|3.35|2014-12-29 17:33:00|80.805842308733688|1|2840005597|27|35.055736922602016|0|49|199|-80.850065|31|35.030252|DIPS & SALSAS|0.35|1|TOSTITOS RESTRNT  STYLE SALSA|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00028400089364|SNACKS|G1 GROCERY|-80.8062|80.80620613079445|470|1
35.037115|b2977c8613eaaf62962bb34103a14e0b399750a5|7.49|2014-10-26 12:05:00|1.4091206135396188|1|2840000288|27|0.611513017149893|0|47|205|-80.8062|31|35.037115|REMAINING SNACKS|0.5|1|FRITOLAY CLASSIC 20 CTN|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|0.61242566243833529|00028400002882|SNACKS|G1 GROCERY|-80.8062|1.4103342460250419|27|1
35.037115|f7c885687d7789932cbc4482bd9dc227f72c8f49|4.99|2015-02-04 19:04:00|80.805842308733688|1|2410044068|27|35.055736922291381|0|49|87|-80.770346|13|35.052812|CHEESE CRACKERS|2.5|1|CHEEZ-IT DUOZ CHEDDAR/PARMESAN|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00024100788958|CRACKERS|G1 GROCERY|-80.8062|80.806207405918826|40|1
35.037115|381c07990b91d50d36f98fe8987b75a09df861a6|2.59|2014-09-15 14:46:00|80.805842308733688|1|3620000250|27|35.055736922338575|0|49|1221|-80.847383|275|35.024464|PASTA SC VALUE|0.4|1|RAGU SC OWS WITH MEAT|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00036200003008|PASTA SAUCES|G1 GROCERY|-80.8062|80.806207226728617|317|1
35.037115|184d89808fda8ee151a1f574ae3ef3cbb645663d|5.18|2014-09-28 20:02:00|80.805842308733688|1|3620000250|27|35.055736921285323|0|49|1221|-80.771677|275|35.066546|PASTA SC VALUE|1.3|1|RAGU SC OWS WITH MEAT|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00036200003008|PASTA SAUCES|G1 GROCERY|-80.8062|80.806210523851107|45|2
35.037115|df12180dc72399ee9edc3d6a7692002b03c5bf9e|5.99|2015-01-07 14:25:00|80.805842308733688|1|7580582046|27|35.055736922338575|0|49|2021|-80.847383|505|35.024464|FRESH CHEESE|2.0|6|STELLA BLUE CHEESE CRUMBLES|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00075805820467|SPECIALTY CHEESE|DELI|-80.8062|80.806207226728617|317|1
35.037115|322fd6f3cddceca061c4aa1f9b7d76b50a77b80e|6.55|2014-12-05 17:50:00|1.4091206135396188|1|7570616502|27|0.611513017149893|0|47|254|-80.8062|892|35.037115|PREMIUM PIZZA|0.57|5|PALERMOS PEPPERONI PIZZA|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|0.61242566243833529|00075706165018|FROZEN PIZZA|FROZEN|-80.8062|1.4103342460250419|27|1
35.037115|618c9a11f1981def3ff26722af6a4fb04768ef15|0.87|2014-11-24 16:29:00|80.805842308733688|1|7203608080|27|35.055736922602016|0|49|120|-80.850065|15|35.030252|COATINGS & BREADERS|0.0|1|HT BREAD CRUMBS PLAIN|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00072036080806|FLOUR|G1 GROCERY|-80.8062|80.80620613079445|470|1
35.037115|a5dd57be62abd7e7e2ed7c6a09595c597f1332a2|1.69|2014-12-08 16:32:00|80.805842308733688|1|7203688003|27|35.055736922602016|0|49|527|-80.850065|64|35.030252|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00072036880031|FRESH PRODUCE|PRODUCE|-80.8062|80.80620613079445|470|1
35.037115|7a4ebb5b650d8c1b711ffe1e759cae00d86f9c45|1.69|2015-02-02 18:35:00|80.805842308733688|1|7203688003|27|35.055736922602016|0|49|527|-80.850065|64|35.030252|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00072036880031|FRESH PRODUCE|PRODUCE|-80.8062|80.80620613079445|470|1
35.037115|36f0a06e833058d82f12f6b8909003b2ab34628c|1.69|2015-01-25 12:25:00|80.805842308733688|1|7203688003|27|35.05573692327409|0|49|527|-80.848528|64|35.053394|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00072036880031|FRESH PRODUCE|PRODUCE|-80.8062|80.806200491266651|11|1
35.037115|7bb6e559e3e862187ea9b1a2ec39a0c5b1b976ca|1.69|2015-01-18 09:56:00|80.805842308733688|1|7203688003|27|35.05573692327409|0|49|527|-80.848528|64|35.053394|FRESH CARROTS|0.0|4|HT BABY CARROTS 1LB BAG|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00072036880031|FRESH PRODUCE|PRODUCE|-80.8062|80.806200491266651|11|1
35.037115|86ed17cb04e793d9d86f2e6caa77951c2a82c2f8|3.99|2014-11-23 15:46:00|80.805842308733688|1|7203697785|27|35.055736922338575|0|49|2022|-80.847383|505|35.024464|BLUE VEINED CHEESE|0.0|6|HT BLUE CHEESE CRMBLD|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00072036977854|SPECIALTY CHEESE|DELI|-80.8062|80.806207226728617|317|1
35.037115|7342e18f2cf065e7db927a105c388ca917617da0|10.19|2015-02-15 15:34:00|80.805842308733688|1|20596200000|27|35.055736922602016|0|49|1821|-80.850065|410|35.030252|BH TURKEY|1.02|6|BOARS HEAD MAPLE HONEY TURKEY|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00205962000000|BH MEAT|DELI|-80.8062|80.80620613079445|470|1
35.037115|605ca16566b5c0262324226a0cdc77a07f5ff0c2|9.99|2014-09-28 16:13:00|80.805842308733688|1|20596200000|27|35.055736922338575|0|49|1821|-80.847383|410|35.024464|BH TURKEY|1.0|6|BOARS HEAD MAPLE HONEY TURKEY|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00205962000000|BH MEAT|DELI|-80.8062|80.806207226728617|317|1
35.037115|688aca8e13840684911fc26911eaf33424da9cd3|17.45|2014-10-17 21:25:00|80.805842308733688|1|20138900000|27|35.055736922602016|0|49|296|-80.850065|49|35.030252|RANCHER BEEF|4.85|2|BEEF TENDERLOIN FILET MIGNON|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00201389000005|BEEF|MEAT|-80.8062|80.80620613079445|470|1
35.037115|9a3ba4cf29f618b541de35ee4e996ee7afbbbcf6|4.08|2015-02-01 17:19:00|80.805842308733688|1||27|35.05573692327409|0|49|500|-80.848528|64|35.053394|FRESH APPLES|0.0|4|RED DEL APPLE, WA  48|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00233284000002|FRESH PRODUCE|PRODUCE|-80.8062|80.806200491266651|11|1
35.037115|8fbae7317ed34b5546562458d4a2519dfc905553|6.49|2014-12-14 14:01:00|80.805842308733688|1|7430000071|27|35.055736922937022|0|49|5188|-80.816172|1305|35.059823|BABY OINTMENTS|0.0|17|DESITIN OINTMENT     -00071|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00074300000718|BABY HBC|HBC|-80.8062|80.806204355605288|66|1
35.037115|2a28680cecd31bb241616827708ad3a93603a9e2|5.98|2014-10-12 14:10:00|80.805842308733688|1|4470036113|27|35.055736922338575|0|49|659|-80.847383|103|35.024464|CHILDRENS LUNCH SNACKS|0.0|19|FUNPACK LUNCHABLE NACHO|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00044700006795|LUNCH SNACKS|CASE READY MEATS|-80.8062|80.806207226728617|317|2
35.037115|4a30cc6e2c61ab3214145d8e8e378baa6523fc56|8.99|2014-12-21 17:15:00|80.805842308733688|1|4242116030|27|35.055736917200093|0|49|1855|-80.732725|430|35.082768|BH SALAMI/CHUBBS|4.0|6|BH BIANCO D'ORO SALAME CHUBS|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00042421160307|SPECIALTY MEAT|DELI|-80.8062|80.806218378140883|147|1
35.037115|ac44674b2507b20abec65665ead519423dce6206|2.79|2015-03-09 18:28:00|80.805842308733688|1|3800035900|27|35.055736922338575|0|49|42|-80.847383|6|35.024464|GRANOLA/YOGURT BARS|0.29|1|KLG NUTRI GRN BAR FC APPLE COB|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00038000724145|BREAKFAST FOODS|G1 GROCERY|-80.8062|80.806207226728617|317|1
35.037115|90682993229c6e4c9fe621372aff0aa548135fd6|1.67|2014-09-21 12:12:00|80.805842308733688|1|4000029476|27|35.055736922937022|0|49|53|-80.816172|7|35.059823|THEATER BOX|0.0|1|M&M PLAIN THEATER BOX|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00040000294764|CANDY|G1 GROCERY|-80.8062|80.806204355605288|66|1
35.037115|aa95c835d075563b001f7ae842bcb202be724c4a|4.85|2014-12-24 17:37:00|80.805842308733688|1|7790011553|27|35.055736922291381|0|49|361|-80.770346|105|35.052812|BREAKFAST SAUSAGE|1.51|19|JIMMY DEAN MILD SAUSAGE|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00077900115530|BREAKFAST SAUSAGE|CASE READY MEATS|-80.8062|80.806207405918826|40|1
35.037115|760458e234c6ce5d59bbd3345dcac39a44c15959|14.97|2015-02-18 16:51:00|80.805842308733688|1|8136300100|27|35.055736922602016|0|49|1981|-80.850065|480|35.030252|CHIPS|8.97|6|NY STYLE SEA SALT BAGEL CHIPS|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00081363002009|DRY GOODS|DELI|-80.8062|80.80620613079445|470|3
35.037115|7fc7e628f08f472a1ad9d30d3ab22f6a49f81b4c|2.99|2014-09-26 18:48:00|1.4091206135396188|1|7203697784|27|0.611513017149893|0|47|2020|-80.8062|505|35.037115|CHEESE SPECIALTIES|0.0|6|HT FETA CHEESE CRMBLD|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|0.61242566243833529|00072036977847|SPECIALTY CHEESE|DELI|-80.8062|1.4103342460250419|27|1
35.037115|6cbb0e5e863f19fd3fede2bc71cf1789156ed5ea|5.99|2014-10-22 19:40:00|80.805842308733688|1|8143403135|27|35.055736922602016|0|49|9940|-80.850065|885|35.030252|NFS POP SYRAH/SHIRAZ|0.0|13|REX GOLIATH SHIRAZ|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00081434031358|POPULAR (4-$7.99)|WINE|-80.8062|80.80620613079445|470|1
35.037115|8145ff0bd75b016572d57ac6e1a0891df5b20ed1|5.99|2014-09-22 19:49:00|80.805842308733688|1|8143403130|27|35.055736922338575|0|49|9939|-80.847383|885|35.024464|NFS POP PINOT NOIR|0.0|13|REX GOLIATH PINOT NOIR|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00081434031303|POPULAR (4-$7.99)|WINE|-80.8062|80.806207226728617|317|1
35.037115|29a1adadc5d05bd0f3fb0da9d91c98293f87cf38|17.98|2014-12-01 21:27:00|1.4091206135396188|1|8500001227|27|0.611513017149893|0|47|9952|-80.8062|886|35.037115|NFS-PREM-PINOT NOIR|0.0|13|MIRASSOU PINOT NOIR|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|0.61242566243833529|00085000012277|PREMIUM ($8-$10.99)|WINE|-80.8062|1.4103342460250419|27|2
35.037115|ebe2a0e7933e9f92177050a671b941c325c7bee5|23.96|2015-02-13 16:30:00|80.805842308733688|1|8143403130|27|35.055736922291381|0|49|9939|-80.770346|885|35.052812|NFS POP PINOT NOIR|0.0|13|REX GOLIATH PINOT NOIR|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00081434031303|POPULAR (4-$7.99)|WINE|-80.8062|80.806207405918826|40|4
35.037115|804952ef487f55aceda525f95d332d6de62065f9|10.0|2014-10-15 18:27:00|80.805842308733688|1|8143403130|27|35.055736922291381|0|49|9939|-80.770346|885|35.052812|NFS POP PINOT NOIR|0.0|13|REX GOLIATH PINOT NOIR|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00081434031303|POPULAR (4-$7.99)|WINE|-80.8062|80.806207405918826|40|2
35.037115|c7ed1fef049f27d1acab29df8c06c3025a86cf75|2.99|2015-02-27 17:42:00|1.4091206135396188|1|70601011292|27|0.611513017149893|0|47|1219|-80.8062|275|35.037115|PASTA SC CORE|2.99|1|BARILLA SC TRADITIONAL.|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|0.61242566243833529|00076808003031|PASTA SAUCES|G1 GROCERY|-80.8062|1.4103342460250419|27|1
35.037115|1ad39e490e13fc08fbd00a7afe55c76de0c2cc1e|4.29|2014-10-11 22:33:00|1.4091206135396188|1|4900005235|27|0.611513017149893|0|47|55|-80.8062|8|35.037115|REGULAR|0.79|23|SEAGRAMS G' ALE 8PK 7.5 OZ CAN|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|0.61242566243833529|00072979004198|CARBONATED BEVERAGES|BEVERAGE|-80.8062|1.4103342460250419|27|1
35.037115|0a11d7acf776431aa97faac48737f2c83f6e19bb|2.29|2014-11-10 21:33:00|80.805842308733688|1|1900008501|27|35.055736921285323|0|49|50|-80.771677|7|35.066546|PEG CANDY|0.0|1|LIFE SAVERS GUMMIS 5 FLAVOR|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00019000083425|CANDY|G1 GROCERY|-80.8062|80.806210523851107|45|1
35.037115|e38c404d46cb0c2866c11904a2b12c02700e09d1|4.99|2014-10-27 16:29:00|80.805842308733688|1|85706300242|27|35.055736922602016|0|49|1218|-80.850065|273|35.030252|ASIAN OTHER|1.0|1|SAFFRON CHICKPEAS FALAFEL|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00857063002461|ASIAN PREP. FOODS|G1 GROCERY|-80.8062|80.80620613079445|470|1
35.037115|b8f1a5f9fa03a4a9f83ca6632ce8f3e6de0af7d3|5.99|2015-01-20 18:58:00|80.805842308733688|1|7203663044|27|35.055736922291381|0|49|974|-80.770346|201|35.052812|FRESH TURKEY|2.0|2|HT 93% LEAN GROUND TURKEY|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00072036630445|POULTRY|MEAT|-80.8062|80.806207405918826|40|1
35.037115|bf90c4c3405bd3ed4222cce834449b8c275afc2c|3.29|2014-11-11 18:59:00|80.805842308733688|1|1204403891|27|35.055736922291381|0|49|3876|-80.770346|1070|35.052812|SOLID-MALE|0.8|17|OLD SPICE HI ENDR PLAY MAKER|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00012044017906|DEODORANT|HBC|-80.8062|80.806207405918826|40|1
35.037115|307806d51464cf13c03a7901167e6da624aca20e|3.99|2015-01-08 19:54:00|80.805842308733688|1|7464100997|27|35.055736922937022|0|49|562|-80.816172|64|35.059823|FRESH CUT FRUIT|0.0|4|MULTIPACK APPLES & CARAMEL|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00074641009975|FRESH PRODUCE|PRODUCE|-80.8062|80.806204355605288|66|1
35.037115|f0284fb774d4e29525a399d24c1eee6b680b232f|4.39|2014-09-21 12:13:00|80.805842308733688|1|6843738350|27|35.055736922937022|0|49|46|-80.816172|7|35.059823|PKG CHOC|0.89|1|BROOKSDE POMEGRANATE|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00068437389082|CANDY|G1 GROCERY|-80.8062|80.806204355605288|66|1
35.037115|28194fa6767965cc360d7847437af0145dd78148|10.38|2014-10-12 18:59:00|1.4091206135396188|1|1204401560|27|0.611513017149893|0|47|3816|-80.8062|1070|35.037115|INVISIBLE-MALE|0.0|17|OLD SPICE FRSH COL AP/DEO FIJI|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|0.61242566243833529|00012044015605|DEODORANT|HBC|-80.8062|1.4103342460250419|27|2
35.037115|8a123dc5799fa6611e01aada6b00876201e8b745|9.99|2015-01-21 15:02:00|80.805842308733688|1|7203661016|27|35.055736922291381|0|49|297|-80.770346|49|35.052812|GROUND BEEF|1.52|2|GROUND CHUCK 80% LEAN 2 LB|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00072036610164|BEEF|MEAT|-80.8062|80.806207405918826|40|1
35.037115|5065ddb215d5677a196ce66bfeba04ca7d715cee|10.98|2014-12-14 12:53:00|80.805842308733688|1|1410009589|27|35.05573692327409|0|49|1255|-80.848528|13|35.053394|LUNCH BOX CRACKERS|0.0|1|PP PF MULTIPACK GOLDFISH CHEDR|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00014100095897|CRACKERS|G1 GROCERY|-80.8062|80.806200491266651|11|2
35.037115|60afa510b676acf2e89215ea6b061124608a0be6|3.99|2014-11-26 16:19:00|80.805842308733688|1|89504500026|27|35.055736922291381|0|49|3177|-80.770346|1010|35.052812|MAKE UP REMOVER|0.0|17|EXFOLIATING DLY CLNS TOWELETTE|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00895045000265|NAIL CARE|HBC|-80.8062|80.806207405918826|40|1
35.037115|2fff5844b7a8847a482ad4cb6b244e91f0301e8a|1.69|2014-10-15 12:31:00|80.805842308733688|1|4900000044|27|35.055736900681048|0|49|54|-80.826724|8|35.195689|DIET|0.0|23|CB DIET DR PEPPER 20OZ NR|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00078000083408|CARBONATED BEVERAGES|BEVERAGE|-80.8062|80.806235435475955|412|1
35.037115|11a5ef03bb1bd035fa87fc6b10722632d36e0386|1.69|2014-10-10 12:55:00|80.805842308733688|1|4900000044|27|35.055736900681048|0|49|54|-80.826724|8|35.195689|DIET|0.0|23|CB DIET DR PEPPER 20OZ NR|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00078000083408|CARBONATED BEVERAGES|BEVERAGE|-80.8062|80.806235435475955|412|1
35.037115|4f5cbcb2e55b506c8f977a2727039d446abd44a1|1.34|2014-11-18 18:40:00|80.805842308733688|1|7203624012|27|35.055736922291381|0|49|149|-80.770346|23|35.052812|WHSE PASTA CORE|0.0|1|HT PASTA ANGEL HAIR|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00072036240125|PASTA|G1 GROCERY|-80.8062|80.806207405918826|40|1
35.037115|d9e397e40b2dda6f1b3559188a3801493acde392|15.99|2015-02-17 17:19:00|80.805842308733688|1|2249480502|27|35.05573692327409|0|49|5867|-80.848528|1538|35.053394|CUTLERY|0.0|18|(PLR) THCK BEECHWD CHSE SLICR|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00022494805022|KITCHEN GADGETS|GM|-80.8062|80.806200491266651|11|1
35.037115|03d1e8cf4fee30e87f9ea850137df9cf956bb407|1.69|2014-12-15 11:17:00|80.805842308733688|1|1200000129|27|35.055736922937022|0|49|54|-80.816172|8|35.059823|DIET|0.0|23|CB DIET PEPSI 20 OZ NR|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00012000001307|CARBONATED BEVERAGES|BEVERAGE|-80.8062|80.806204355605288|66|1
35.037115|668a1dbd4d35d9887a5c6d2eac8b6c785b61f755|2.99|2014-10-06 12:12:00|80.805842308733688|1|7203601870|27|35.055736900681048|0|49|1895|-80.826724|450|35.195689|TEA|0.0|6|FFM RASPBERRY TEA|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00072036018755|BEVERAGES|DELI|-80.8062|80.806235435475955|412|1
35.037115|293fcdd11b39990cdce5174cab047e8a9d3bb58b|2.99|2014-09-26 12:19:00|80.805842308733688|1|7203601870|27|35.055736900681048|0|49|1895|-80.826724|450|35.195689|TEA|0.0|6|FFM RASPBERRY TEA|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00072036018755|BEVERAGES|DELI|-80.8062|80.806235435475955|412|1
35.037115|dcfda695b9334547a46b5f510d9f526c33c3198b|4.49|2014-09-17 13:37:00|80.805842308733688|1|2301290007|27|35.055736900681048|0|49|1483|-80.826724|485|35.195689|SUSHI ROLL AND WRAP|0.0|6|SUMMER ROLL|cb7ffbbf89cee48586a1658eacb9cf9760f3ad91|1.2867299282047586|35.053350220983141|00023012900076|SUSHI|DELI|-80.8062|80.806235435475955|412|1
35.204336|7db7e7ab46fa5bb010f4538b31b0a5c4b043be97|2.65|2015-01-07 12:38:00|80.843945456961976|4|4119691401|61|35.216652491781247|0|59|1201|-80.85013|33|35.175855|RTS CANNED|2.65|1|PROG RICH HRT CHCKEN WILD RICE|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|35.232478750868765|00041196453850|SOUP|G1 GROCERY|-80.844274|80.84427886456406|218|1
35.204336|4959fb937886bea9e2a68d3fb0d0d9c199ec9a13|2.29|2015-02-04 14:26:00|80.843945456961976|4|1450001098|61|35.216652491781247|0|59|1275|-80.85013|50|35.175855|BOX VEG|0.31|5|BE STEAMFRESH MIXED VEGES|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|35.232478750868765|00014500011282|VEGETABLES-FROZEN|FROZEN|-80.844274|80.84427886456406|218|1
35.204336|cb79d4a4ea738437a64b5fa984e28037e1afd7e1|11.59|2014-10-25 21:00:00|1.4094857484078087|4|20202100000|61|0.6144315741783704|0|26|299|-80.844274|49|35.204336|ANGUS BEEF|0.0|2|ANGUS BEEF THIN RIBEYE STEAK|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|0.61471665291522548|00202021000001|BEEF|MEAT|-80.844274|1.4109987626844462|61|1
35.204336|da9654ba7ce866358c9769c8deefb8c0418a143b|10.14|2014-10-11 15:08:00|80.843945456961976|4|20202100000|61|35.216652491781247|0|59|299|-80.85013|49|35.175855|ANGUS BEEF|3.5|2|ANGUS BEEF THIN RIBEYE STEAK|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|35.232478750868765|00202021000001|BEEF|MEAT|-80.844274|80.84427886456406|218|1
35.204336|1862d5f0973559fa52f09ef48ed302701bd60c80|1.95|2015-01-26 17:44:00|80.843945456961976|4||61|35.216652492421872|0|59|502|-80.826724|64|35.195689|FRESH BANANAS|0.0|4|BANANAS, YELLOW|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|35.232478750868765|00204011000008|FRESH PRODUCE|PRODUCE|-80.844274|80.844274157525618|412|1
35.204336|48bd76fe19c323a8d9683856a36e46691f5e2689|4.42|2014-11-11 19:17:00|80.843945456961976|4|2580002020|61|35.216652491781247|0|59|1278|-80.85013|48|35.175855|SINGLE SERVE NUTRITIONAL|0.0|5|WW SMART ONES CHICKN ENCHILADA|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|35.232478750868765|00025800019656|FROZEN MEALS|FROZEN|-80.844274|80.84427886456406|218|2
35.204336|a43fc7bf2a9a3e0e7f4abed52ba2e625dd73088b|5.49|2014-12-14 14:54:00|1.4094857484078087|4|20600100000|61|0.6144315741783704|0|26|1802|-80.844274|400|35.204336|FFM HAM|1.65|6|VIRGINIA BAKED HAM|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|0.61471665291522548|00206001000005|FFM MEAT|DELI|-80.844274|1.4109987626844462|61|1
35.204336|4e28555138bcf8d1c16bacb4f97e82ae7d2503ae|7.01|2014-09-20 12:15:00|1.4094857484078087|4|20039000000|61|0.6144315741783704|0|26|1801|-80.844274|400|35.204336|FFM TURKEY|1.56|6|HONEY SMOKED TURKEY BREAST|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|0.61471665291522548|00200397000007|FFM MEAT|DELI|-80.844274|1.4109987626844462|61|1
35.204336|7063d4c27895504d5ffbad254d5e731a7e171ef2|6.38|2014-09-28 10:09:00|80.843945456961976|4|20191900000|61|35.216652491781247|0|59|655|-80.85013|49|35.175855|STR MDE VALUE ADDED BEEF|0.71|2|SKEWERD BEEF KABOB W/VEGTABLES|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|35.232478750868765|00201919000000|BEEF|MEAT|-80.844274|80.84427886456406|218|1
35.204336|1e21404fdd21b08c427d721b6ec54e4f1296d216|5.49|2015-01-18 18:51:00|1.4094857484078087|4|20600200000|61|0.6144315741783704|0|26|1802|-80.844274|400|35.204336|FFM HAM|2.75|6|HONEY CURED HAM|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|0.61471665291522548|00206002000004|FFM MEAT|DELI|-80.844274|1.4109987626844462|61|1
35.204336|5e795108e3ecbb6f120afb2aa4ad86a46e7d682b|4.9|2014-12-04 21:09:00|80.843945456961976|4|20600200000|61|35.216652491781247|0|59|1802|-80.85013|400|35.175855|FFM HAM|2.45|6|HONEY CURED HAM|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|35.232478750868765|00206002000004|FFM MEAT|DELI|-80.844274|80.84427886456406|218|2
35.204336|891d3198dd91c7458a8997ce797afe5aae280ef8|4.17|2015-02-17 18:17:00|80.843945456961976|4|6414404551|61|35.216652491781247|0|59|179|-80.85013|27|35.175855|CANNED PASTA|1.47|1|CBRD WG ABC 123|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|35.232478750868765|00064144041350|PREPARED FOODS-RTS|G1 GROCERY|-80.844274|80.84427886456406|218|3
35.204336|5bb751649f9024485a171b230709206b4334c90d|2.69|2014-10-08 19:12:00|80.843945456961976|4|7203663996|61|35.216652491781247|0|59|342|-80.85013|57|35.175855|FRESH MILK|0.0|3|HARRIS TEETER 2%   MILK|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|35.232478750868765|00072036639998|MILK|DAIRY|-80.844274|80.84427886456406|218|1
35.204336|a0571e2bec5b7a210257a95ab721a4a4729e02ab|1.47|2015-02-01 15:24:00|1.4094857484078087|4|4142051960|61|0.6144315741783704|0|26|727|-80.844274|7|35.204336|SEASONAL CANDY-SINGLE FAC|0.72|1|I/O(V15)BRACH SM CONV HRT BX|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|0.61471665291522548|00041420519604|CANDY|G1 GROCERY|-80.844274|1.4109987626844462|61|3
35.204336|84e1e41433e12b1f188c63710beb8e12827dcb21|3.97|2014-12-14 15:00:00|1.4094857484078087|4|3040077377|61|0.6144315741783704|0|26|427|-80.844274|72|35.204336|NFS-TOILET TISSUE|0.0|1|ANGEL SOFT SOFT/STRONG 12DR|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|0.61471665291522548|00030400773778|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.844274|1.4109987626844462|61|1
35.204336|06e6a791f785b9b0c2547998c05c273233318d6e|1.69|2015-03-08 17:18:00|1.4094857484078087|4|2840005509|61|0.6144315741783704|0|26|201|-80.844274|31|35.204336|POTATO CHIPS|0.0|1|LAYS STAX CHEDDAR|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|0.61471665291522548|00028400055116|SNACKS|G1 GROCERY|-80.844274|1.4109987626844462|61|1
35.204336|52cf4264dd0ba2142725c4aea74cfa45a4a84569|5.99|2014-11-09 18:24:00|1.4094857484078087|4|7203688215|61|0.6144315741783704|0|26|500|-80.844274|64|35.204336|FRESH APPLES|1.02|4|HT GALA APPLE 5LB|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|0.61471665291522548|00072036882158|FRESH PRODUCE|PRODUCE|-80.844274|1.4109987626844462|61|1
35.204336|db1733b8a1b228dedd050550a6bdbd9d213f20f2|4.99|2015-02-16 17:51:00|1.4094857484078087|4|71575620002|61|0.6144315741783704|0|26|504|-80.844274|64|35.204336|FRESH BERRIES|2.5|4|STRAWBERRIES 1LB CLAM|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|0.61471665291522548|00846391005039|FRESH PRODUCE|PRODUCE|-80.844274|1.4109987626844462|61|1
35.204336|5d03be4a6035e6f86dfe95b3ef3352fb6942feec|13.58|2014-12-30 21:29:00|80.843945456961976|4|4900002890|61|35.216652450238506|0|59|54|-80.893784|8|35.478031|DIET|3.6|23|DT SPRITE ZERO 12PK FRIDGEPKCN|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|35.232478750868765|00049000037111|CARBONATED BEVERAGES|BEVERAGE|-80.844274|80.844313453841011|179|2
35.204336|6f81ae160a44baa359248a65e5801088e2bf4a9a|2.39|2015-02-28 10:01:00|80.843945456961976|4|7357013000|61|35.216652488252173|0|59|1267|-80.824767|53|35.116751|DIPS AND SPREADS|1.2|3|HELUVA GOOD FRENCH ONION DIP|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|35.232478750868765|00073570130002|CULTURES|DAIRY|-80.844274|80.844286405166315|294|1
35.204336|4ed7e7cae44f1e6739cbbfb1f23f7469eddf57d5|12.0|2014-11-19 18:21:00|80.843945456961976|4|66440177739|61|35.216652491781247|0|59|1165|-80.85013|87|35.175855|NFS-FRESH CONSUMER BUNCH|0.0|9|BUNCH- JUMBO SUNFLOWER 3 ST|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|35.232478750868765|00664401777390|FLORAL|FLORAL|-80.844274|80.84427886456406|218|3
35.204336|18ef59f568410fad7a503adaddbe5e8c31f28471|4.29|2014-11-06 17:17:00|1.4094857484078087|4|70897111899|61|0.6144315741783704|0|26|1703|-80.844274|387|35.204336|SEASONAL COOKIES|0.8|14|HARVEST ORANGE FRSTD SGR COOK|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|0.61471665291522548|00708971118990|COOKIES|BAKERY|-80.844274|1.4109987626844462|61|1
35.204336|7d1caafd45088dbe9e09426a3aa026204009b775|3.6|2014-10-05 17:12:00|80.843945456961976|4||61|35.216652492421872|0|59|531|-80.826724|64|35.195689|FRESH CORN|0.0|4|COO WHITE CORN|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|35.232478750868765|00204077000004|FRESH PRODUCE|PRODUCE|-80.844274|80.844274157525618|412|6
35.204336|16cd1a11ccbefcb6676477ebe6258d9b9d93f026|3.29|2015-01-17 16:59:00|1.4094857484078087|4|2840004768|61|0.6144315741783704|0|26|202|-80.844274|31|35.204336|PRETZELS|1.65|1|ROLD GOLD PRETZEL TINY TWIST|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|0.61471665291522548|00028400047685|SNACKS|G1 GROCERY|-80.844274|1.4109987626844462|61|1
35.204336|4a9e248e7fe11ebab82de9c2442f2da9e8d728f6|3.99|2014-11-05 14:06:00|80.843945456961976|4|4812121657|61|35.216652491781247|0|59|1036|-80.85013|164|35.175855|BREAKFAST BAGELS|2.0|7|THOMAS BLUBRY MINI  BGLS PP|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|35.232478750868765|00048121216764|BREAKFAST|COMMERCIAL BAKERY|-80.844274|80.84427886456406|218|1
35.204336|0c1c54cc135d46169858ac3650a92791e064c749|9.98|2014-09-21 18:12:00|80.843945456961976|4|2301290130|61|35.216652491781247|0|59|1477|-80.85013|485|35.175855|SUSHI HYBRID|0.0|6|CALIFORNIA ROLL SP|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|35.232478750868765|00023012901301|SUSHI|DELI|-80.844274|80.84427886456406|218|2
35.204336|43b2bb0135392f68dc4751df20b6ca20b466964b|4.99|2015-01-21 18:11:00|80.843945456961976|4|2301290130|61|35.216652491781247|0|59|1477|-80.85013|485|35.175855|SUSHI HYBRID|0.0|6|CALIFORNIA ROLL SP|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|35.232478750868765|00023012901301|SUSHI|DELI|-80.844274|80.84427886456406|218|1
35.204336|ed106a39e474ca579b63ab369e8eb56f3ab1439d|9.98|2014-12-22 17:20:00|1.4094857484078087|4|2301290130|61|0.6144315741783704|0|26|1477|-80.844274|485|35.204336|SUSHI HYBRID|0.0|6|CALIFORNIA ROLL SP|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|0.61471665291522548|00023012901301|SUSHI|DELI|-80.844274|1.4109987626844462|61|2
35.204336|9543e373b8b759d50a9a6829ba630dee04220c91|7.35|2015-02-15 18:08:00|80.843945456961976|4|4470002268|61|35.216652491781247|0|59|358|-80.85013|100|35.175855|REGULAR BACON|3.68|19|OSCAR MAYER THICK SLIC BACON|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|35.232478750868765|00044700019900|BACON|CASE READY MEATS|-80.844274|80.84427886456406|218|1
35.204336|a6a06aee0203a512d31354734b8f6059140984b0|6.99|2014-10-19 17:00:00|80.843945456961976|4|2301200046|61|35.216652492421872|0|59|1475|-80.826724|485|35.195689|SUSHI CLASSIC|0.0|6|CALIFORNIA ROLL (BROWN RICE)|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|35.232478750868765|00023012000462|SUSHI|DELI|-80.844274|80.844274157525618|412|1
35.204336|b21e7c4e6647374f41e24da165fbf418d168010e|4.99|2014-09-29 08:19:00|1.4094857484078087|4|7468210722|61|0.6144315741783704|0|26|139|-80.844274|20|35.204336|REMAINING SHELF STABLE JUICES|0.0|1|KNUDSEN JUICE MORNING BLEND|d1084d93d2f0e09baec1ee751c5c66b545b35033|0.8510398831336001|0.61471665291522548|00074682107227|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.844274|1.4109987626844462|61|1
35.585842|3c4145e20844bf69f9330b9ac64c5626b343942a|9.99|2014-10-18 16:39:00|1.4102725052409182|1|7962100001|99|0.6210901099944839|0|1|1489|-80.875654|100|35.585842|STACK PACK BACON|0.0|19|WRIGHTS HICKORY SMOKED BACON|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00079621461002|BACON|CASE READY MEATS|-80.875654|1.411546447003722|99|1
35.585842|e42025c21aef11d426d52c3f1d6de6e40df6b676|4.95|2015-01-19 12:09:00|1.4102725052409182|1|7447024102|99|0.6210901099944839|0|1|6789|-80.875654|1568|35.585842|MAGAZINES QUARTERLY|0.0|18|CHARLESTON DESIGN|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00074470241027|MAGAZINES|GM|-80.875654|1.411546447003722|99|1
35.585842|288fbe7897fc0fa08105f978328c46cc32fc834f|3.99|2014-11-14 09:45:00|1.4102725052409182|1|3000005620|99|0.6210901099944839|0|1|228|-80.875654|36|35.585842|TABLE SYRUP|1.0|1|AUNT JEMIMA ORIGINAL SYRUP|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00030000059708|TABLE SYRUPS|G1 GROCERY|-80.875654|1.411546447003722|99|1
35.585842|9e8c102088b562bef4c288a6ffc099dd0add5bd2|2.49|2015-02-14 13:06:00|1.4102725052409182|1|2529300224|99|0.6210901099944839|0|1|341|-80.875654|57|35.585842|CREAMERS|0.0|3|SILK ALMOND VANILLA CREAMER|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00025293002241|MILK|DAIRY|-80.875654|1.411546447003722|99|1
35.585842|2403301007a38ac54fd65009e41e5a580f4f931a|16.99|2014-09-19 16:50:00|1.4102725052409182|1|1820096721|99|0.6210901099944839|0|1|455|-80.875654|82|35.585842|DOMESTIC PREMIUM 12PK&>|0.0|16|MICHELOB ULTRA 18PK 12OZ CANS|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00018200967214|DOMESTIC BEER|BEER|-80.875654|1.411546447003722|99|1
35.585842|526a3115026bb9960b6e5e7049abdfeb01828b52|16.99|2015-02-28 15:17:00|1.4102725052409182|1|1820096721|99|0.6210901099944839|0|1|455|-80.875654|82|35.585842|DOMESTIC PREMIUM 12PK&>|0.0|16|MICHELOB ULTRA 18PK 12OZ CANS|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00018200967214|DOMESTIC BEER|BEER|-80.875654|1.411546447003722|99|1
35.585842|b4dc6bd6f1d86d80aed0bdc5ad35fabd8e82ac95|21.4|2015-02-08 13:11:00|1.4102725052409182|1|20898900000|99|0.6210901099944839|0|1|1421|-80.875654|201|35.585842|SMART CHICKEN VEGETABLE FED|0.0|2|SMART CHICKEN BONELESS BREAST|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00208989000008|POULTRY|MEAT|-80.875654|1.411546447003722|99|2
35.585842|5eeecea4b246bd618491ff5a868ed9089bdc1378|26.700000000000003|2015-01-24 16:26:00|1.4102725052409182|1|20898900000|99|0.6210901099944839|0|1|1421|-80.875654|201|35.585842|SMART CHICKEN VEGETABLE FED|2.9699999999999998|2|SMART CHICKEN BONELESS BREAST|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00208989000008|POULTRY|MEAT|-80.875654|1.411546447003722|99|3
35.585842|5a12368425f2a662a2937dfdd1d18a3042813aae|2.29|2014-09-24 11:42:00|1.4102725052409182|1|7225100105|99|0.6210901099944839|0|1|238|-80.875654|38|35.585842|RICE FLAVORED|0.29|1|NEAR EAST RICE SPANISH|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00072251000306|RICE GRAINS AND BEANS|G1 GROCERY|-80.875654|1.411546447003722|99|1
35.585842|c15b5cd0d670fe73c9511d5fd4254e46f9e991f3|3.39|2014-12-27 11:50:00|1.4102725052409182|1|1312000286|99|0.6210901099944839|0|1|1469|-80.875654|278|35.585842|REGULAR CUT FRIES|0.0|5|ORE-IDA ZESTIES|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00013120004841|FROZEN POTATO|FROZEN|-80.875654|1.411546447003722|99|1
35.585842|537e5ead9a18daf9b88e566135fc5bffc03af45b|2.35|2015-02-19 13:05:00|1.4102725052409182|1|1480000010|99|0.6210901099944839|0|1|104|-80.875654|16|35.585842|APPLESAUCE-CUPS|0.0|1|MOTTS 6PK APLSC SWEETENED|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00014800000108|FRUIT-CAN/JAR|G1 GROCERY|-80.875654|1.411546447003722|99|1
35.585842|4aa195524b604df41f7a6fd6105e41c5589a55bb|3.19|2014-09-13 15:37:00|1.4102725052409182|1|1800081778|99|0.6210901099944839|0|1|326|-80.875654|54|35.585842|COOKIES/BROWNIES-REFRIGERATED|0.69|3|PILLSURY RTB SUGAR|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00018000817726|DOUGH PRODUCTS|DAIRY|-80.875654|1.411546447003722|99|1
35.585842|f440d1651234877a00088b02c9a3fe4339a481e8|8.49|2014-09-15 16:38:00|1.4102725052409182|1|4173601014|99|0.6210901099944839|0|1|194|-80.875654|30|35.585842|OLIVE OIL|2.0|1|FILIPPO BERIO EX VIRGIN OLIVE|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00041736010147|SHORTENING/OIL|G1 GROCERY|-80.875654|1.411546447003722|99|1
35.585842|5034325b6f1260b12576a61d3a36444fd744254c|3.93|2014-11-26 16:31:00|1.4102725052409182|1|20394300000|99|0.6210901099944839|0|1|643|-80.875654|137|35.585842|PORK OFFALS-FROZEN|0.0|2|MORTY PRIDE SMOKED HOCKS|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00203943000001|PORK|MEAT|-80.875654|1.411546447003722|99|1
35.585842|c7222fcb539faf65c1ac792aa29810e334844947|4.58|2015-02-15 15:55:00|1.4102725052409182|1|4112907700|99|0.6210901099944839|0|1|1219|-80.875654|275|35.585842|PASTA SC CORE|0.0|1|CLASSICO SC FIRE RSTD TOM GAR|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00041129077009|PASTA SAUCES|G1 GROCERY|-80.875654|1.411546447003722|99|2
35.585842|25a147539d9ad332636c50766e9279c1c78acd0a|2.99|2014-10-12 16:25:00|1.4102725052409182|1||99|0.6210901099944839|0|1|561|-80.875654|64|35.585842|FR PROD ORGANIC PRODUCE|1.0|4|ORG CELERY|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00294070000002|FRESH PRODUCE|PRODUCE|-80.875654|1.411546447003722|99|1
35.585842|8f574d2e6dbd3a69625e5eb9f939f950c0f3157a|1.39|2014-11-23 15:01:00|1.4102725052409182|1|4144310303|99|0.6210901099944839|0|1|242|-80.875654|39|35.585842|CANNED BEANS|0.0|1|M HOLMES SND PINTO BEANS|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00041443119539|VEGETABLES-CAN/JAR|G1 GROCERY|-80.875654|1.411546447003722|99|1
35.585842|7916103dd95923877b2eff05ab2b0dc65bef6dd6|2.59|2014-11-17 16:47:00|1.4102725052409182|1|7203663996|99|0.6210901099944839|0|1|342|-80.875654|57|35.585842|FRESH MILK|0.0|3|HARRIS TEETER 2%   MILK|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00072036639998|MILK|DAIRY|-80.875654|1.411546447003722|99|1
35.585842|6556caafff802004fb7ca56f6a7ef93544df4e42|2.99|2015-02-22 15:45:00|1.4102725052409182|1|38137004666|99|0.6210901099944839|0|1|4816|-80.875654|1235|35.585842|FIRST AID ADHESIVE BANDG|0.0|17|BAND AID CLEAR SPOTS|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00381370047087|FIRST AID|HBC|-80.875654|1.411546447003722|99|1
35.585842|ebbec5234d1f5b5d04e0cc70680756523bf2e3f6|4.99|2014-10-26 11:48:00|1.4102725052409182|1|71575620002|99|0.6210901099944839|0|1|504|-80.875654|64|35.585842|FRESH BERRIES|2.5|4|STRAWBERRIES 1LB CLAM|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00715756200023|FRESH PRODUCE|PRODUCE|-80.875654|1.411546447003722|99|1
35.585842|b317e8f1342398ae36663651d9ec9ade1dec7000|7.34|2015-01-11 13:00:00|1.4102725052409182|1||99|0.6210901099944839|0|1|503|-80.875654|64|35.585842|FRESH GRAPES|0.0|4|GREEN GRAPES, SEEDLESS 12/16|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00204022000004|FRESH PRODUCE|PRODUCE|-80.875654|1.411546447003722|99|1
35.585842|93928049f0e60865470df9e8dfb1dedac74734f7|2.89|2014-10-21 12:42:00|1.4102725052409182|1|3800040260|99|0.6210901099944839|0|1|1269|-80.875654|41|35.585842|BREAKFAST SYRUP CARRIER|0.0|5|EGGO BUTTERMILK WAFFLES|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00038000402906|BREAKFAST FOODS FROZEN|FROZEN|-80.875654|1.411546447003722|99|1
35.585842|05043b3b2fe948aad899d5f9581ae35834b624e2|2.89|2014-11-09 16:52:00|1.4102725052409182|1|7203663125|99|0.6210901099944839|0|1|1262|-80.875654|57|35.585842|HALF N HALF WHIPPING CREAM|0.0|3|HT HEAVY WHIPPING CREAM|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00072036630988|MILK|DAIRY|-80.875654|1.411546447003722|99|1
35.585842|8f6fb1a7dbe29058e4555a8c42258f5eb4107f58|3.29|2014-10-28 17:12:00|1.4102725052409182|1|7203695076|99|0.6210901099944839|0|1|1609|-80.875654|371|35.585842|TAKE & BAKE BREAD|0.0|14|TAKE & BAKE SMALL WHEAT FRENCH|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00072036950765|BREAD|BAKERY|-80.875654|1.411546447003722|99|1
35.585842|b98ac4151b958765cc6589d6de8c5c4e025de734|4.99|2014-11-26 12:07:00|1.4102725052409182|1|7002500010|99|0.6210901099944839|0|1|361|-80.875654|105|35.585842|BREAKFAST SAUSAGE|0.0|19|NEESE COUNTRY SAUSAGE HOT|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00070025000118|BREAKFAST SAUSAGE|CASE READY MEATS|-80.875654|1.411546447003722|99|1
35.585842|f95864264d37106a513876a229304ac2bf27e878|4.39|2014-11-02 14:08:00|1.4102725052409182|1|5480001008|99|0.6210901099944839|0|1|239|-80.875654|38|35.585842|RICE-PACKAGED & BULK|0.0|1|UNCLE BENS RICE CONVERTED 32|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00054800010080|RICE GRAINS AND BEANS|G1 GROCERY|-80.875654|1.411546447003722|99|1
35.585842|463f4b8738cd639cb52eb20771f90598d031fc71|2.39|2015-02-23 18:43:00|1.4102725052409182|1|2529360040|99|0.6210901099944839|0|1|341|-80.875654|57|35.585842|CREAMERS|0.72|3|SILK FRENCH VANILLA CREAMER|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00025293600430|MILK|DAIRY|-80.875654|1.411546447003722|99|1
35.585842|c23a7ef7162ca16a32645cb458b31662f61442f8|9.58|2014-10-09 10:58:00|1.4102725052409182|1|20165500000|99|0.6210901099944839|0|1|297|-80.875654|49|35.585842|GROUND BEEF|0.0|2|HT PREMIUM GRND BEEF 80% LEAN|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00201655000005|BEEF|MEAT|-80.875654|1.411546447003722|99|2
35.585842|fef190da84d976a38984f37e27ed61ae82e04577|7.69|2014-12-03 16:04:00|1.4102725052409182|1|30045025708|99|0.6210901099944839|0|1|4236|-80.875654|1200|35.585842|DEX ADULT/CHILDREN|2.7|17|TYL COLD M/S NIGHTTIME LIQUID|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00300450269089|COUGH/COLD/SINUS|HBC|-80.875654|1.411546447003722|99|1
35.585842|07d896bf6acf43c2f42240260d602cd75cd7fc1e|3.15|2014-11-03 20:26:00|1.4102725052409182|1|7225003706|99|0.6210901099944839|0|1|1026|-80.875654|162|35.585842|WHEAT|0.86|7|NATOWN HONEYWHEAT BRD|d543107d523bc1e850f259734a1320fbf9bb84f1|3.4838838961298753|0.61833652052202714|00072250037068|SLICED BREAD|COMMERCIAL BAKERY|-80.875654|1.411546447003722|99|1
35.444615|77db651442ec47560c3a2a41e291b3031861e3a5|3.89|2014-09-28 17:53:00|1.4102725052409182|4|7184005080|340|0.6186252338517699|0|1|580|-80.861571|136|35.444615|OTHER MERCH DRESSINGS|0.0|4|MARIES COLE SLAW DRESSING|d6a98e608896c62f0f3e530d95d1b73d167efcc0|1.8509290874421198|0.61833652052202714|00071840043304|OTHER MERCHANDISE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|f6acf7bcf394b7082b645f0bc6ec6191d39aaec3|5.49|2014-12-21 16:11:00|1.4102725052409182|4|2900001628|340|0.6186252338517699|0|1|1244|-80.861571|21|35.444615|OTHER NUTS|1.0|1|PLANTERS BRITTLE NUT MEDLEY|d6a98e608896c62f0f3e530d95d1b73d167efcc0|1.8509290874421198|0.61833652052202714|00029000016286|NUTS|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.444615|97f0c6590acb5418bd3c4f25f305c1bcd0a1ab40|25.96|2014-12-05 17:21:00|80.86161257435397|4|1200080994|340|35.471402174227137|0|36|55|-80.893784|8|35.478031|REGULAR|0.0|23|PEPSI FRIDGEMATE|d6a98e608896c62f0f3e530d95d1b73d167efcc0|1.8509290874421198|35.472272108304431|00012000809941|CARBONATED BEVERAGES|BEVERAGE|-80.861571|80.861577580668666|179|4
35.444615|891380d6e37be5ed629ba0c3e6d787f2f29c07e1|2.65|2014-10-12 15:44:00|1.4102725052409182|4|1600026460|340|0.6186252338517699|0|1|42|-80.861571|6|35.444615|GRANOLA/YOGURT BARS|0.0|1|NV BAR SWT SLTY ALMND.|d6a98e608896c62f0f3e530d95d1b73d167efcc0|1.8509290874421198|0.61833652052202714|00016000277069|BREAKFAST FOODS|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.444615|0b2205cf1c7dc0cc3e99f5d673f27b2915c711a9|1.79|2015-01-27 18:35:00|1.4102725052409182|4|1800000261|340|0.6186252338517699|0|1|325|-80.861571|54|35.444615|BISCUITS-REFRIGERATED|0.0|3|GRANDS FLAKY BISCUITS|d6a98e608896c62f0f3e530d95d1b73d167efcc0|1.8509290874421198|0.61833652052202714|00018000002610|DOUGH PRODUCTS|DAIRY|-80.861571|1.4113006522851637|340|1
35.444615|92e5483c3e7bcbbba522144bfc27fe93f8625f33|13.98|2014-12-13 17:06:00|1.4102725052409182|4|1820005989|340|0.6186252338517699|0|1|455|-80.861571|82|35.444615|DOMESTIC PREMIUM 12PK&>|0.0|16|MICHELOB ULTRA 6PK 12OZ  BTL|d6a98e608896c62f0f3e530d95d1b73d167efcc0|1.8509290874421198|0.61833652052202714|00018200059896|DOMESTIC BEER|BEER|-80.861571|1.4113006522851637|340|2
35.444615|71cf9802a440ed0b4173c1e720a2eb7bb101ac6b|1.29|2014-12-01 13:19:00|80.86161257435397|4|8379152001|340|35.471402174227137|0|36|1981|-80.893784|480|35.478031|CHIPS|0.0|6|DIRTY POTATO CHIP SOUR CRM|d6a98e608896c62f0f3e530d95d1b73d167efcc0|1.8509290874421198|35.472272108304431|00083791520094|DRY GOODS|DELI|-80.861571|80.861577580668666|179|1
35.444615|f2577b7dd2b21656193c55262a5679952a20769d|1.29|2014-10-23 13:12:00|80.86161257435397|4|8379152001|340|35.471402174227137|0|36|1981|-80.893784|480|35.478031|CHIPS|0.0|6|DIRTY POTATO CHIP SOUR CRM|d6a98e608896c62f0f3e530d95d1b73d167efcc0|1.8509290874421198|35.472272108304431|00083791520094|DRY GOODS|DELI|-80.861571|80.861577580668666|179|1
35.444615|1df54290fac742c65c94a0a74bff68805fc05bb1|2.69|2015-02-01 14:21:00|1.4102725052409182|4|70935100013|340|0.6186252338517699|0|1|556|-80.861571|64|35.444615|PACKAGED VEGETABLES|0.0|4|APIO BROCCOLI & CAULIFLOWER|d6a98e608896c62f0f3e530d95d1b73d167efcc0|1.8509290874421198|0.61833652052202714|00709351000263|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|5c4822043aaa645cc51219497178678b7ad22260|0.75|2015-01-05 18:32:00|1.4102725052409182|4||340|0.6186252338517699|0|1|500|-80.861571|64|35.444615|FRESH APPLES|0.0|4|ROME APPLE EASTERN|d6a98e608896c62f0f3e530d95d1b73d167efcc0|1.8509290874421198|0.61833652052202714|00204171000009|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|a077a975cf5fba8019e5920a0a87d8bfdf8c55c4|6.58|2014-09-21 19:59:00|80.86161257435397|4|3746608323|340|35.471402174227137|0|36|62|-80.893784|7|35.478031|SPECIALTY BAR/BOX CHOCOLATE|3.3|1|LINDT BAR EXCEL CHOC COCONUT|d6a98e608896c62f0f3e530d95d1b73d167efcc0|1.8509290874421198|35.472272108304431|00037466062266|CANDY|G1 GROCERY|-80.861571|80.861577580668666|179|2
35.444615|8f507cdb6969d2ba967ed422c25fe607bff12328|3.59|2015-03-07 15:16:00|1.4102725052409182|4|1660000071|340|0.6186252338517699|0|1|207|-80.861571|32|35.444615|COCKTAIL MIXES|0.0|1|ROSES LIME JUICE-12 OZ PLASTIC|d6a98e608896c62f0f3e530d95d1b73d167efcc0|1.8509290874421198|0.61833652052202714|00016600000043|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.861571|1.4113006522851637|340|1
35.444615|d156415e51f886d6a36abb369a8ae92cd9f06833|5.0|2014-11-24 15:32:00|1.4102725052409182|4|8500001581|340|0.6186252338517699|0|1|9943|-80.861571|885|35.444615|NFS POP RIESLING|0.0|13|BAREFOOT RIESLING|d6a98e608896c62f0f3e530d95d1b73d167efcc0|1.8509290874421198|0.61833652052202714|00085000015810|POPULAR (4-$7.99)|WINE|-80.861571|1.4113006522851637|340|1
35.444615|465c30feecf636377a7b0154ec2e6844bbea9a5e|2.99|2015-01-18 15:02:00|1.4102725052409182|4|20443000000|340|0.6186252338517699|0|1|510|-80.861571|64|35.444615|FRESH PINEAPPLE|0.0|4|GOLD PINEAPPLES|d6a98e608896c62f0f3e530d95d1b73d167efcc0|1.8509290874421198|0.61833652052202714|00643126072003|FRESH PRODUCE|PRODUCE|-80.861571|1.4113006522851637|340|1
35.444615|e7a9d936335cd19da13c8540118f8aeb346304b5|5.79|2014-10-17 17:28:00|80.86161257435397|4|78978501962|340|35.471402174227137|0|36|273|-80.893784|43|35.478031|PREMIUM NOVELTIES|0.0|5|SKINNYCOW BEST OF BOTH SWIRLED|d6a98e608896c62f0f3e530d95d1b73d167efcc0|1.8509290874421198|35.472272108304431|00789785020013|FROZEN NOVELTIES|FROZEN|-80.861571|80.861577580668666|179|1
35.41832|c551ded77a7974c9d3e5a7c0c138dc81a9c17835|4.59|2015-02-17 16:39:00|1.4102725052409182|3|3377601795|190|0.6181662995249579|0|1|313|-80.746334|51|35.41832|MARGARINE|2.3|3|SMART BAL SPRDABL BUTTER 15 OZ|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00033776017958|BUTTER & MARGARINE|DAIRY|-80.746334|1.409289387215043|190|1
35.41832|50160eea14a2a124b83f9d1a5198b7dccb6d3b93|4.58|2014-10-10 18:30:00|1.4102725052409182|3|7203653023|190|0.6181662995249579|0|1|1273|-80.746334|50|35.41832|BAG VEG NON STEAM|0.58|5|HT CUT GREEN BEANS|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036530356|VEGETABLES-FROZEN|FROZEN|-80.746334|1.409289387215043|190|2
35.41832|28264d59de340c1db2db293ebb2181652093a4c0|2.99|2015-02-01 08:53:00|1.4102725052409182|3|7203653055|190|0.6181662995249579|0|1|1273|-80.746334|50|35.41832|BAG VEG NON STEAM|0.0|5|HT BABY LIMA BEANS|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036530554|VEGETABLES-FROZEN|FROZEN|-80.746334|1.409289387215043|190|1
35.41832|2f454a0a674223ebb180aec1fa0dd0d21ec8d930|15.98|2014-11-16 16:59:00|1.4102725052409182|3|7005700210|190|0.6181662995249579|0|1|670|-80.746334|146|35.41832|CRAB PACKAGED|0.0|12|PHILLIPS CLAW CRABMEAT PAST|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00070057002104|CRAB|SEAFOOD|-80.746334|1.409289387215043|190|2
35.41832|1998286175fd97c2f60b53bfdfb4f5c70cf2980b|3.55|2014-12-02 12:23:00|1.4102725052409182|3|7332100027|190|0.6181662995249579|0|1|251|-80.746334|43|35.41832|NON-DAIRY NOVELTIES|1.78|5|LUIGI'S ITALIAN ICE LEMON|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00073321000271|FROZEN NOVELTIES|FROZEN|-80.746334|1.409289387215043|190|1
35.41832|35a87da3429a793b8eec47e7819c80dc474a334a|2.49|2014-11-23 15:34:00|1.4102725052409182|3|7203688048|190|0.6181662995249579|0|1|526|-80.746334|64|35.41832|FRESH MUSHROOMS|0.0|4|HT SLICED BABY BELLAS|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036880482|FRESH PRODUCE|PRODUCE|-80.746334|1.409289387215043|190|1
35.41832|6cb6ffca5756642fdb1c3b1bd5c3bc775b27f9aa|5.78|2014-11-07 14:30:00|1.4102725052409182|3|7203697887|190|0.6181662995249579|0|1|61|-80.746334|9|35.41832|RTE CEREAL ADULT|0.92|1|HT CER CRUNCH GRAN RAISIN BRAN|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036978899|CEREAL|G1 GROCERY|-80.746334|1.409289387215043|190|2
35.41832|e5b5f908178440f7b7af9d732a0fbf5e7330299e|8.67|2014-10-19 12:46:00|1.4102725052409182|3|7203697887|190|0.6181662995249579|0|1|61|-80.746334|9|35.41832|RTE CEREAL ADULT|0.92|1|HT CER CRUNCH GRAN RAISIN BRAN|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036978899|CEREAL|G1 GROCERY|-80.746334|1.409289387215043|190|3
35.41832|161faa9eb9215a219de659f4f1d7c0c174da8ca8|2.89|2014-10-28 21:27:00|1.4102725052409182|3|7203697887|190|0.6181662995249579|0|1|61|-80.746334|9|35.41832|RTE CEREAL ADULT|0.92|1|HT CER CRUNCH GRAN RAISIN BRAN|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036978899|CEREAL|G1 GROCERY|-80.746334|1.409289387215043|190|1
35.41832|c5d866eb433f92bdbd7ffad68a1067bc6b4f8051|5.78|2014-09-27 11:33:00|1.4102725052409182|3|7203697887|190|0.6181662995249579|0|1|61|-80.746334|9|35.41832|RTE CEREAL ADULT|1.39|1|HT CER CRUNCH GRAN RAISIN BRAN|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036978899|CEREAL|G1 GROCERY|-80.746334|1.409289387215043|190|2
35.41832|00da597ea4121d6abd193cbd24872c01317e7120|2.5|2014-10-05 10:28:00|1.4102725052409182|3|7203671406|190|0.6181662995249579|0|1|61|-80.746334|9|35.41832|RTE CEREAL ADULT|0.23|1|HT CER RAISIN BRAN|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036520364|CEREAL|G1 GROCERY|-80.746334|1.409289387215043|190|1
35.41832|f51d120e46b23e40875ae1a8f1c79b965e351014|3.59|2014-11-16 17:06:00|1.4102725052409182|3|7225006580|190|0.6181662995249579|0|1|1033|-80.746334|163|35.41832|HAMBURGER|0.6|7|CBC SESAME TWIST HAMBURGER BUN|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072250065801|BUNS/ROLLS|COMMERCIAL BAKERY|-80.746334|1.409289387215043|190|1
35.41832|95dca4804ec56e10f519b6a545a55e8e993525e3|6.78|2014-09-21 15:37:00|1.4102725052409182|3|20668800000|190|0.6181662995249579|0|1|1830|-80.746334|415|35.41832|FFM SLICING CHEESE|0.0|6|HT YELLOW AMERICAN|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00206687000009|SLICING CHEESE|DELI|-80.746334|1.409289387215043|190|1
35.41832|0b62f833259dab3f9280c1e7cbaa47476a6d4f5a|8.39|2015-01-13 07:25:00|1.4102725052409182|3|20668800000|190|0.6181662995249579|0|1|1830|-80.746334|415|35.41832|FFM SLICING CHEESE|0.0|6|HT YELLOW AMERICAN|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00206687000009|SLICING CHEESE|DELI|-80.746334|1.409289387215043|190|1
35.41832|088af66eba7b93988ed5ca9a5eb0b57429f7b515|6.92|2014-11-13 18:15:00|1.4102725052409182|3|20668800000|190|0.6181662995249579|0|1|1830|-80.746334|415|35.41832|FFM SLICING CHEESE|0.99|6|HT YELLOW AMERICAN|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00206687000009|SLICING CHEESE|DELI|-80.746334|1.409289387215043|190|1
35.41832|dcabdaee4531a66f8cda237aa85fc652022e2840|6.98|2015-02-20 16:15:00|1.4102725052409182|3|20967400000|190|0.6181662995249579|0|1|669|-80.746334|146|35.41832|CRAB VALUE ADDED|0.0|12|MARYLAND STYLE CRAB CAKES 4 OZ|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00209674000006|CRAB|SEAFOOD|-80.746334|1.409289387215043|190|1
35.41832|2fef6286df504403c0f269a04239e5ca0de27ed6|9.17|2014-12-15 17:19:00|1.4102725052409182|3|20541200000|190|0.6181662995249579|0|1|1832|-80.746334|415|35.41832|BH SLICING CHEESE|0.0|6|BOARS HEAD YELLOW AMER CHEESE|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00205412000000|SLICING CHEESE|DELI|-80.746334|1.409289387215043|190|1
35.41832|8fb4bb6c009d8a6ff47737dc2387dc6a3e9aedfe|1.97|2015-02-15 09:20:00|80.749667378538092|3|7203629075|190|35.437367625817508|0|3|1211|-80.762919|272|35.442529|HISP SALSA/DIPS|0.0|1|HT PICANTE MEDIUM|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|35.465179900649026|00072036290724|HISPANIC PREP. FOODS|G1 GROCERY|-80.746334|80.74633811067487|471|1
35.41832|15d429c4b69fc5c7fd1822e7f198eacd9eafda82|2.89|2014-11-21 07:53:00|1.4102725052409182|3|7203663102|190|0.6181662995249579|0|1|339|-80.746334|57|35.41832|EGGNOGS/DRINKS|0.39|3|I/O HARRIS TEETER EGG NOG|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036631022|MILK|DAIRY|-80.746334|1.409289387215043|190|1
35.41832|8ad6b3614ea15deba289eb5fe9a53236063b4891|3.67|2015-01-14 17:17:00|1.4102725052409182|3|7203655019|190|0.6181662995249579|0|1|332|-80.746334|52|35.41832|STRING/SNACK|0.0|3|HT STRING CHEESE|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036550194|CHEESE|DAIRY|-80.746334|1.409289387215043|190|1
35.41832|4244f536e31c18eb6d8ec6a6a76913e85649f374|2.58|2015-01-06 18:15:00|1.4102725052409182|3|7203678692|190|0.6181662995249579|0|1|1208|-80.746334|23|35.41832|WHSE PASTA VALUE ADD|0.0|1|HTO WW SPAGHETTI|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036786920|PASTA|G1 GROCERY|-80.746334|1.409289387215043|190|2
35.41832|74e1136440063c765b43eec5c5b0894d58a17ffb|2.38|2015-02-24 18:58:00|1.4102725052409182|3|7488007017|190|0.6181662995249579|0|1|80|-80.746334|34|35.41832|SEASONING PACKETS|0.38|1|SUNBIRD STIR FRY MIX|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00074880070040|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.746334|1.409289387215043|190|2
35.41832|a5f10d8616583f80d940b30694f4d0b343936ac7|0.8|2014-10-18 08:49:00|1.4102725052409182|3||190|0.6181662995249579|0|1|502|-80.746334|64|35.41832|FRESH BANANAS|0.0|4|BANANAS, YELLOW|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.746334|1.409289387215043|190|1
35.41832|2be6129738f4454f07260efd9746abde50137567|1.19|2015-02-18 18:44:00|1.4102725052409182|3|73801577713|190|0.6181662995249579|0|1|545|-80.746334|64|35.41832|FRESH SPROUTS|0.0|4|BEAN SPROUTS,  PKG|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00738015777135|FRESH PRODUCE|PRODUCE|-80.746334|1.409289387215043|190|1
35.41832|80490f5991e459c0b2c2b9efc6d6c557c125bf7c|1.19|2015-01-21 16:49:00|1.4102725052409182|3|73801577713|190|0.6181662995249579|0|1|545|-80.746334|64|35.41832|FRESH SPROUTS|0.0|4|BEAN SPROUTS,  PKG|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00738015777135|FRESH PRODUCE|PRODUCE|-80.746334|1.409289387215043|190|1
35.41832|4b808099d682bb3087177a88b6e4b4360e192058|9.06|2015-01-05 07:44:00|1.4102725052409182|3||190|0.6181662995249579|0|1|561|-80.746334|64|35.41832|FR PROD ORGANIC PRODUCE|0.0|4|ORG HH BUNCH TOMATOES|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00294664000005|FRESH PRODUCE|PRODUCE|-80.746334|1.409289387215043|190|1
35.41832|021df77b39cbe33e7631ec92abc2772c76f2610d|0.55|2014-10-20 19:52:00|1.4102725052409182|3||190|0.6181662995249579|0|1|545|-80.746334|64|35.41832|FRESH SPROUTS|0.0|4|COO BEAN SPROUTS, BULK|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00204536000002|FRESH PRODUCE|PRODUCE|-80.746334|1.409289387215043|190|1
35.41832|0c1dc2ebbc259782d2a5f832fc27520733e812b7|2.54|2015-01-13 21:06:00|1.4102725052409182|3||190|0.6181662995249579|0|1|535|-80.746334|64|35.41832|FRESH GREENS|0.0|4|COO TURNIP GREENS, BULK|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00204619000004|FRESH PRODUCE|PRODUCE|-80.746334|1.409289387215043|190|1
35.41832|c930b2895a3a1c6bee4c348cb4507cbac3a52338|1.25|2014-09-11 20:11:00|80.749667378538092|3||190|35.437367625817508|0|3|502|-80.762919|64|35.442529|FRESH BANANAS|0.0|4|BANANAS, YELLOW|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|35.465179900649026|00204011000008|FRESH PRODUCE|PRODUCE|-80.746334|80.74633811067487|471|1
35.41832|5fc9e4f43f1214e15d288277d4e551eab33e8203|4.49|2014-11-10 07:39:00|1.4102725052409182|3|2570071147|190|0.6181662995249579|0|1|442|-80.746334|76|35.41832|NFS-COOKING-STORAGE BAGS|1.49|1|ZIPLOC SANDWICH BAGS|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00025700003915|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.746334|1.409289387215043|190|1
35.41832|c0aaec03a6b8dd6e546409a84bdc3c45964cb62e|0.8|2014-10-12 22:54:00|1.4102725052409182|3|7047000100|190|0.6181662995249579|0|1|687|-80.746334|61|35.41832|BLENDED|0.3|3|YOPLAIT VANILLA CUSTARD|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00070470001128|YOGURT|DAIRY|-80.746334|1.409289387215043|190|1
35.41832|fc73aafc06a0d41d93841dec524fc090c7b2d076|3.29|2014-11-30 19:25:00|1.4102725052409182|3|2840004768|190|0.6181662995249579|0|1|202|-80.746334|31|35.41832|PRETZELS|0.29|1|ROLD GOLD PRETZEL CLASSIC THIN|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00028400047678|SNACKS|G1 GROCERY|-80.746334|1.409289387215043|190|1
35.41832|1f07066db6893687965aeb58bf847ef3777359c7|3.29|2014-10-19 19:20:00|1.4102725052409182|3|2840004768|190|0.6181662995249579|0|1|202|-80.746334|31|35.41832|PRETZELS|0.79|1|ROLD GOLD PRETZEL CLASSIC THIN|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00028400047678|SNACKS|G1 GROCERY|-80.746334|1.409289387215043|190|1
35.41832|11d013b05fa716cabee6655de545a086f3156b1f|2.99|2014-09-20 12:42:00|80.749667378538092|3||190|35.437367625817508|0|3|542|-80.762919|64|35.442529|FRESH VEGETABLES REMAIN|0.0|4|RED BUN BEETS (RPC)|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|35.465179900649026|00204539000009|FRESH PRODUCE|PRODUCE|-80.746334|80.74633811067487|471|1
35.41832|6dfe485845beed60dccd7bc95875a936de088426|5.97|2014-12-17 06:10:00|1.4102725052409182|3|7203676359|190|0.6181662995249579|0|1|345|-80.746334|57|35.41832|ORGANIC MILK|0.0|3|HTO ORGANIC 1% MILK GAL|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036763617|MILK|DAIRY|-80.746334|1.409289387215043|190|1
35.41832|26f074c03039fcc4f7222486046a9ceb2738e064|20.55|2015-02-17 18:05:00|1.4102725052409182|3|20897500000|190|0.6181662995249579|0|1|977|-80.746334|201|35.41832|FRESH HT CHICKEN|10.3|2|FRESH BONELESS CHICKEN BREAST|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00208975000005|POULTRY|MEAT|-80.746334|1.409289387215043|190|1
35.41832|7285dab6ce55aa3748c92889068428456cde2594|0.56|2014-10-12 16:10:00|1.4102725052409182|3||190|0.6181662995249579|0|1|534|-80.746334|64|35.41832|FRESH CHILI PEPPERS|0.0|4|COO ORANGE HABANERO CHILI|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00204711000001|FRESH PRODUCE|PRODUCE|-80.746334|1.409289387215043|190|1
35.41832|1f629ee28941922db0a2893b6b6fe995c7afb0f7|6.0|2015-01-12 08:40:00|80.749667378538092|3|20966900000|190|35.437367625817508|0|3|669|-80.762919|146|35.442529|CRAB VALUE ADDED|0.0|12|THE CHARLESTON CRABCAKE4 OZ EA|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|35.465179900649026|00209669000004|CRAB|SEAFOOD|-80.746334|80.74633811067487|471|1
35.41832|ef46a312602a9ebc13f2daa225cb3ea45e7930d8|3.99|2014-09-23 17:07:00|1.4102725052409182|3|3260190020|190|0.6181662995249579|0|1|561|-80.746334|64|35.41832|FR PROD ORGANIC PRODUCE|0.49|4|EBF ORG SPINACH CLAM 5 OZ|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00032601900205|FRESH PRODUCE|PRODUCE|-80.746334|1.409289387215043|190|1
35.41832|7b7f7229ed51ccf029b745895db1017c74365788|3.0|2015-02-20 16:41:00|80.749667378538092|3|7203688157|190|35.437367622138417|0|3|556|-80.782849|64|35.372142|PACKAGED VEGETABLES|0.0|4|HT RV BRUSSEL SPROUTS|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|35.465179900649026|00072036881656|FRESH PRODUCE|PRODUCE|-80.746334|80.746349099124998|122|1
35.41832|0ccbe94a2fc8df61393c88c20282b390b5e5fadf|3.49|2014-10-02 18:44:00|1.4102725052409182|3|7225003712|190|0.6181662995249579|0|1|1026|-80.746334|162|35.41832|WHEAT|1.2|7|NATOWN 100% WHEAT BRD|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072250037129|SLICED BREAD|COMMERCIAL BAKERY|-80.746334|1.409289387215043|190|1
35.41832|aa123680db360ed7c00a29a332e21bf43f734926|6.3|2014-11-15 18:58:00|1.4102725052409182|3|7225003712|190|0.6181662995249579|0|1|1026|-80.746334|162|35.41832|WHEAT|1.58|7|NATOWN 100% WHEAT BRD|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072250037129|SLICED BREAD|COMMERCIAL BAKERY|-80.746334|1.409289387215043|190|2
35.41832|4b88712549f990ca8137662d769c85389c22e11a|2.99|2015-02-28 21:14:00|1.4102725052409182|3|7203698526|190|0.6181662995249579|0|1|201|-80.746334|31|35.41832|POTATO CHIPS|0.8|1|HT TRADER KETTLE CHIP REG|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036985279|SNACKS|G1 GROCERY|-80.746334|1.409289387215043|190|1
35.41832|7c8b4189ecdc8c5ae63f0a2b336d7e701b6ca82c|2.29|2014-09-18 20:56:00|1.4102725052409182|3|7660655611|190|0.6181662995249579|0|1|76|-80.746334|11|35.41832|MEAT SAUCES|0.0|1|TROPICAL PEPPER SCOTCH BONNET|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00076606556111|CONDIMENTS|G1 GROCERY|-80.746334|1.409289387215043|190|1
35.41832|8dce4a5b74df5513af82bb43ccc26beba4f8aaad|4.99|2014-10-02 20:35:00|1.4102725052409182|3|7203697885|190|0.6181662995249579|0|1|200|-80.746334|31|35.41832|MICROWAVE POPCORN|0.0|1|HTN ORGANIC POPCORN YELLOW|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036978851|SNACKS|G1 GROCERY|-80.746334|1.409289387215043|190|1
35.41832|eb84ee82089746a3569709ff265a6d79149511fa|1.88|2015-03-05 20:00:00|80.749667378538092|3||190|35.437367625817508|0|3|561|-80.762919|64|35.442529|FR PROD ORGANIC PRODUCE|0.21|4|ORG BANANAS|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|35.465179900649026|00294011000009|FRESH PRODUCE|PRODUCE|-80.746334|80.74633811067487|471|1
35.41832|a03b8846135e94e704766b68e28954063f3d9773|2.99|2014-11-23 13:26:00|1.4102725052409182|3|5844977731|190|0.6181662995249579|0|1|61|-80.746334|9|35.41832|RTE CEREAL ADULT|0.0|1|NAT PATH ORG CER HERITAG FLAKE|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00058449770206|CEREAL|G1 GROCERY|-80.746334|1.409289387215043|190|1
35.41832|ab6258a8993ed4828e59cb91059d987cb34c1d45|2.99|2015-02-12 08:08:00|1.4102725052409182|3|5844977731|190|0.6181662995249579|0|1|61|-80.746334|9|35.41832|RTE CEREAL ADULT|0.0|1|NAT PATH ORG CER HERITAG FLAKE|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00058449770206|CEREAL|G1 GROCERY|-80.746334|1.409289387215043|190|1
35.41832|04ebde488806c26807fe3470553e5d878ae52e29|2.99|2014-11-27 11:45:00|1.4102725052409182|3|5844977731|190|0.6181662995249579|0|1|61|-80.746334|9|35.41832|RTE CEREAL ADULT|0.0|1|NAT PATH ORG GRAN FLX PUMPK|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00058449890072|CEREAL|G1 GROCERY|-80.746334|1.409289387215043|190|1
35.41832|6aa64a8d7d457a6f5859a659e0b660c49e3ec866|0.37|2014-10-27 18:08:00|1.4102725052409182|3|7203659035|190|0.6181662995249579|0|1|688|-80.746334|61|35.41832|LIGHT|0.0|3|HT NONFAT PLAIN YOGURT|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036040299|YOGURT|DAIRY|-80.746334|1.409289387215043|190|1
35.41832|ba3b33e32c3711b4264b7d292a0b69ad769d1df6|2.74|2015-01-19 15:26:00|80.749667378538092|3|7203690021|190|35.437367625817508|0|3|1033|-80.762919|163|35.442529|HAMBURGER|0.0|7|H T HAMBURGER BUNS|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|35.465179900649026|00072036900210|BUNS/ROLLS|COMMERCIAL BAKERY|-80.746334|80.74633811067487|471|2
35.41832|6086b6e8916f06564ff8d62dbdb6eaecea0683f1|2.79|2014-10-25 10:17:00|1.4102725052409182|3|7203688035|190|0.6181662995249579|0|1|522|-80.746334|64|35.41832|FRESH TOMATOES|0.0|4|HT SLICING TOMATO 4 PK|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036880352|FRESH PRODUCE|PRODUCE|-80.746334|1.409289387215043|190|1
35.41832|6b882e171ffa19a71f3bea27ecfc8c6acd8c7f59|3.29|2014-12-01 22:02:00|1.4102725052409182|3|7203688035|190|0.6181662995249579|0|1|522|-80.746334|64|35.41832|FRESH TOMATOES|0.0|4|HT SLICING TOMATO 4 PK|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036880352|FRESH PRODUCE|PRODUCE|-80.746334|1.409289387215043|190|1
35.41832|ba9ee21b223b56299e61e003fd6992c634f92c1f|1.97|2014-10-05 14:39:00|1.4102725052409182|3|7203629075|190|0.6181662995249579|0|1|1211|-80.746334|272|35.41832|HISP SALSA/DIPS|0.0|1|HT SALSA MILD|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036290748|HISPANIC PREP. FOODS|G1 GROCERY|-80.746334|1.409289387215043|190|1
35.41832|39d4272bd45079bf933dd360ab707edcabce3752|1.97|2014-10-04 17:07:00|1.4102725052409182|3|7203629075|190|0.6181662995249579|0|1|1211|-80.746334|272|35.41832|HISP SALSA/DIPS|0.0|1|HT SALSA MILD|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036290748|HISPANIC PREP. FOODS|G1 GROCERY|-80.746334|1.409289387215043|190|1
35.41832|4667e3865218d5256acf9aa48835c3d0adf9f248|3.39|2015-01-09 08:27:00|1.4102725052409182|3|2529300098|190|0.6181662995249579|0|1|1265|-80.746334|57|35.41832|ALMOND MILK|0.39|3|SILK PURE ALMOND ORIGINAL|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00025293000988|MILK|DAIRY|-80.746334|1.409289387215043|190|1
35.41832|c94333ac84b443210f8a4dd41dd7fe7dcbca31a6|2.99|2015-01-18 11:07:00|1.4102725052409182|3|5844977731|190|0.6181662995249579|0|1|61|-80.746334|9|35.41832|RTE CEREAL ADULT|0.49|1|NAT PATH ORG GRAN CHIA COCONT|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00058449890331|CEREAL|G1 GROCERY|-80.746334|1.409289387215043|190|1
35.41832|e1dbf93e2b4715e33753b1d7166ffcf44b3c4d9d|4.74|2014-09-10 12:53:00|1.4102725052409182|3|7203670412|190|0.6181662995249579|0|1|252|-80.746334|45|35.41832|PREMIUM ICE CREAM|0.0|5|HIGHLAND CREST STRAWBERRY IC|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036704153|ICE CREAM|FROZEN|-80.746334|1.409289387215043|190|2
35.41832|f6147f75c70c1828f33a9f2bb3a7e3feae67c472|2.32|2014-11-02 20:35:00|1.4102725052409182|3||190|0.6181662995249579|0|1|522|-80.746334|64|35.41832|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00204664000004|FRESH PRODUCE|PRODUCE|-80.746334|1.409289387215043|190|1
35.41832|e4a52b7afcefb5a682b1c111dce03afe13333833|2.38|2015-01-25 17:23:00|1.4102725052409182|3||190|0.6181662995249579|0|1|522|-80.746334|64|35.41832|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00204664000004|FRESH PRODUCE|PRODUCE|-80.746334|1.409289387215043|190|1
35.41832|aabbcd280418dbb66547e8cc3b703e319b6f234f|2.99|2015-02-12 17:26:00|1.4102725052409182|3|7203659032|190|0.6181662995249579|0|1|321|-80.746334|53|35.41832|RICOTTA/FARMERS CHEESE|0.0|3|HT FAT FREE RICOTTA CHEESE|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036590336|CULTURES|DAIRY|-80.746334|1.409289387215043|190|1
35.41832|419241159373b7615447fbd324c6f3fab6a36cc3|5.38|2015-02-18 19:15:00|1.4102725052409182|3|2548400005|190|0.6181662995249579|0|1|579|-80.746334|136|35.41832|SOY/MEATLESS PRODUCTS|0.0|4|NASOYA EGG ROLL WRAPPER|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00025484000056|OTHER MERCHANDISE|PRODUCE|-80.746334|1.409289387215043|190|2
35.41832|26ff8e8c4fbcac38f732f973380c767a00242f23|2.99|2015-02-06 22:13:00|1.4102725052409182|3|5844977731|190|0.6181662995249579|0|1|61|-80.746334|9|35.41832|RTE CEREAL ADULT|0.0|1|NAT PATH ORG CER OPTIMUM BLBRY|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00058449777007|CEREAL|G1 GROCERY|-80.746334|1.409289387215043|190|1
35.41832|cddb0390065a75043f064e1871936a902a503b47|2.0|2014-09-14 19:28:00|1.4102725052409182|3|2840000210|190|0.6181662995249579|0|1|204|-80.746334|31|35.41832|TORTILLA CHIPS|0.0|1|SANTITAS WHITE CORN|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00028400002103|SNACKS|G1 GROCERY|-80.746334|1.409289387215043|190|1
35.41832|69c2f89c82d6d58616a50402cd4d4b8344b6f21b|2.0|2014-11-09 18:16:00|1.4102725052409182|3|2840000210|190|0.6181662995249579|0|1|204|-80.746334|31|35.41832|TORTILLA CHIPS|0.0|1|SANTITAS WHITE CORN|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00028400002103|SNACKS|G1 GROCERY|-80.746334|1.409289387215043|190|1
35.41832|629ad08075f812255074241711ff0722c343f0cd|0.89|2015-01-21 17:10:00|1.4102725052409182|3|20406800000|190|0.6181662995249579|0|1|524|-80.746334|64|35.41832|FRESH PROD FRESH ONIONS|0.0|4|GREEN ONIONS|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00033383605005|FRESH PRODUCE|PRODUCE|-80.746334|1.409289387215043|190|1
35.41832|1b3b9a3974198117b7efdab8fd2abd57c4cada88|5.97|2014-10-28 08:38:00|1.4102725052409182|3|7203676359|190|0.6181662995249579|0|1|345|-80.746334|57|35.41832|ORGANIC MILK|0.0|3|HTO ORGANIC FF SKIM GAL|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036763624|MILK|DAIRY|-80.746334|1.409289387215043|190|1
35.41832|e80358fa2f25d65102741f153c756c7bc9497d59|5.97|2014-10-10 08:54:00|1.4102725052409182|3|7203676359|190|0.6181662995249579|0|1|345|-80.746334|57|35.41832|ORGANIC MILK|0.0|3|HTO ORGANIC FF SKIM GAL|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036763624|MILK|DAIRY|-80.746334|1.409289387215043|190|1
35.41832|ac57ac390efa8412f80c8e0e438fb55f85a248dc|2.69|2015-03-04 19:35:00|80.749667378538092|3|7203663217|190|35.437367625817508|0|3|330|-80.762919|55|35.442529|EGGS|0.69|3|HT GRADE A LARGE EGGS 18 CT|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|35.465179900649026|00072036632173|EGGS FRESH|DAIRY|-80.746334|80.74633811067487|471|1
35.41832|4eaf91ee2478ea95a59617610e27d56f95875c20|1.99|2014-12-06 16:58:00|1.4102725052409182|3|7203600004|190|0.6181662995249579|0|1|1026|-80.746334|162|35.41832|WHEAT|0.0|7|HT HONEY WHEAT BRD|d7d54ae57897e7eccd6a0643cec77514075147af|1.3161449659704718|0.61833652052202714|00072036000040|SLICED BREAD|COMMERCIAL BAKERY|-80.746334|1.409289387215043|190|1
35.103409|b0f9f278f3d1eaeb453b0bdae1f70c6f5c0ae09b|3.29|2015-01-09 19:53:00|1.4132775322775095|4|2840018382|88|0.6126700657242101|0|58|201|-80.992182|31|35.103409|POTATO CHIPS|0.29|1|BAKED RUFFLES REGULAR|d8122272c740cad216fc6c038a5e0bceb6f36cac|4.083641674536447|0.61177642288969325|00028400184793|SNACKS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|3e92e2c6ac7ab8bad4eb4cbe8dd7cf804d19f880|3.29|2014-10-19 17:57:00|80.992238315890603|4|2840018382|88|35.162508618182244|0|22|201|-80.97058|31|35.03469|POTATO CHIPS|0.79|1|BAKED RUFFLES REGULAR|d8122272c740cad216fc6c038a5e0bceb6f36cac|4.083641674536447|35.131650835559327|00028400184793|SNACKS|G1 GROCERY|-80.992182|80.992226625110703|82|1
35.103409|afa506530778145cb9f8b5a28893ae01463309c6|3.29|2015-02-07 12:47:00|80.992238315890603|4|2840014741|88|35.162508618182244|0|22|205|-80.97058|31|35.03469|REMAINING SNACKS|0.79|1|SUNCHIPS REGULAR|d8122272c740cad216fc6c038a5e0bceb6f36cac|4.083641674536447|35.131650835559327|00028400147415|SNACKS|G1 GROCERY|-80.992182|80.992226625110703|82|1
35.103409|163a24c8bd947957fa9a5f8b417566b66c2694f0|4.19|2014-11-20 18:59:00|1.4132775322775095|4|2100000201|88|0.6126700657242101|0|58|317|-80.992182|52|35.103409|CHUNK AND BAR CHEESE|1.69|3|KRAFT NY EXTRA SHARP CHEESE|d8122272c740cad216fc6c038a5e0bceb6f36cac|4.083641674536447|0.61177642288969325|00021000001989|CHEESE|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|1098e18d0181c63ad216f87862e7ba7798535441|8.55|2015-02-21 17:42:00|1.4132775322775095|4|7510121065|88|0.6126700657242101|0|58|37|-80.992182|10|35.103409|PODS/CUPS/SINGLES|2.56|1|FOLGER GOURM CARM DRIZLE K-CUP|d8122272c740cad216fc6c038a5e0bceb6f36cac|4.083641674536447|0.61177642288969325|00025500201061|COFFEE|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|3a1a6841ba760056946dcc0279fee9210199df7d|5.58|2015-03-08 14:23:00|1.4132775322775095|4|7173000720|88|0.6126700657242101|0|58|150|-80.992182|23|35.103409|NOODLES/DUMPLINGS-DRY|1.4|1|NO YOLKS DUMPLINGS|d8122272c740cad216fc6c038a5e0bceb6f36cac|4.083641674536447|0.61177642288969325|00071730007201|PASTA|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|3bc13292fd7bbb61e7dc6defe907ba970b284108|6.9399999999999995|2014-12-14 14:09:00|1.4132775322775095|4|20165500000|88|0.6126700657242101|0|58|297|-80.992182|49|35.103409|GROUND BEEF|0.0|2|HT PREMIUM GRND BEEF 80% LEAN|d8122272c740cad216fc6c038a5e0bceb6f36cac|4.083641674536447|0.61177642288969325|00201655000005|BEEF|MEAT|-80.992182|1.413580244274486|88|2
35.103409|c0a14448100245c2c32bc8dc87a1419f979cc2d8|7.62|2015-02-15 17:59:00|1.4132775322775095|4|20165500000|88|0.6126700657242101|0|58|297|-80.992182|49|35.103409|GROUND BEEF|0.0|2|HT PREMIUM GRND BEEF 80% LEAN|d8122272c740cad216fc6c038a5e0bceb6f36cac|4.083641674536447|0.61177642288969325|00201655000005|BEEF|MEAT|-80.992182|1.413580244274486|88|2
35.103409|1c7ab3585b1cc602a76aa1664ed55a072dc53b23|0.25|2014-11-28 21:37:00|1.4132775322775095|4|4178900211|88|0.6126700657242101|0|58|1203|-80.992182|33|35.103409|RAMEN|0.0|1|MARUCHAN RAMEN CHICKEN|d8122272c740cad216fc6c038a5e0bceb6f36cac|4.083641674536447|0.61177642288969325|00041789002113|SOUP|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|7b89298263daf681a99424ea327565bba1e2dbc8|3.79|2015-01-24 18:31:00|80.992238315890603|4|4400002854|88|35.162508623604175|0|22|1248|-80.994596|12|35.061685|SANDWICH COOKIES|0.29|1|OREO DOUBLE STUFF|d8122272c740cad216fc6c038a5e0bceb6f36cac|4.083641674536447|35.131650835559327|00044000028541|COOKIES|G1 GROCERY|-80.992182|80.992214143493342|475|1
35.103409|0c4a1a267b81398515874e21cf9d3fca869102a0|3.99|2014-12-26 15:26:00|80.992238315890603|4|4400002854|88|35.162508618182244|0|22|1248|-80.97058|12|35.03469|SANDWICH COOKIES|1.49|1|OREO DOUBLE STUFF|d8122272c740cad216fc6c038a5e0bceb6f36cac|4.083641674536447|35.131650835559327|00044000028541|COOKIES|G1 GROCERY|-80.992182|80.992226625110703|82|1
35.103409|61c0365bf473780bb53066418b20db466e4c66ed|2.69|2014-11-16 16:37:00|1.4132775322775095|4|7294570544|88|0.6126700657242101|0|58|1025|-80.992182|162|35.103409|WHITE|0.2|7|SL S&S  W.G. WHITE BREAD|d8122272c740cad216fc6c038a5e0bceb6f36cac|4.083641674536447|0.61177642288969325|00072945705449|SLICED BREAD|COMMERCIAL BAKERY|-80.992182|1.413580244274486|88|1
35.103409|f9f49ea04bb0324a34eaad5f2424f6d2ab98e0c8|2.69|2015-01-04 16:03:00|1.4132775322775095|4|7294570544|88|0.6126700657242101|0|58|1025|-80.992182|162|35.103409|WHITE|0.0|7|SL S&S  W.G. WHITE BREAD|d8122272c740cad216fc6c038a5e0bceb6f36cac|4.083641674536447|0.61177642288969325|00072945705449|SLICED BREAD|COMMERCIAL BAKERY|-80.992182|1.413580244274486|88|1
35.103409|b7706585bbc33dc2da5389054e59a3fc7c62a817|2.59|2015-02-01 14:17:00|1.4132775322775095|4|1480000034|88|0.6126700657242101|0|58|128|-80.992182|20|35.103409|APPLE JUICE-SHELF|0.0|1|MOTTS FOR TOTS APPLE JUICE|d8122272c740cad216fc6c038a5e0bceb6f36cac|4.083641674536447|0.61177642288969325|00014800318203|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|df2c0979237b39389737f9679697207908f15e78|2.15|2014-11-01 17:39:00|80.992238315890603|4|3800030110|88|35.162508618182244|0|22|44|-80.97058|6|35.03469|TOASTER PASTRIES-SHELF STABLE|0.15|1|KELL POPTART COOKIES CREME|d8122272c740cad216fc6c038a5e0bceb6f36cac|4.083641674536447|35.131650835559327|00038000235948|BREAKFAST FOODS|G1 GROCERY|-80.992182|80.992226625110703|82|1
35.103409|066b0b4ad665076a10fc13fb984b3327cad918f4|3.59|2014-11-08 15:36:00|80.992238315890603|4|4127100908|88|35.162508618182244|0|22|341|-80.97058|57|35.03469|CREAMERS|0.59|3|I/O ITNAT'L WHITE CHOC RASP|d8122272c740cad216fc6c038a5e0bceb6f36cac|4.083641674536447|35.131650835559327|00041271009088|MILK|DAIRY|-80.992182|80.992226625110703|82|1
35.103409|8edee08b7a6724662e4d19d676f04809e4b2f4be|1.99|2015-02-03 19:25:00|1.4132775322775095|4|4142001998|88|0.6126700657242101|0|58|727|-80.992182|7|35.103409|SEASONAL CANDY-SINGLE FAC|1.0|1|I/O(V15)BRACH SM CONV HEARTS|d8122272c740cad216fc6c038a5e0bceb6f36cac|4.083641674536447|0.61177642288969325|00041420019982|CANDY|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|2c70ed7fd161cd20554d9a1a22380459de001419|3.99|2015-02-12 17:30:00|1.4132775322775095|4|7316826801|88|0.6126700657242101|0|58|6975|-80.992182|1600|35.103409|VALENTINE CARDS IMP|1.0|18|WOODLAND CREATURES VAL CARDS|d8122272c740cad216fc6c038a5e0bceb6f36cac|4.083641674536447|0.61177642288969325|00073168268018|SEASONAL MERCHANDISE|GM|-80.992182|1.413580244274486|88|1
35.103409|d686b6708a89d30157e8313be3fe3c8035f8d4b8|7.79|2015-01-10 13:11:00|80.992238315890603|4|30045027125|88|35.162508618182244|0|22|4195|-80.97058|1200|35.03469|COUGH & COLD REMEDY-ADULT|1.8|17|TYL COLD HEAD CONG CAPLETS|d8122272c740cad216fc6c038a5e0bceb6f36cac|4.083641674536447|35.131650835559327|00300450261250|COUGH/COLD/SINUS|HBC|-80.992182|80.992226625110703|82|1
35.103409|aaf4c5d44bfd3a996362728c6f4dbf4ed12bfa96|13.58|2014-12-26 15:27:00|80.992238315890603|4|1200080994|88|35.162508618182244|0|22|55|-80.97058|8|35.03469|REGULAR|3.6|23|DR. PEPPER FRIDGEMATE|d8122272c740cad216fc6c038a5e0bceb6f36cac|4.083641674536447|35.131650835559327|00078000082166|CARBONATED BEVERAGES|BEVERAGE|-80.992182|80.992226625110703|82|2
35.103409|603db14a3cb4b01237dd5d85b2410afa56667b02|7.99|2015-03-07 19:14:00|80.992238315890603|4|63598560611|88|35.162508618182244|0|22|464|-80.97058|84|35.03469|HARD LEMONADE|0.0|16|MIKES CRANBERRY LEMONADE 6PK|d8122272c740cad216fc6c038a5e0bceb6f36cac|4.083641674536447|35.131650835559327|00635985606116|SPECIALTY|BEER|-80.992182|80.992226625110703|82|1
35.323246|08a4f518a2c96bcdeb88ce992bd9645698739c7a|23.7|2015-01-11 12:44:00|1.4102725052409182|4|20896900000|166|0.6165069451919168|0|1|657|-80.945176|201|35.323246|STR MDE VALUE ADD POLTRY|13.56|2|HNY GINGER MARINATED CHKN BRST|debab8cb01b12495d1fb25d083e0202924ab0219|3.0895476464389655|0.61833652052202714|00208969000004|POULTRY|MEAT|-80.945176|1.4127598348062935|166|1
35.323246|872ac204c28f0d58310b8153030c22f784858613|2.29|2014-10-10 13:07:00|1.4102725052409182|4|1900008501|166|0.6165069451919168|0|1|50|-80.945176|7|35.323246|PEG CANDY|0.29|1|LIFESAVERS GUMMI WILDBERRIES|debab8cb01b12495d1fb25d083e0202924ab0219|3.0895476464389655|0.61833652052202714|00019000083449|CANDY|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|5fbd98dbea613db4af97a146bcb441454019b0fd|3.98|2015-02-10 13:51:00|1.4102725052409182|4|7680828073|166|0.6165069451919168|0|1|149|-80.945176|23|35.323246|WHSE PASTA CORE|0.49|1|BARILLA PASTA RIGATONI|debab8cb01b12495d1fb25d083e0202924ab0219|3.0895476464389655|0.61833652052202714|00076808502947|PASTA|G1 GROCERY|-80.945176|1.4127598348062935|166|2
35.323246|72805bef0f837826410027f370251d80ab498a5c|1.37|2014-10-19 10:52:00|1.4102725052409182|4|1122509483|166|0.6165069451919168|0|1|192|-80.945176|30|35.323246|COOKING SPRAYS|0.0|1|VALU TME VEGETABLE COOKNG SPRY|debab8cb01b12495d1fb25d083e0202924ab0219|3.0895476464389655|0.61833652052202714|00011225094835|SHORTENING/OIL|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|9f5566586a37c7cf5bd7c5414559c78dc06411b7|38.97|2015-02-13 10:45:00|1.4102725052409182|4|7203695587|166|0.6165069451919168|0|1|1707|-80.945176|387|35.323246|MESSAGE|9.0|14|12 INCH MESSAGE COOKIE|debab8cb01b12495d1fb25d083e0202924ab0219|3.0895476464389655|0.61833652052202714|00072036955876|COOKIES|BAKERY|-80.945176|1.4127598348062935|166|3
35.323246|1b688380aa1e795de27d4a159c3c767dea291c57|2.98|2015-02-27 13:33:00|1.4102725052409182|4|7618316363|166|0.6165069451919168|0|1|99|-80.945176|32|35.323246|LIQUID TEA|0.98|1|SNAPPLE KIWI STRAWBERRY|debab8cb01b12495d1fb25d083e0202924ab0219|3.0895476464389655|0.61833652052202714|00076183163634|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.945176|1.4127598348062935|166|2
35.323246|42e061a028eb5cda80768d08698fa63f9ec305b5|15.96|2015-02-10 14:27:00|1.4102725052409182|4|7203688076|166|0.6165069451919168|0|1|523|-80.945176|64|35.323246|FRESH POTATOES|1.96|4|HT RUSSET POTATO 5LB BAG|debab8cb01b12495d1fb25d083e0202924ab0219|3.0895476464389655|0.61833652052202714|00072036880765|FRESH PRODUCE|PRODUCE|-80.945176|1.4127598348062935|166|4
35.323246|201329c11c341b864ab177684224e20b22d5b362|9.99|2015-02-02 14:01:00|1.4102725052409182|4|3700086527|166|0.6165069451919168|0|1|427|-80.945176|72|35.323246|NFS-TOILET TISSUE|4.0|1|CHARMIN BATH ULTRA SOFT 6MR|debab8cb01b12495d1fb25d083e0202924ab0219|3.0895476464389655|0.61833652052202714|00037000868019|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|699179988b04d2965ca8764e8b169cce13b1a783|7.97|2015-01-08 14:33:00|1.4102725052409182|4|3700009614|166|0.6165069451919168|0|1|3774|-80.945176|1070|35.323246|CLINICAL-FEMALE|0.0|17|SECRET ADV SOLID SERENCTRS|debab8cb01b12495d1fb25d083e0202924ab0219|3.0895476464389655|0.61833652052202714|00037000850519|DEODORANT|HBC|-80.945176|1.4127598348062935|166|1
35.323246|188424e8a92249bf1c611bbb354fdc4c473ae92b|7.79|2015-01-02 17:51:00|80.945255278477163|4|30045027125|166|35.367958781918247|0|13|4236|-80.782849|1200|35.372142|DEX ADULT/CHILDREN|0.0|17|TYL SEVERE COLD/FLU CAPLETS|debab8cb01b12495d1fb25d083e0202924ab0219|3.0895476464389655|35.37387923947206|00300450270269|COUGH/COLD/SINUS|HBC|-80.945176|80.945244231968658|122|1
35.323246|3df01c4adb3fec294087056361ddcf2cb02581a8|8.99|2014-09-12 14:23:00|1.4102725052409182|4|76211120604|166|0.6165069451919168|0|1|36|-80.945176|10|35.323246|PREMIUM GROUND|2.0|1|STARBUCKS ITALIAN ROAST GROUND|debab8cb01b12495d1fb25d083e0202924ab0219|3.0895476464389655|0.61833652052202714|00762111622853|COFFEE|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|19d73cb1c2a3dbfaddf6af81d9b77e55742be4aa|1.0|2015-01-16 08:47:00|80.945255278477163|4|4000000435|166|35.3679588117256|0|13|47|-80.810056|7|35.219587|REGISTER BARS|0.0|1|(FE)M&M PEANUT CANDY|debab8cb01b12495d1fb25d083e0202924ab0219|3.0895476464389655|35.37387923947206|00040000000327|CANDY|G1 GROCERY|-80.945176|80.945201480489615|401|1
35.323246|8282b90f9b115ee5744e156d96cf3a02ecef83d5|29.58|2015-03-08 19:57:00|1.4102725052409182|4|3700086522|166|0.6165069451919168|0|1|427|-80.945176|72|35.323246|NFS-TOILET TISSUE|5.6|1|CHARMIN BATH ULTRA SOFT 9MR|debab8cb01b12495d1fb25d083e0202924ab0219|3.0895476464389655|0.61833652052202714|00037000868033|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.945176|1.4127598348062935|166|2
35.323246|de9ae5d854c1c4f8e48160c4b555b630a8dbbb16|5.49|2015-01-11 12:32:00|1.4102725052409182|4|8500001846|166|0.6165069451919168|0|1|9925|-80.945176|883|35.323246|NFS-ECONOMY GLASS|0.0|13|TISDALE SWEET RED|debab8cb01b12495d1fb25d083e0202924ab0219|3.0895476464389655|0.61833652052202714|00085000018460|ECONOMY (GLASS 3L & UP)|WINE|-80.945176|1.4127598348062935|166|1
35.323246|b943d18fa2dd5be48b4be199240835545d159db9|5.98|2015-01-02 13:47:00|1.4102725052409182|4|5208333816|166|0.6165069451919168|0|1|1976|-80.945176|475|35.323246|COLD PIZZA OTHER|0.0|6|PREMIUM PIZZA DOUGH BALLS|debab8cb01b12495d1fb25d083e0202924ab0219|3.0895476464389655|0.61833652052202714|00052083338167|PIZZA|DELI|-80.945176|1.4127598348062935|166|2
35.323246|2f121c25b3406720dbad67b92dd330671bf87e86|1.19|2015-02-10 13:52:00|1.4102725052409182|4|7203653022|166|0.6165069451919168|0|1|1273|-80.945176|50|35.323246|BAG VEG NON STEAM|0.0|5|HT BROCCOLI CUTS|debab8cb01b12495d1fb25d083e0202924ab0219|3.0895476464389655|0.61833652052202714|00072036530721|VEGETABLES-FROZEN|FROZEN|-80.945176|1.4127598348062935|166|1
35.219587|d0c116c835e005bf2e94177b380fbd2f1ddd259e|1.34|2014-10-23 12:53:00|80.810069425230125|4|7203670897|401|35.259897368416716|0|23|214|-80.995484|33|35.444064|BROTH|0.34|1|HT FF BEEF BROTH|df39f4df1b401289af1c63c58339b6330006f515|2.785352203287377|35.240679762029046|00072036708991|SOUP|G1 GROCERY|-80.810056|80.810129537296135|121|2
35.219587|d2b33f2fdc8dfb053ac0e259ff36e335b95ed83e|3.1799999999999997|2014-10-05 16:54:00|80.810069425230125|4|1708289781|401|35.259897368416716|0|23|206|-80.995484|31|35.444064|FRONT END SNACKS|0.0|1|JLINKS SASQUATCH ORIG BIG STK|df39f4df1b401289af1c63c58339b6330006f515|2.785352203287377|35.240679762029046|00017082897817|SNACKS|G1 GROCERY|-80.810056|80.810129537296135|121|2
35.219587|a714a0eee0eb82c1724e709e8737ddade55eb4e1|4.99|2014-10-05 16:57:00|80.810069425230125|4|67569050122|401|35.259897368416716|0|23|3919|-80.995484|1075|35.444064|DISPOSABLE RAZOR-WOMEN|2.0|17|NOXEMA 12CT DISPOSABLE RAZORS|df39f4df1b401289af1c63c58339b6330006f515|2.785352203287377|35.240679762029046|00675690501221|SHAVING NEEDS/MEN HAIR|HBC|-80.810056|80.810129537296135|121|1
35.219587|fc8f436e7572a3b69f55edfaadc7de3829f9316c|4.99|2014-09-30 13:03:00|80.810069425230125|4|67569050122|401|35.259897368416716|0|23|3919|-80.995484|1075|35.444064|DISPOSABLE RAZOR-WOMEN|2.0|17|NOXEMA 12CT DISPOSABLE RAZORS|df39f4df1b401289af1c63c58339b6330006f515|2.785352203287377|35.240679762029046|00675690501221|SHAVING NEEDS/MEN HAIR|HBC|-80.810056|80.810129537296135|121|1
35.219587|f12fac172538594cec90d57c5835fffeca066a8c|6.49|2014-11-19 10:16:00|80.810069425230125|4|1200080994|401|35.259897387220398|0|23|55|-80.737839|8|35.297134|REGULAR|1.5|23|CF PEPSI FRIDGEMATE|df39f4df1b401289af1c63c58339b6330006f515|2.785352203287377|35.240679762029046|00012000810022|CARBONATED BEVERAGES|BEVERAGE|-80.810056|80.810111992540072|258|1
35.219587|31da0c8407675c1f9ab3a7fc5381ea638b1cd7a3|1.69|2014-11-18 15:40:00|80.810069425230125|4|3660207290|401|35.259897368416716|0|23|4207|-80.995484|1200|35.444064|COUGH DROP-ADULT|0.84|17|RICOLA NATURAL HERB -07917|df39f4df1b401289af1c63c58339b6330006f515|2.785352203287377|35.240679762029046|00036602079175|COUGH/COLD/SINUS|HBC|-80.810056|80.810129537296135|121|1
35.43259|6f054b136e5230aa6576ee89001c86ebb31a6cc1|3.38|2015-01-16 14:18:00|1.4057311447477159|3|65153806700|202|0.6184153580092175|0|52|99|-80.605588|32|35.43259|LIQUID TEA|0.0|1|SWT LEAF HONEY GREEN TEA|e0e89f173013ea67aa270afbacc8f6a37face17e|10.34758948264388|0.6209993146566879|00651538067012|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.605588|1.406832906106031|202|2
35.43259|926e0fc31625d8793ec96428f0ec41f216a33af3|1.58|2014-11-11 10:32:00|80.606823361882718|3||202|35.582343017272365|0|57|532|-80.66939|64|35.28326|FRESH CUCUMBERS|0.2|4|COO CUCUMBERS S/S|e0e89f173013ea67aa270afbacc8f6a37face17e|10.34758948264388|35.500309569604553|00204062000002|FRESH PRODUCE|PRODUCE|-80.605588|80.605927585243435|46|2
35.43259|bd3f8dd3541e44b4d2c3597ed7656a2c7c42ca41|1.95|2014-10-14 13:43:00|80.606823361882718|3|4470002410|202|35.582343255719771|0|57|659|-80.662946|103|35.412407|CHILDRENS LUNCH SNACKS|0.0|19|BASIC LUNCHABLE TURKEY STACKER|e0e89f173013ea67aa270afbacc8f6a37face17e|10.34758948264388|35.500309569604553|00044700360019|LUNCH SNACKS|CASE READY MEATS|-80.605588|80.605674865811338|68|1
35.43259|b3f0d61aaad55c7cc0b1552630cda61dad27f0af|0.99|2014-12-22 16:03:00|80.606823361882718|3|4300020001|202|35.582343017272365|0|57|93|-80.66939|14|35.28326|GELATIN MIXES|0.24|1|KOOL AID GELATIN CHERRY|e0e89f173013ea67aa270afbacc8f6a37face17e|10.34758948264388|35.500309569604553|00043000063880|DESSERTS/GELS/SYRUPS|G1 GROCERY|-80.605588|80.605927585243435|46|1
35.43259|a5af577312f05ae173a19269eb2c9b64c986a93b|4.99|2014-10-26 11:42:00|80.606823361882718|3||202|35.582343255719771|0|57|500|-80.662946|64|35.412407|FRESH APPLES|0.55|4|RED DEL APPLE, WA  48|e0e89f173013ea67aa270afbacc8f6a37face17e|10.34758948264388|35.500309569604553|00233284000002|FRESH PRODUCE|PRODUCE|-80.605588|80.605674865811338|68|1
35.43259|cb71abc59b46b8cfcee1969273a7127319154548|24.28|2015-01-29 14:16:00|80.606823361882718|3|20138900000|202|35.582343255719771|0|57|296|-80.662946|49|35.412407|RANCHER BEEF|6.75|2|BEEF TENDERLOIN FILET MIGNON|e0e89f173013ea67aa270afbacc8f6a37face17e|10.34758948264388|35.500309569604553|00201389000005|BEEF|MEAT|-80.605588|80.605674865811338|68|2
35.43259|9f9a26f99bf057af229dba2eac686f43053b2501|7.18|2014-10-07 14:29:00|80.606823361882718|3|20252400000|202|35.582343255719771|0|57|299|-80.662946|49|35.412407|ANGUS BEEF|0.0|2|ANGUS BF TENDERIZED CUBED STK|e0e89f173013ea67aa270afbacc8f6a37face17e|10.34758948264388|35.500309569604553|00202524000003|BEEF|MEAT|-80.605588|80.605674865811338|68|2
35.43259|c56f1443efdbf23b92399c2cd482588dde630da8|4.99|2014-11-18 14:29:00|80.606823361882718|3|4950800823|202|35.582343255719771|0|57|1980|-80.662946|480|35.412407|CHOCOLATES|1.0|6|DARK CHOC PRETZEL CRISPS|e0e89f173013ea67aa270afbacc8f6a37face17e|10.34758948264388|35.500309569604553|00049508008231|DRY GOODS|DELI|-80.605588|80.605674865811338|68|1
35.43259|a7ab5367a63c0bee3b730108b5ec8eceb4451e4c|27.96|2015-01-31 15:58:00|80.606823361882718|3|4900002890|202|35.582343017272365|0|57|55|-80.66939|8|35.28326|REGULAR|6.99|23|CLASSIC 12OZ 12PK FRIDGE CAN|e0e89f173013ea67aa270afbacc8f6a37face17e|10.34758948264388|35.500309569604553|00049000028904|CARBONATED BEVERAGES|BEVERAGE|-80.605588|80.605927585243435|46|4
35.23102|a2be286be7c9d452fe770feda616592bfaee8e03|5.07|2014-10-25 11:15:00|80.843809562956082|4||205|35.256925665302894|0|37|524|-80.810056|64|35.219587|FRESH PROD FRESH ONIONS|0.0|4|COO VIDALIA SWEET BULB ONION|e423eef1085fdde6ed985fd515033f0e9aa71e6c|1.7900189135238365|35.255745041786184|00204824000004|FRESH PRODUCE|PRODUCE|-80.8438|80.843801079620974|401|3
35.23102|cc296d5692c3e0b52eda00c036d5f9b5363b2191|0.97|2015-01-22 11:14:00|80.843809562956082|4|7203608052|205|35.256925646665785|0|37|76|-80.780702|11|35.318911|MEAT SAUCES|0.0|1|HT WORCESTERSHIRE SAUCE|e423eef1085fdde6ed985fd515033f0e9aa71e6c|1.7900189135238365|35.255745041786184|00072036080523|CONDIMENTS|G1 GROCERY|-80.8438|80.843838063827206|167|1
35.23102|97e361a9fd33b43eafe5e80c0c6238cc642108fc|4.59|2014-12-21 16:02:00|80.843809562956082|4|7140300004|205|35.256925646596507|0|37|67|-80.814133|10|35.333742|SOLUBLE INSTANT|0.0|1|FERRARA ESPRESSO INSTANT|e423eef1085fdde6ed985fd515033f0e9aa71e6c|1.7900189135238365|35.255745041786184|00071403000041|COFFEE|G1 GROCERY|-80.8438|80.843838134456263|472|1
35.23102|ecf544a4cb711c4a92d45d8443b4a817ca66b182|2.98|2015-01-27 11:10:00|80.843809562956082|4|85245300200|205|35.256925646665785|0|37|508|-80.780702|64|35.318911|FRESH GRAPEFRUIT|0.0|4|RED GRAPEFRUIT 3LB BAG|e423eef1085fdde6ed985fd515033f0e9aa71e6c|1.7900189135238365|35.255745041786184|00033383911120|FRESH PRODUCE|PRODUCE|-80.8438|80.843838063827206|167|2
35.23102|58f602d3c01453c346f642f4991dc9efd9d14a4b|7.58|2015-03-04 11:07:00|80.843809562956082|4|4850002013|205|35.256925646665785|0|37|335|-80.780702|56|35.318911|ORANGE JUICE-REGRIGERATED|1.58|3|TROPICANA PP ORIGINAL|e423eef1085fdde6ed985fd515033f0e9aa71e6c|1.7900189135238365|35.255745041786184|00048500301029|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.8438|80.843838063827206|167|2
35.23102|3d6424a27bfef0ebdf0beb90b5950e4710660cbd|0.75|2014-10-04 13:21:00|80.843809562956082|4|7203641160|205|35.256925646665785|0|37|247|-80.780702|39|35.318911|VEGETABLES-FLANKER|0.0|1|HT BEETS CUT|e423eef1085fdde6ed985fd515033f0e9aa71e6c|1.7900189135238365|35.255745041786184|00072036410818|VEGETABLES-CAN/JAR|G1 GROCERY|-80.8438|80.843838063827206|167|1
35.23102|b3003a0d847b644570f79794d480fd3cbb48e56d|3.85|2014-12-24 13:53:00|80.843809562956082|4|2100060464|205|35.256925646665785|0|37|315|-80.780702|52|35.318911|CHEESE-PROCESSED-SLICED|0.0|3|KRAFT WHITE AMERICAN|e423eef1085fdde6ed985fd515033f0e9aa71e6c|1.7900189135238365|35.255745041786184|00021000604654|CHEESE|DAIRY|-80.8438|80.843838063827206|167|1
35.43259|c3b6072052cfa531d34a21975c4e4b95b6093897|5.99|2014-11-17 09:48:00|1.4057311447477159|4|7203695643|202|0.6184153580092175|0|52|1663|-80.605588|381|35.43259|CREME CAKE|0.0|14|44 OZ CHOC CREME CAKE|e493b47d791a206988bd474918d6e2ae3732aeb7|3.7766321979927717|0.6209993146566879|00072036956644|CAKES|BAKERY|-80.605588|1.406832906106031|202|1
35.43259|9cd1599d8434c487a8a96969575b6d13dbcaca32|0.51|2014-12-11 13:08:00|80.606823361882718|4||202|35.487246494474263|0|57|502|-80.662946|64|35.412407|FRESH BANANAS|0.0|4|BANANAS, YELLOW|e493b47d791a206988bd474918d6e2ae3732aeb7|3.7766321979927717|35.500309569604553|00204011000008|FRESH PRODUCE|PRODUCE|-80.605588|80.605619666494704|68|1
35.43259|47a8b51581b5dd1ce92653ad53f22cd147a0588b|7.99|2015-02-25 12:04:00|1.4057311447477159|4|8500000704|202|0.6184153580092175|0|52|9925|-80.605588|883|35.43259|NFS-ECONOMY GLASS|0.0|13|CARLO ROSSI CHABLIS 1.5L|e493b47d791a206988bd474918d6e2ae3732aeb7|3.7766321979927717|0.6209993146566879|00085000007044|ECONOMY (GLASS 3L & UP)|WINE|-80.605588|1.406832906106031|202|1
35.43259|2c20688f28954ddbc60f78f6671d3005c613fd6b|4.99|2014-11-17 09:49:00|1.4057311447477159|4|20165500000|202|0.6184153580092175|0|52|297|-80.605588|49|35.43259|GROUND BEEF|0.0|2|HT PREMIUM GRND BEEF 80% LEAN|e493b47d791a206988bd474918d6e2ae3732aeb7|3.7766321979927717|0.6209993146566879|00201655000005|BEEF|MEAT|-80.605588|1.406832906106031|202|1
35.43259|cbfd9a29d00943afbd9b5154e99bb87bc5488331|7.99|2014-11-20 11:31:00|1.4057311447477159|4|8500000480|202|0.6184153580092175|0|52|9925|-80.605588|883|35.43259|NFS-ECONOMY GLASS|0.0|13|CARLO ROSSI CHARDONNAY 1.5L|e493b47d791a206988bd474918d6e2ae3732aeb7|3.7766321979927717|0.6209993146566879|00085000004807|ECONOMY (GLASS 3L & UP)|WINE|-80.605588|1.406832906106031|202|1
35.43259|06dbab393de95442f7b8b6cbdd5e8fa4dc175ce6|3.89|2015-02-23 09:30:00|1.4057311447477159|4|3010054073|202|0.6184153580092175|0|52|1249|-80.605588|12|35.43259|CHOCOLATE CHIP COOKIES|1.94|1|CHIPS DELUXE RAINBOW|e493b47d791a206988bd474918d6e2ae3732aeb7|3.7766321979927717|0.6209993146566879|00030100100379|COOKIES|G1 GROCERY|-80.605588|1.406832906106031|202|1
35.43259|c80ddaa97158daa16bbdc74bbcda3736327878c7|1.39|2014-12-19 10:59:00|1.4057311447477159|4|7203602056|202|0.6184153580092175|0|52|78|-80.605588|11|35.43259|MUSTARD|0.7|1|HT MUSTARD YELLOW 14 OZ|e493b47d791a206988bd474918d6e2ae3732aeb7|3.7766321979927717|0.6209993146566879|00072036020567|CONDIMENTS|G1 GROCERY|-80.605588|1.406832906106031|202|1
35.43259|eb2e536f0ebe7200035ee4f4b46263ce3e5d1a01|8.0|2014-09-14 12:03:00|1.4057311447477159|4|84115200732|202|0.6184153580092175|0|52|1165|-80.605588|87|35.43259|NFS-FRESH CONSUMER BUNCH|0.0|9|BUNCH- 3/$12 DAISY BUNCHES|e493b47d791a206988bd474918d6e2ae3732aeb7|3.7766321979927717|0.6209993146566879|00841152007321|FLORAL|FLORAL|-80.605588|1.406832906106031|202|2
35.43259|e2b9e02f2fd96a3a95caf23446958548bb5d7e84|11.98|2014-12-15 11:10:00|1.4057311447477159|4|7203695643|202|0.6184153580092175|0|52|1663|-80.605588|381|35.43259|CREME CAKE|0.0|14|44 OZ MARBLE CREME CAKE|e493b47d791a206988bd474918d6e2ae3732aeb7|3.7766321979927717|0.6209993146566879|00072036956637|CAKES|BAKERY|-80.605588|1.406832906106031|202|2
35.43259|568a97ac9a75dbc3e9b8b77cc08472a2c6db7d3d|5.99|2014-12-15 11:11:00|1.4057311447477159|4|7203695643|202|0.6184153580092175|0|52|1663|-80.605588|381|35.43259|CREME CAKE|0.0|14|44 OZ VANILLA CREME CAKE|e493b47d791a206988bd474918d6e2ae3732aeb7|3.7766321979927717|0.6209993146566879|00072036956439|CAKES|BAKERY|-80.605588|1.406832906106031|202|1
35.667941|3d72eff4dfc8e245a10ce648afa02aadb9a17cd0|7.78|2015-01-04 11:59:00|1.4057311447477159|3|5450019352|178|0.6225230078570788|0|52|359|-80.497332|101|35.667941|MEAT WIENERS|1.78|19|BALL PARK BUN SIZE MEAT FRANK|e7b6658229af085da8e586939d1319971ea11620|8.628164382726366|0.6209993146566879|00054500193274|WIENERS|CASE READY MEATS|-80.497332|1.4049434824709919|178|2
35.667941|feb34c38fd2a67b2b46d7ab3f99d432192d18630|1.49|2014-12-10 16:04:00|80.497482303704658|3|20406100000|178|35.792808932682277|0|6|525|-80.764523|64|35.341927|FRESH LETTUCE|0.0|4|ICEBERG LETTUCE|e7b6658229af085da8e586939d1319971ea11620|8.628164382726366|35.699188602026126|00033383650203|FRESH PRODUCE|PRODUCE|-80.497332|80.49804149348752|220|1
35.667941|0989ac76e50fe84d9ab462abebcb0d0794578d87|2.79|2015-01-21 13:06:00|80.497482303704658|3|1600015110|178|35.792808932682277|0|6|205|-80.764523|31|35.341927|REMAINING SNACKS|1.39|1|CHEX SNACK MIX - BOLD PARTY BL|e7b6658229af085da8e586939d1319971ea11620|8.628164382726366|35.699188602026126|00016000159402|SNACKS|G1 GROCERY|-80.497332|80.49804149348752|220|1
35.667941|939c34cd02b33b623056cdf2feff66bb855e4534|9.4|2014-09-18 15:55:00|80.497482303704658|3||178|35.792808932682277|0|6|503|-80.764523|64|35.341927|FRESH GRAPES|5.7|4|GREEN GRAPES, SEEDLESS 12/16|e7b6658229af085da8e586939d1319971ea11620|8.628164382726366|35.699188602026126|00204022000004|FRESH PRODUCE|PRODUCE|-80.497332|80.49804149348752|220|1
35.667941|49b9f9564584e8c6f0b8deb803f18a541a3e2560|3.25|2015-02-19 12:54:00|1.4057311447477159|3|7203656080|178|0.6225230078570788|0|52|318|-80.497332|52|35.667941|SHREDDED/GRATED CHEESE|0.0|3|HT SHREDDED MOZZ/PROVLONE|e7b6658229af085da8e586939d1319971ea11620|8.628164382726366|0.6209993146566879|00072036705174|CHEESE|DAIRY|-80.497332|1.4049434824709919|178|1
35.667941|a09c94084b6c5762708a98f0c3b7ead258195e3c|1.49|2014-11-21 18:00:00|1.4057311447477159|3|87218100501|178|0.6225230078570788|0|52|47|-80.497332|7|35.667941|REGISTER BARS|0.2|1|(FE)TURTLES 3PC|e7b6658229af085da8e586939d1319971ea11620|8.628164382726366|0.6209993146566879|00872181005019|CANDY|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|e4c6d365fda0d2fad9c04608a1959b9be8075c60|6.55|2014-12-07 12:34:00|1.4057311447477159|3|7570616502|178|0.6225230078570788|0|52|254|-80.497332|892|35.667941|PREMIUM PIZZA|0.57|5|PALERMOS HT PEPPERONI PIZZA|e7b6658229af085da8e586939d1319971ea11620|8.628164382726366|0.6209993146566879|00075706148035|FROZEN PIZZA|FROZEN|-80.497332|1.4049434824709919|178|1
35.667941|aca5ca159e6f1a574461dfebe0a7ab04d4b3f2e0|0.97|2015-02-25 16:37:00|80.497482303704658|3|7203688002|178|35.792808932682277|0|6|527|-80.764523|64|35.341927|FRESH CARROTS|0.0|4|HT WHOLE CARROTS 2LB BAG|e7b6658229af085da8e586939d1319971ea11620|8.628164382726366|35.699188602026126|00072036880024|FRESH PRODUCE|PRODUCE|-80.497332|80.49804149348752|220|1
35.667941|aa662c120552578c571f9698d71d58a8e78c943b|2.37|2015-03-07 16:05:00|1.4057311447477159|3|7203608050|178|0.6225230078570788|0|52|76|-80.497332|11|35.667941|MEAT SAUCES|0.0|1|HT STEAK SAUCE|e7b6658229af085da8e586939d1319971ea11620|8.628164382726366|0.6209993146566879|00072036080509|CONDIMENTS|G1 GROCERY|-80.497332|1.4049434824709919|178|1
35.667941|3732b40f4ecab036ba380ad4de94244df8102de8|6.55|2015-01-11 12:27:00|1.4057311447477159|3|7570616502|178|0.6225230078570788|0|52|254|-80.497332|892|35.667941|PREMIUM PIZZA|3.27|5|PALERMOS PEPPERONI PIZZA|e7b6658229af085da8e586939d1319971ea11620|8.628164382726366|0.6209993146566879|00075706165018|FROZEN PIZZA|FROZEN|-80.497332|1.4049434824709919|178|1
35.667941|b040088753d33614e2ef9044af0c0c116338966b|7.99|2014-11-23 12:34:00|1.4057311447477159|3|8857370002|178|0.6225230078570788|0|52|458|-80.497332|82|35.667941|CRAFT BEER|0.0|16|SHINER FAMILY REUNION 6PK|e7b6658229af085da8e586939d1319971ea11620|8.628164382726366|0.6209993146566879|00088573700022|DOMESTIC BEER|BEER|-80.497332|1.4049434824709919|178|1
35.667941|2f49ba58af8592fa1edb530f4e54ae0454ec7b87|3.49|2015-02-02 16:43:00|80.497482303704658|3|20455000000|178|35.792808932682277|0|6|542|-80.764523|64|35.341927|FRESH VEGETABLES REMAIN|0.0|4|BRUSSEL SPROUTS 1LB (RPC)|e7b6658229af085da8e586939d1319971ea11620|8.628164382726366|35.699188602026126|00094922577160|FRESH PRODUCE|PRODUCE|-80.497332|80.49804149348752|220|1
35.667941|cdaa82ff7d556179a588fcc2db53e430dc1dbc71|11.99|2014-11-17 12:25:00|1.4057311447477159|3|8769201103|178|0.6225230078570788|0|52|458|-80.497332|82|35.667941|CRAFT BEER|0.0|16|SAM ADAMS SEASONAL 12PK|e7b6658229af085da8e586939d1319971ea11620|8.628164382726366|0.6209993146566879|00087692011033|DOMESTIC BEER|BEER|-80.497332|1.4049434824709919|178|1
35.667941|2ae1d957ef2f1f47bbeae3ebe059564fa518f198|3.49|2014-11-07 09:49:00|80.497482303704658|3|2068500089|178|35.792809185197051|0|6|197|-80.8955|31|35.4437|POPPED POPCORN|0.99|1|CAPE COD SEA SALT POPCORN|e7b6658229af085da8e586939d1319971ea11620|8.628164382726366|35.699188602026126|00020685000874|SNACKS|G1 GROCERY|-80.497332|80.497970501392103|272|1
35.667941|5ea1bb8b9117803e225e7ec18d5abcfe0341fc94|5.13|2014-10-04 12:48:00|1.4057311447477159|3||178|0.6225230078570788|0|52|523|-80.497332|64|35.667941|FRESH POTATOES|1.19|4|COO SWEET POTATOES, BULK|e7b6658229af085da8e586939d1319971ea11620|8.628164382726366|0.6209993146566879|00204091000004|FRESH PRODUCE|PRODUCE|-80.497332|1.4049434824709919|178|1
35.23102|fff8fd27d440d3e6ba85492777cbf51fc424494a|2.5|2015-03-01 18:04:00|80.843945456961976|2|78142100610|205|35.233522162802032|0|59|1601|-80.70901|371|35.17335|BRANDED BREAD|1.51|14|LA BREA WHEAT BAGUETTE|e829a323ff38f07bbea130697026b25eeedc25a3|0.17289340712391948|35.232478750868765|00781421521182|BREAD|BAKERY|-80.8438|80.843800034139889|174|1
35.23102|cdcdaf90d3e460550006d1a18d106b48c4370920|4.99|2015-02-07 12:32:00|80.843945456961976|2|6827493471|205|35.233522162802032|0|59|31|-80.70901|4|35.17335|NON CARBONATED WATER|2.0|1|NESTLE PURE LIFE .5L 24PK|e829a323ff38f07bbea130697026b25eeedc25a3|0.17289340712391948|35.232478750868765|00068274934711|BOTTLED WATER|G1 GROCERY|-80.8438|80.843800034139889|174|1
35.23102|714dde64e829d34645a34d5f674fc34c5d4b5778|8.21|2015-01-28 14:29:00|80.843945456961976|2|20249700000|205|35.233522162802032|0|59|297|-80.70901|49|35.17335|GROUND BEEF|0.41|2|NY STRIP STEAKBURGER 80% LEAN|e829a323ff38f07bbea130697026b25eeedc25a3|0.17289340712391948|35.232478750868765|00202497000000|BEEF|MEAT|-80.8438|80.843800034139889|174|1
35.23102|f17b589db981ba7eda7612fc9250871b1b243a46|7.39|2014-10-10 17:15:00|80.843945456961976|2|3500068048|205|35.233522162802032|0|59|4056|-80.70901|1080|35.17335|TOOTH BRUSH-PREMIUM|2.39|17|COLG 360 OPTC WH TB CP SFT 247|e829a323ff38f07bbea130697026b25eeedc25a3|0.17289340712391948|35.232478750868765|00035000680488|ORAL HYGIENE|HBC|-80.8438|80.843800034139889|174|1
35.23102|98cc76716e1d4f670ad9a5849bff4fa4e904695a|4.29|2014-11-28 20:33:00|80.843945456961976|2|2840016014|205|35.233522162802032|0|59|201|-80.70901|31|35.17335|POTATO CHIPS|0.29|1|LAYS DUAF CHEESY GARLIC BREAD|e829a323ff38f07bbea130697026b25eeedc25a3|0.17289340712391948|35.232478750868765|00028400150101|SNACKS|G1 GROCERY|-80.8438|80.843800034139889|174|1
35.23102|35b5cee3c1934989fd3d20c4f1d6253fd61063c1|3.55|2015-01-10 19:32:00|80.843945456961976|2|3800039125|205|35.233522162802032|0|59|81|-80.70901|9|35.17335|RTE CEREAL KIDS|0.0|1|KELLOGG FROOT LOOPS 8.7|e829a323ff38f07bbea130697026b25eeedc25a3|0.17289340712391948|35.232478750868765|00038000391255|CEREAL|G1 GROCERY|-80.8438|80.843800034139889|174|1
35.23102|35d3de2d4a5b7ed2bce778cc83b72958f7bd8772|4.39|2014-10-22 17:49:00|80.843945456961976|2|3800057074|205|35.233522162802032|0|59|81|-80.70901|9|35.17335|RTE CEREAL KIDS|0.0|1|KELLOGG KRAVE CHOCOLATE|e829a323ff38f07bbea130697026b25eeedc25a3|0.17289340712391948|35.232478750868765|00038000570742|CEREAL|G1 GROCERY|-80.8438|80.843800034139889|174|1
35.23102|633a635d2ccd2302af892b772b9c35380f233db7|2.29|2014-11-16 18:07:00|80.843945456961976|2|7203695175|205|35.233522162802032|0|59|1607|-80.70901|371|35.17335|FROZEN DOUGH (BREAD)|1.3|14|FRESH LRG FRENCH BREAD|e829a323ff38f07bbea130697026b25eeedc25a3|0.17289340712391948|35.232478750868765|00072036951755|BREAD|BAKERY|-80.8438|80.843800034139889|174|1
35.23102|d4c68442cc640c144541d4255395dea88aa29dc0|1.99|2014-12-02 19:33:00|80.843945456961976|2|7203688097|205|35.233522162802032|0|59|526|-80.70901|64|35.17335|FRESH MUSHROOMS|0.0|4|HT BUTTON MUSHROOMS|e829a323ff38f07bbea130697026b25eeedc25a3|0.17289340712391948|35.232478750868765|00072036880970|FRESH PRODUCE|PRODUCE|-80.8438|80.843800034139889|174|1
35.23102|31d3f8565535dc657671293d9a69f6f92a3aa987|5.99|2014-09-16 19:19:00|1.4094857484078087|2|7203663044|205|0.6148972978359727|0|26|974|-80.8438|201|35.23102|FRESH TURKEY|2.0|2|HT 93% LEAN GROUND TURKEY|e829a323ff38f07bbea130697026b25eeedc25a3|0.17289340712391948|0.61471665291522548|00072036630445|POULTRY|MEAT|-80.8438|1.4109904898237917|205|1
35.23102|0c25f1e028f1fb2df64d2d3e50611b92edfd238e|3.89|2014-11-13 16:48:00|80.843945456961976|2|7203663092|205|35.233522162802032|0|59|1263|-80.70901|57|35.17335|GOOD FOR YOU MILK|0.5|3|HARRIS TEETER FAT FREE LACTOSE|e829a323ff38f07bbea130697026b25eeedc25a3|0.17289340712391948|35.232478750868765|00072036630940|MILK|DAIRY|-80.8438|80.843800034139889|174|1
35.23102|42feb2b0a7662c002d079137854f4eff37ac86b4|1.29|2014-11-29 22:16:00|80.843945456961976|2|7203657030|205|35.233522162802032|0|59|322|-80.70901|53|35.17335|SOUR CREAM|0.0|3|HT LIGHT SOUR CREAM|e829a323ff38f07bbea130697026b25eeedc25a3|0.17289340712391948|35.232478750868765|00072036600349|CULTURES|DAIRY|-80.8438|80.843800034139889|174|1
35.23102|db7c89e4cba58bf73cafaee24707002c0d829cd4|0.5|2014-09-24 15:28:00|80.843945456961976|2|4178900211|205|35.233522162496101|0|59|1203|-80.709466|33|35.124987|RAMEN|0.12|1|MARUCHAN RAMEN CHICKEN|e829a323ff38f07bbea130697026b25eeedc25a3|0.17289340712391948|35.232478750868765|00041789002113|SOUP|G1 GROCERY|-80.8438|80.843801515180928|157|2
35.23102|ee3af061cefc4a69c827465ca9e5b35580ecf6ce|3.19|2014-10-29 12:23:00|80.843945456961976|2|4060034500|205|35.233522162802032|0|59|313|-80.70901|51|35.17335|MARGARINE|0.0|3|ICBINB SPREAD BOWL|e829a323ff38f07bbea130697026b25eeedc25a3|0.17289340712391948|35.232478750868765|00040600345002|BUTTER & MARGARINE|DAIRY|-80.8438|80.843800034139889|174|1
35.23102|a50fa4b052579fd99e2f86c0d44bbcab27d8b514|2.29|2014-12-31 21:08:00|80.843945456961976|2|3890000407|205|35.233522162802032|0|59|105|-80.70901|16|35.17335|FRUIT CUPS AND GELS|0.29|1|DOLE 4PK PEACH LS|e829a323ff38f07bbea130697026b25eeedc25a3|0.17289340712391948|35.232478750868765|00038900029708|FRUIT-CAN/JAR|G1 GROCERY|-80.8438|80.843800034139889|174|1
35.23102|cb41a55f0fbe68dfacc994c9222869943cf867cb|0.6|2014-09-16 14:35:00|1.4094857484078087|2|7047000641|205|0.6148972978359727|0|26|688|-80.8438|61|35.23102|LIGHT|0.0|3|YOPLAIT LIGHT BLUEBERRY|e829a323ff38f07bbea130697026b25eeedc25a3|0.17289340712391948|0.61471665291522548|00070470006529|YOGURT|DAIRY|-80.8438|1.4109904898237917|205|1
35.23102|3fa991ea3e94ab114f42aeef2f4ae92725dc5541|2.69|2015-01-19 12:27:00|80.843945456961976|2|7294570544|205|35.233522162802032|0|59|1025|-80.70901|162|35.17335|WHITE|0.4|7|SL S&S  W.G. WHITE BREAD|e829a323ff38f07bbea130697026b25eeedc25a3|0.17289340712391948|35.232478750868765|00072945705449|SLICED BREAD|COMMERCIAL BAKERY|-80.8438|80.843800034139889|174|1
35.23102|d57072c4764a900d0f324f570b79a2c49ea58fe1|4.65|2014-09-17 17:31:00|1.4094857484078087|2|3000006119|205|0.6148972978359727|0|26|74|-80.8438|9|35.23102|RTE CEREAL ALL FAMILY|2.15|1|QUAKER CINNAMON LIFE|e829a323ff38f07bbea130697026b25eeedc25a3|0.17289340712391948|0.61471665291522548|00030000060834|CEREAL|G1 GROCERY|-80.8438|1.4109904898237917|205|1
35.23102|326f81073996dfd19cfb7b1d9fc9ad41d9528be3|2.69|2014-11-27 13:36:00|80.843945456961976|2|70935100013|205|35.233522162802032|0|59|556|-80.70901|64|35.17335|PACKAGED VEGETABLES|0.19|4|APIO BROCCOLI & CAULIFLOWER|e829a323ff38f07bbea130697026b25eeedc25a3|0.17289340712391948|35.232478750868765|00709351000263|FRESH PRODUCE|PRODUCE|-80.8438|80.843800034139889|174|1
35.23102|a4c5ec123b65c34a81f41dadd24515f3c18330a6|4.57|2015-02-27 20:39:00|80.843945456961976|2|5000062264|205|35.233522162802032|0|59|326|-80.70901|54|35.17335|COOKIES/BROWNIES-REFRIGERATED|0.0|3|NESTLE CHOCOLATE CHIP TUB|e829a323ff38f07bbea130697026b25eeedc25a3|0.17289340712391948|35.232478750868765|00050000622641|DOUGH PRODUCTS|DAIRY|-80.8438|80.843800034139889|174|1
35.23102|c4f2939c635e28594b7392f5ecddae5792bf656a|6.0|2014-11-08 17:32:00|80.843945456961976|2||205|35.233522162802032|0|59|511|-80.70901|64|35.17335|FRESH AVOCADOS|0.75|4|AVOCADOS, HASS XL 36CT|e829a323ff38f07bbea130697026b25eeedc25a3|0.17289340712391948|35.232478750868765|00204770000004|FRESH PRODUCE|PRODUCE|-80.8438|80.843800034139889|174|3
35.23102|4c3cf78b05801e3f2daf667b60bcbdba3e7d9341|4.99|2014-10-22 22:24:00|80.843945456961976|2|3022100607|205|35.233522162802032|0|59|6249|-80.70901|1550|35.17335|SMALL HAND TOOLS|1.5|18|"MS FIX-IT 6"" ADJUSTABLE WRENCH"|e829a323ff38f07bbea130697026b25eeedc25a3|0.17289340712391948|35.232478750868765|00030221006079|HARDWARE|GM|-80.8438|80.843800034139889|174|1
35.341927|96c69c4ee3a6ec6a1952532bd6976db322db87cb|1.89|2014-12-26 16:15:00|1.4102725052409182|4|7033050604|220|0.6168329901494819|0|1|6586|-80.764523|1564|35.341927|CORRECTION SUPPLY|0.0|18|BIC WHT OUT PL QUK DRY (50604)|ea46c6964444e258858a5c34bc74182113b6a30d|1.009591131086844|0.61833652052202714|00070330506046|SCHOOL & OFFICE SUPPLY|GM|-80.764523|1.4096068451526882|220|1
35.341927|35be7711f1359d3096f9118004556002bb1ca328|2.29|2014-12-01 10:17:00|1.4102725052409182|4|7800023046|220|0.6168329901494819|0|1|54|-80.764523|8|35.341927|DIET|1.29|23|CANADA DRY DT CRNBRY GINGR ALE|ea46c6964444e258858a5c34bc74182113b6a30d|1.009591131086844|0.61833652052202714|00078000141467|CARBONATED BEVERAGES|BEVERAGE|-80.764523|1.4096068451526882|220|1
35.103409|b22d2982cb9b591f70b675b695b80614983b30a2|5.38|2015-03-05 15:17:00|80.992238315890603|0|79357321453|88|35.170216455913774|0|22|4778|-80.847383|1230|35.024464|BARS-PROTEIN|0.19|17|QUEST CHOCCHIP COOKIEDOUGH BAR|ebaac8b3b89528060acccebaa81997b075ad044d|4.6162339350461075|35.131650835559327|00793573214539|SPORTS NUTRITIONAL|HBC|-80.992182|80.992195776110293|317|2
35.103409|09c11422042cec0f0dcbeb30a909db24711dbb7b|5.38|2015-03-01 19:57:00|1.4132775322775095|0|79357321453|88|0.6126700657242101|0|58|4778|-80.992182|1230|35.103409|BARS-PROTEIN|0.19|17|QUEST COOKIES & CREAM BAR|ebaac8b3b89528060acccebaa81997b075ad044d|4.6162339350461075|0.61177642288969325|00793573238467|SPORTS NUTRITIONAL|HBC|-80.992182|1.413580244274486|88|2
35.372142|d250873e349d8202ae33643e2e040ac4aad65fc5|8.99|2015-02-01 16:18:00|1.4102725052409182|2|7203695312|122|0.617360341382972|0|1|1970|-80.782849|475|35.372142|COLD PRE-MADE|3.0|6|SUPREME PIZZA|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00072036953124|PIZZA|DELI|-80.782849|1.4099266941914086|122|1
35.372142|b1f4d6a388d30bb3c0be3e2105bdde44a1a28f4c|3.29|2015-02-13 21:03:00|1.4102725052409182|2|3000005040|122|0.617360341382972|0|1|12|-80.782849|2|35.372142|PANCAKE MIXES|0.0|1|AJEMIMA PANCAKE MIX|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00030000050408|BAKING MIXES|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|613297d3ad83f17741f79b128782a451224c45ce|9.99|2015-02-07 21:15:00|1.4102725052409182|2|3700086527|122|0.617360341382972|0|1|427|-80.782849|72|35.372142|NFS-TOILET TISSUE|2.0|1|CHARMIN BATH SENSITIVE 6MR|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00037000857365|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|543f7d3a61a3c542f0f5f5ec21d19e4c12f903bf|9.99|2015-02-23 13:00:00|1.4102725052409182|2|3700086527|122|0.617360341382972|0|1|427|-80.782849|72|35.372142|NFS-TOILET TISSUE|0.0|1|CHARMIN BATH SENSITIVE 6MR|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00037000857365|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|f7934c9c13e556dc61d8dab212a872d1ca43ad08|9.69|2014-11-20 17:36:00|80.779636304526477|2|3700086527|122|35.397000260101713|0|17|427|-80.764523|72|35.341927|NFS-TOILET TISSUE|0.0|1|CHARMIN BATH SENSITIVE 6MR|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|35.392509581117899|00037000857365|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.782849|80.78285603145379|220|1
35.372142|f8458e8c6ccff351d139d406a79da579c308c6ac|1.29|2014-11-19 16:30:00|1.4102725052409182|2|2700039014|122|0.617360341382972|0|1|257|-80.782849|39|35.372142|TOMATOES|0.0|1|HUNTS TOMATO SAUCE 15|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00027000390146|VEGETABLES-CAN/JAR|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|a5b86b18de15d6236957110622118957c7592128|7.99|2015-01-08 18:37:00|1.4102725052409182|2|2840000288|122|0.617360341382972|0|1|205|-80.782849|31|35.372142|REMAINING SNACKS|2.0|1|FRITOLAY FLAVOR 20 CTN|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00028400002899|SNACKS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|2b6bf667386885b2098980368ba56f4da8da1d81|7.49|2014-12-03 17:39:00|1.4102725052409182|2|2840000288|122|0.617360341382972|0|1|205|-80.782849|31|35.372142|REMAINING SNACKS|0.5|1|FRITOLAY FLAVOR 20 CTN|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00028400002899|SNACKS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|8afc77aefc648e1185ab5745813274d980f59d8d|4.99|2014-11-09 17:45:00|1.4102725052409182|2|7495618054|122|0.617360341382972|0|1|492|-80.782849|101|35.372142|KOSHER WIENERS|0.49|19|HEBREW NATIONAL BUN BEEF FRANK|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00074956284005|WIENERS|CASE READY MEATS|-80.782849|1.4099266941914086|122|1
35.372142|44c9ac237c46b13c0d8c6aecca66a67dbffcd4b1|11.38|2015-02-08 14:55:00|1.4102725052409182|2|7495618054|122|0.617360341382972|0|1|492|-80.782849|101|35.372142|KOSHER WIENERS|2.84|19|HEBREW NATIONAL BUN BEEF FRANK|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00074956284005|WIENERS|CASE READY MEATS|-80.782849|1.4099266941914086|122|2
35.372142|d4e4dccb06800c38b6bd93fc231cf28aba82f7a5|5.49|2014-12-28 15:19:00|1.4102725052409182|2|7495618054|122|0.617360341382972|0|1|492|-80.782849|101|35.372142|KOSHER WIENERS|0.99|19|HEBREW NATIONAL BUN BEEF FRANK|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00074956284005|WIENERS|CASE READY MEATS|-80.782849|1.4099266941914086|122|1
35.372142|7ef7ba2589a90f1c5c81bff9e78d1616ad19b29c|1.49|2014-11-11 17:43:00|1.4102725052409182|2||122|0.617360341382972|0|1|525|-80.782849|64|35.372142|FRESH LETTUCE|0.0|4|ICEBERG LETTUCE|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00204061000003|FRESH PRODUCE|PRODUCE|-80.782849|1.4099266941914086|122|1
35.372142|2a4de187209c3b60cf0d1b317806eeea675137c3|3.1|2015-01-28 13:56:00|1.4102725052409182|2|8000051306|122|0.617360341382972|0|1|189|-80.782849|29|35.372142|TUNA-POUCH|1.1|1|STARKIST CREATION LEMON PEPPER|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00080000513090|SEAFOOD-CANNED|G1 GROCERY|-80.782849|1.4099266941914086|122|2
35.372142|edfecdabb3df7789970540a88e96930be8ad226f|9.98|2015-02-17 11:01:00|1.4102725052409182|2|7203658011|122|0.617360341382972|0|1|484|-80.782849|101|35.372142|BEEF WIENERS|2.5|19|HT BUNSIZE BEEF FRANKS|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00072036580115|WIENERS|CASE READY MEATS|-80.782849|1.4099266941914086|122|2
35.372142|0febbafd54d7692cb1140b19e1fdbef428d334c0|9.98|2014-09-27 15:38:00|1.4102725052409182|2|7203658011|122|0.617360341382972|0|1|484|-80.782849|101|35.372142|BEEF WIENERS|0.0|19|HT BUNSIZE BEEF FRANKS|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00072036580115|WIENERS|CASE READY MEATS|-80.782849|1.4099266941914086|122|2
35.372142|11399e8bc2aa14c07ba592539dffe651741c4b5d|3.69|2014-10-12 16:12:00|1.4102725052409182|2|7203678062|122|0.617360341382972|0|1|238|-80.782849|38|35.372142|RICE FLAVORED|0.0|1|HT TRADER RISOTTO GAR HERB|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00072036780645|RICE GRAINS AND BEANS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|7dc92399aa213fd2c177f70b1ec8256c274c7d85|7.38|2015-01-17 18:24:00|1.4102725052409182|2|7203678062|122|0.617360341382972|0|1|238|-80.782849|38|35.372142|RICE FLAVORED|2.38|1|HT TRADER RISOTTO GAR HERB|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00072036780645|RICE GRAINS AND BEANS|G1 GROCERY|-80.782849|1.4099266941914086|122|2
35.372142|f6942cc0537e543510ef781cec5d44b5f430ba00|1.79|2014-12-09 14:02:00|1.4102725052409182|2|20406100000|122|0.617360341382972|0|1|525|-80.782849|64|35.372142|FRESH LETTUCE|0.0|4|ICEBERG LETTUCE|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00033383650203|FRESH PRODUCE|PRODUCE|-80.782849|1.4099266941914086|122|1
35.372142|9d8479ab03dab80822438e0978bed2750c1ab664|3.29|2015-01-10 15:54:00|1.4102725052409182|2|2840011895|122|0.617360341382972|0|1|204|-80.782849|31|35.372142|TORTILLA CHIPS|0.0|1|TOSTITOS CANTINA TRADITIONAL|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00028400118958|SNACKS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|ea258996318fc3985c495d52eb7c99e723269d8b|3.29|2015-03-02 18:14:00|1.4102725052409182|2|2840011895|122|0.617360341382972|0|1|204|-80.782849|31|35.372142|TORTILLA CHIPS|0.79|1|TOSTITOS CANTINA TRADITIONAL|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00028400118958|SNACKS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|37f328b96d626f6afcb944a342241f8d2a728b75|3.49|2015-02-16 15:18:00|1.4102725052409182|2|2700049016|122|0.617360341382972|0|1|200|-80.782849|31|35.372142|MICROWAVE POPCORN|0.0|1|OR REDENBUDER MOVIE 3 CT BOWL|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00027000490167|SNACKS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|783d0129847ee0a90b89ddbbca7c52005647d5a2|13.12|2015-03-07 17:44:00|1.4102725052409182|2|20332600000|122|0.617360341382972|0|1|641|-80.782849|137|35.372142|PREMIUM PORK|1.89|2|VALUE PK BONE-IN PORK CHOPS|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00203326000000|PORK|MEAT|-80.782849|1.4099266941914086|122|1
35.372142|76de5bb6ffc2d7f67703fe17225eb4c1766b06c1|1.99|2015-02-22 13:51:00|80.779636304526477|2|7680828073|122|35.397000260101713|0|17|149|-80.764523|23|35.341927|WHSE PASTA CORE|0.49|1|BARILLA PASTA ELBOWS|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|35.392509581117899|00076808516135|PASTA|G1 GROCERY|-80.782849|80.78285603145379|220|1
35.372142|c5887619a7d9199f44900f5218afed9fb2448f57|15.42|2015-02-24 17:31:00|80.779636304526477|2|20332600000|122|35.397000260101713|0|17|641|-80.764523|137|35.341927|PREMIUM PORK|2.23|2|VALUE PK BONE-IN PORK CHOPS|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|35.392509581117899|00203326000000|PORK|MEAT|-80.782849|80.78285603145379|220|1
35.372142|34942fb36f092234a53b28bb8ee435e6176e8212|1.49|2015-01-11 09:08:00|1.4102725052409182|2|7053801184|122|0.617360341382972|0|1|50|-80.782849|7|35.372142|PEG CANDY|0.0|1|BOB'S SWEET STRIPE MINT|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00070538011847|CANDY|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|7694986c36317702e156d824c1d9ef703edf1959|4.3|2014-11-23 15:30:00|1.4102725052409182|2|7092047449|122|0.617360341382972|0|1|1147|-80.782849|229|35.372142|HOT COCOA MIX|0.65|1|SWISS MISS MARSHMALLOW 10 CT|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00070920474502|COCOAS CREAMERS SYRUPS|G1 GROCERY|-80.782849|1.4099266941914086|122|2
35.372142|bb21100bfaf318c95dd5e538e8bb6b5dba3f837a|3.99|2014-10-04 18:11:00|1.4102725052409182|2|5210000647|122|0.617360341382972|0|1|1245|-80.782849|34|35.372142|SINGLE SPICES|0.0|1|MC ONION POWDER|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00052100006475|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|f834730d88109b0d0c9f66a0cef53a442907b939|1.95|2014-09-26 15:04:00|1.4102725052409182|2|4300000953|122|0.617360341382972|0|1|272|-80.782849|307|35.372142|TOPPINGS FROZEN|0.0|5|COOL WHIP WHIPPED TOPPING|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00043000009536|DESSERTS FROZEN|FROZEN|-80.782849|1.4099266941914086|122|1
35.372142|0d268024b1522ede27183a936da5885a733a1dc3|8.78|2014-12-22 20:27:00|1.4102725052409182|2|4133310310|122|0.617360341382972|0|1|8460|-80.782849|1769|35.372142|BATTERY-ELECTRONICS|0.0|18|DURACELL MED 2032 1PK|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00041333103105|BATTERY & FLASHLIGHT|GM|-80.782849|1.4099266941914086|122|2
35.372142|76d3ab30a34e801c34c8ed150748fc3fe29d4b54|16.41|2014-09-28 14:02:00|1.4102725052409182|2|20188000000|122|0.617360341382972|0|1|299|-80.782849|49|35.372142|ANGUS BEEF|0.0|2|ANGUS BEEF BNLS CHUCK ROAST|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00201880000009|BEEF|MEAT|-80.782849|1.4099266941914086|122|1
35.372142|08345a1142650a1b25b5e7e3684473eb090c7940|7.49|2014-12-26 21:09:00|1.4102725052409182|2|31031032503|122|0.617360341382972|0|1|4026|-80.782849|1080|35.372142|ORAL HYGI ORAL MEDICATN|0.0|17|ORAJEL SEVERE TOOTHACHE GEL|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00310310325039|ORAL HYGIENE|HBC|-80.782849|1.4099266941914086|122|1
35.372142|1455dcb6bdb852bae3637240a1f4f98280ee68e1|39.92|2014-09-20 10:56:00|80.779636304526477|2|4124400006|122|35.397000260101713|0|17|128|-80.764523|20|35.341927|APPLE JUICE-SHELF|0.0|1|MARTINELLI SPARKLING CIDER|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|35.392509581117899|00041244000067|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.782849|80.78285603145379|220|8
35.372142|1e0e70cc1d6f8798f7393ecb91eb61017e3a625b|1.39|2014-10-22 16:44:00|1.4102725052409182|2|4100002253|122|0.617360341382972|0|1|1439|-80.782849|274|35.372142|DRY DINNERS|0.39|1|KNORR PASTA BUTTER HERB|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00041000022517|PREP FOODS DINNERS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|0f8d249f83e79cb1ababd61d8df33f522dd46229|1.79|2015-01-22 17:33:00|1.4102725052409182|2|3940001614|122|0.617360341382972|0|1|243|-80.782849|39|35.372142|BAKED BEANS|0.0|1|BUSH BKD BEAN W/ONION 28|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00039400016038|VEGETABLES-CAN/JAR|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|23ae661ace06d856156ab0cd0b7cb3d76e4c647a|7.98|2014-09-10 09:39:00|1.4102725052409182|2|3800059644|122|0.617360341382972|0|1|81|-80.782849|9|35.372142|RTE CEREAL KIDS|2.0|1|KELLOGG FROSTED FLAKES 10.5|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00038000596445|CEREAL|G1 GROCERY|-80.782849|1.4099266941914086|122|2
35.372142|ce323e286eab046c624712e69e589c5f430793db|3.65|2015-02-18 10:49:00|80.779636304526477|2|3800059644|122|35.397000260101713|0|17|81|-80.764523|9|35.341927|RTE CEREAL KIDS|1.15|1|KELLOGG FROSTED FLAKES 10.5|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|35.392509581117899|00038000596445|CEREAL|G1 GROCERY|-80.782849|80.78285603145379|220|1
35.372142|d80ebc80183c8a889733d24b2627a66b1b7c0086|2.69|2015-01-19 18:09:00|1.4102725052409182|2|3663202720|122|0.617360341382972|0|1|688|-80.782849|61|35.372142|LIGHT|0.0|3|DANNON L&F STRAWBERRY|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00036632027207|YOGURT|DAIRY|-80.782849|1.4099266941914086|122|1
35.372142|767b178b8bfb2e305ac9a5caed3778f8edd383da|1.79|2015-01-11 17:17:00|1.4102725052409182|2|4150001310|122|0.617360341382972|0|1|76|-80.782849|11|35.372142|MEAT SAUCES|0.0|1|FRENCHS WORCESTERSHIRE 10|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00041500013107|CONDIMENTS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|3b4b417bc51650be24286b8c15af0a6828f617c0|1.81|2014-10-08 21:24:00|80.779636304526477|2||122|35.397000260101713|0|17|502|-80.764523|64|35.341927|FRESH BANANAS|0.0|4|BANANAS, YELLOW|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|35.392509581117899|00204011000008|FRESH PRODUCE|PRODUCE|-80.782849|80.78285603145379|220|1
35.372142|5ce6a0829cc193f6efafa8d1633f0bfc1265123c|1.96|2014-10-06 09:52:00|1.4102725052409182|2||122|0.617360341382972|0|1|502|-80.782849|64|35.372142|FRESH BANANAS|0.0|4|BANANAS, YELLOW|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.782849|1.4099266941914086|122|1
35.372142|ea7923b11482aec14cb40f5df57ba99caa3d402e|1.53|2014-11-23 06:16:00|1.4102725052409182|2||122|0.617360341382972|0|1|502|-80.782849|64|35.372142|FRESH BANANAS|0.0|4|BANANAS, YELLOW|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.782849|1.4099266941914086|122|1
35.372142|3b0190b432ded552d62d0ea4a1e7b3846520c4a3|2.59|2014-11-18 17:38:00|1.4102725052409182|2|7203663996|122|0.617360341382972|0|1|342|-80.782849|57|35.372142|FRESH MILK|0.0|3|HARRIS TEETER 2%   MILK|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00072036639998|MILK|DAIRY|-80.782849|1.4099266941914086|122|1
35.372142|416e5bf972ec334164be9994ac324895b4523916|7.49|2014-12-28 18:46:00|1.4102725052409182|2|35497330981|122|0.617360341382972|0|1|4204|-80.782849|1200|35.372142|COUGH & COLD SYRUPS-CHILD|0.0|17|HYLANDS NT COLD N COUGH 4 KIDS|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00354973309814|COUGH/COLD/SINUS|HBC|-80.782849|1.4099266941914086|122|1
35.372142|f4eebf1bb62be483d517076dbef791d62050b7cc|15.1|2014-09-14 15:26:00|1.4102725052409182|2|20819400000|122|0.617360341382972|0|1|660|-80.782849|154|35.372142|FISH FILLETS WILD CGHT|5.04|12|WC FROZ TILAPIA FILLETS (PA)|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00208194000008|FISH FILLETS/STEAKS|SEAFOOD|-80.782849|1.4099266941914086|122|1
35.372142|7b49194aad86177516d1f6d6bb49b409630293bb|6.68|2014-12-18 16:57:00|1.4102725052409182|2|20889500000|122|0.617360341382972|0|1|648|-80.782849|154|35.372142|FISH FLTS/STK FARM RAISD|0.0|12|FR TILAPIA FILLET|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00208895000000|FISH FILLETS/STEAKS|SEAFOOD|-80.782849|1.4099266941914086|122|1
35.372142|7ffd015397a9f024b03ba183d5148823b2563306|20.21|2014-09-30 18:35:00|1.4102725052409182|2|20889500000|122|0.617360341382972|0|1|648|-80.782849|154|35.372142|FISH FLTS/STK FARM RAISD|7.59|12|FR TILAPIA FILLET|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00208895000000|FISH FILLETS/STEAKS|SEAFOOD|-80.782849|1.4099266941914086|122|1
35.372142|c57a91ae86339f42ca52953fdac7b5bd436994f3|50.120000000000005|2015-03-08 18:05:00|1.4102725052409182|2|20140400000|122|0.617360341382972|0|1|296|-80.782849|49|35.372142|RANCHER BEEF|20.9|2|BEEF LOIN NY STRIP STEAK BNLS|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00201404000003|BEEF|MEAT|-80.782849|1.4099266941914086|122|3
35.372142|af518c1f2bfb9c2f808d9698b3eba93403fca589|8.99|2014-12-07 19:07:00|1.4102725052409182|2|38137003600|122|0.617360341382972|0|1|3202|-80.782849|1015|35.372142|HAND & BODY THERAPEUTIC|1.5|17|AVEENO MOIST LOTION STRESS RLF|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00381370039167|HAND & BODY LOTION/SUN CARE|HBC|-80.782849|1.4099266941914086|122|1
35.372142|8127044bee8504a51b60ab712556bc9f8752fa1e|4.29|2014-10-23 16:06:00|1.4102725052409182|2|2840006399|122|0.617360341382972|0|1|204|-80.782849|31|35.372142|TORTILLA CHIPS|0.29|1|TOSTITOS HINT OF LIME|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00028400064040|SNACKS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|c7d64fa0a700027f50d6fc540dfcffe4484375b5|1.49|2015-01-02 17:59:00|1.4102725052409182|2|2840002819|122|0.617360341382972|0|1|206|-80.782849|31|35.372142|FRONT END SNACKS|0.0|1|LAYS CLASSIC|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00028400027960|SNACKS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|d5c74c94deeedab9b47d2e8d83119319026806b5|2.89|2015-03-05 19:25:00|1.4102725052409182|2|2100065894|122|0.617360341382972|0|1|1441|-80.782849|274|35.372142|MAC AND CHEESE|0.0|1|KRAFT DIN MAC CHS FAMILY|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00021000658947|PREP FOODS DINNERS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|d77c2e3932705b0eb4c95d98b86148e109b3407c|1.59|2014-10-02 17:26:00|1.4102725052409182|2|2200000512|122|0.617360341382972|0|1|48|-80.782849|7|35.372142|REGISTER GUM|0.0|1|(FE) 5 RAIN GUM 15PC|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00022000005144|CANDY|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|eef0b255a768716a0221f6865a4a1fd48ea67daf|8.69|2015-01-30 17:59:00|1.4102725052409182|2|20896400000|122|0.617360341382972|0|1|977|-80.782849|201|35.372142|FRESH HT CHICKEN|0.85|2|HT VALUE PK WING PORTIONS|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00208964000009|POULTRY|MEAT|-80.782849|1.4099266941914086|122|1
35.372142|7301c64394b72387079338249406b132ce18fca0|8.59|2014-11-08 07:39:00|1.4102725052409182|2|76211120604|122|0.617360341382972|0|1|35|-80.782849|10|35.372142|PREMIUM WHOLE BEAN|1.6|1|STARBUCKS BLONDE VERONA WH/BN|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00762111949806|COFFEE|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|4af4dcb63198775d44601dc25602b326da3ab79d|7.65|2015-01-03 08:23:00|1.4102725052409182|2|76211120604|122|0.617360341382972|0|1|35|-80.782849|10|35.372142|PREMIUM WHOLE BEAN|0.0|1|STARBUCKS BLONDE VERONA WH/BN|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00762111949806|COFFEE|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|c15796367e036d4aea3a9a909bd5f1e1a99bc19a|4.99|2014-11-28 20:18:00|1.4102725052409182|2|3917445141|122|0.617360341382972|0|1|7221|-80.782849|1600|35.372142|WINTER GLOVES|1.0|18|I/O LADIES CHENILIE GLOVE|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00039174451417|SEASONAL MERCHANDISE|GM|-80.782849|1.4099266941914086|122|1
35.372142|643bc8dd253726e30e23f03e3bc2e55075f9995b|4.59|2014-12-29 10:19:00|1.4102725052409182|2|3800066330|122|0.617360341382972|0|1|61|-80.782849|9|35.372142|RTE CEREAL ADULT|2.59|1|KELLOGG SMART START CEREAL|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00038000663307|CEREAL|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|f461defeb7fbb83b953b1a68f4d59838916e56af|3.19|2014-11-01 08:04:00|1.4102725052409182|2|3760019991|122|0.617360341382972|0|1|175|-80.782849|27|35.372142|CANNED MEATS|0.0|1|HORMEL MAR KTC ROAST BEEF HASH|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00037600199919|PREPARED FOODS-RTS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|7f187cdbe9897765c31e9a99d73d32e13b6b29f6|7.99|2015-02-15 13:19:00|1.4102725052409182|2|2840000288|122|0.617360341382972|0|1|205|-80.782849|31|35.372142|REMAINING SNACKS|2.0|1|FRITOLAY CLASSIC 20 CTN|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00028400002882|SNACKS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|246dd7b942bb19b0fc358564535c04ad437f8fde|1.59|2014-12-28 15:05:00|80.779636304526477|2|1600043054|122|35.397000260101713|0|17|10|-80.764523|2|35.341927|LAYER CAKE MIX|0.0|1|BC SUPER MOIST RED VELVET MIX|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|35.392509581117899|00016000428997|BAKING MIXES|G1 GROCERY|-80.782849|80.78285603145379|220|1
35.372142|454da762341e6d080424c21b7ec5aa14eee83548|7.75|2014-12-11 17:12:00|1.4102725052409182|2|1258760034|122|0.617360341382972|0|1|443|-80.782849|76|35.372142|NFS-GARBAGE BAGS|0.4|1|GLAD TALL KTCHN DRAWSTG 13GL|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00012587786284|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|2698eefaa5b9b9dd484eb9261bbb1279797303c0|4.85|2014-11-06 10:02:00|80.779636304526477|2|1600048366|122|35.397000260101713|0|17|74|-80.764523|9|35.341927|RTE CEREAL ALL FAMILY|0.0|1|GM CHEERIOS HONEY NUT 21.6|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|35.392509581117899|00016000483668|CEREAL|G1 GROCERY|-80.782849|80.78285603145379|220|1
35.372142|d3d5193940a5a361280bf4b6d4120d3c4b49b031|3.55|2015-03-07 13:02:00|1.4102725052409182|2|3800039125|122|0.617360341382972|0|1|74|-80.782849|9|35.372142|RTE CEREAL ALL FAMILY|0.0|1|KELLOGG RICE KRISPIES 9|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00038000318443|CEREAL|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|17c2539d1811955eef583cefba68bdaa133705d8|9.99|2015-02-13 22:13:00|1.4102725052409182|2|84560401638|122|0.617360341382972|0|1|6984|-80.782849|1600|35.372142|VALENTINE NOVELTY-IMPORT|2.0|18|I/O VAL SPARKLE CHLLER 20OZ|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00845604016381|SEASONAL MERCHANDISE|GM|-80.782849|1.4099266941914086|122|1
35.372142|0ce5e1296d5e5d4f118f70c601bda00e6b2efd25|14.99|2014-09-10 15:38:00|1.4102725052409182|2|8066095615|122|0.617360341382972|0|1|459|-80.782849|83|35.372142|IMPORT BEER|0.0|16|CORONA EXTRA 12PK 12OZ BTL|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00080660956152|IMPORT BEER|BEER|-80.782849|1.4099266941914086|122|1
35.372142|786833f54179238a8a8caba17a5351c7a12d9d7a|1.29|2015-01-13 19:06:00|1.4102725052409182|2|980000761|122|0.617360341382972|0|1|48|-80.782849|7|35.372142|REGISTER GUM|0.0|1|TIC TAC ORANGE BIG PACK|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00009800007639|CANDY|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|b7b12853e9481f5b59a248896ba81c95ecc64873|1.29|2015-01-18 11:01:00|1.4102725052409182|2|980000761|122|0.617360341382972|0|1|48|-80.782849|7|35.372142|REGISTER GUM|0.0|1|TIC TAC ORANGE BIG PACK|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00009800007639|CANDY|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|dc28c7c9d88a16ca8043b7662a0d29b022acaa73|1.29|2015-01-10 15:20:00|1.4102725052409182|2|980000761|122|0.617360341382972|0|1|48|-80.782849|7|35.372142|REGISTER GUM|0.0|1|TIC TAC ORANGE BIG PACK|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00009800007639|CANDY|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|687c91e808bda77c17ca8dfa3c5a1f85a46ce3bd|1.29|2015-01-16 19:26:00|1.4102725052409182|2|980000761|122|0.617360341382972|0|1|48|-80.782849|7|35.372142|REGISTER GUM|0.0|1|TIC TAC ORANGE BIG PACK|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00009800007639|CANDY|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|f5a4f189d11c2c971c094857eb85fc20d042a914|1.79|2014-12-21 07:15:00|1.4102725052409182|2|5100001047|122|0.617360341382972|0|1|212|-80.782849|33|35.372142|CONDENSED SOUP|0.12|1|CAMP COND CREAM OF ONION|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00051000016171|SOUP|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|4b3ab919f442ce60d10ef857b299c5395d6e59e2|4.99|2014-10-08 21:20:00|80.779636304526477|2|6827493471|122|35.397000260101713|0|17|31|-80.764523|4|35.341927|NON CARBONATED WATER|1.2|1|NESTLE PURE LIFE .5L 24PK|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|35.392509581117899|00068274934711|BOTTLED WATER|G1 GROCERY|-80.782849|80.78285603145379|220|1
35.372142|8a8b6a27814f04aba63f68a897e4f74df391489e|4.99|2014-11-03 22:03:00|1.4102725052409182|2|6827493471|122|0.617360341382972|0|1|31|-80.782849|4|35.372142|NON CARBONATED WATER|1.2|1|NESTLE PURE LIFE .5L 24PK|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00068274934711|BOTTLED WATER|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|565b54b4348456284c00fb7383f6e8fcc1e6a237|2.35|2014-10-08 17:57:00|1.4102725052409182|2|2400003409|122|0.617360341382972|0|1|105|-80.782849|16|35.372142|FRUIT CUPS AND GELS|0.0|1|DEL MONTE 4PK NSA PEACH|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00024000393429|FRUIT-CAN/JAR|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|38fe2cf80beb16907cee04f5126df806b03c62ba|4.95|2015-01-10 17:27:00|1.4102725052409182|2|3450015136|122|0.617360341382972|0|1|312|-80.782849|51|35.372142|BUTTER|0.0|3|L O L BUTTER QUARTERS|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00034500151368|BUTTER & MARGARINE|DAIRY|-80.782849|1.4099266941914086|122|1
35.372142|e15c212ad9b26d23d6aeae3ff4356ff09eb22e5f|6.49|2015-03-02 22:04:00|1.4102725052409182|2|7756719329|122|0.617360341382972|0|1|273|-80.782849|43|35.372142|PREMIUM NOVELTIES|0.0|5|MAGNUM MINI ALMOND IC BAR 6PK|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00077567193407|FROZEN NOVELTIES|FROZEN|-80.782849|1.4099266941914086|122|1
35.372142|9c537fbee53955c2f20291fdbdf78770ae92c730|1.89|2014-10-18 17:13:00|1.4102725052409182|2|7203663202|122|0.617360341382972|0|1|1262|-80.782849|57|35.372142|HALF N HALF WHIPPING CREAM|0.0|3|HT WHIPPING CREAM|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00072036632029|MILK|DAIRY|-80.782849|1.4099266941914086|122|1
35.372142|da47fe4da4d601ce53854a2b93f7b32c515f34b5|3.49|2014-10-22 09:42:00|80.779636304526477|2|3800001611|122|35.397000260101713|0|17|61|-80.764523|9|35.341927|RTE CEREAL ADULT|0.0|1|KELLOGG SPECIAL K RED BERRIES|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|35.392509581117899|00038000599231|CEREAL|G1 GROCERY|-80.782849|80.78285603145379|220|1
35.372142|44635f276e49af005d1d3235c1defe17dfc483a0|2.85|2015-01-07 10:12:00|80.779636304526477|2|4400000055|122|35.397000260101713|0|17|88|-80.764523|13|35.341927|FLAKED SODA CRACKERS|0.85|1|NABISCO PREMIUMS|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|35.392509581117899|00044000000578|CRACKERS|G1 GROCERY|-80.782849|80.78285603145379|220|1
35.372142|0cca16bc1e8ec8c12485bf0584ca8aab4399b3b7|1.79|2015-01-01 19:07:00|1.4102725052409182|2|8079380770|122|0.617360341382972|0|1|99|-80.782849|32|35.372142|LIQUID TEA|0.0|1|D FUZE SLENDER TROPICAL PUNCH|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00080793807765|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|d878f6d2fb7b4502bd5b314cc12100fcfe2992bb|1.79|2014-11-01 18:23:00|1.4102725052409182|2|8079380770|122|0.617360341382972|0|1|99|-80.782849|32|35.372142|LIQUID TEA|0.12|1|D FUZE SLENDER TROPICAL PUNCH|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00080793807765|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|2f6bfe1d368c30b045bb5a78ad14e2154f31ceec|1.39|2015-02-11 17:34:00|1.4102725052409182|2|1254667609|122|0.617360341382972|0|1|48|-80.782849|7|35.372142|REGISTER GUM|0.0|1|TRIDENT WHITE PEPPERMINT|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00012546676090|CANDY|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|e6fc63a4e94804733c0a6a0e7a23ca878fa6bb4c|14.99|2015-02-12 15:39:00|1.4102725052409182|2|75444108251|122|0.617360341382972|0|1|663|-80.782849|154|35.372142|FISH FILLETS/STEAKS PKGD|5.02|12|TILAPIA FILLETS|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00664183000617|FISH FILLETS/STEAKS|SEAFOOD|-80.782849|1.4099266941914086|122|1
35.372142|ad2e0506e72ee42409d20bf971ce9028934d82f7|9.31|2014-11-26 16:55:00|1.4102725052409182|2|20896100000|122|0.617360341382972|0|1|977|-80.782849|201|35.372142|FRESH HT CHICKEN|2.9|2|HT VALUE PK CHICKEN DRUMSTICKS|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00208961000002|POULTRY|MEAT|-80.782849|1.4099266941914086|122|1
35.372142|46b4e50973f347d60c66793675ae0639be44c259|1.29|2015-03-07 14:38:00|1.4102725052409182|2|4000000051|122|0.617360341382972|0|1|47|-80.782849|7|35.372142|REGISTER BARS|0.0|1|SKITTLES BITE SIZE|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00040000001607|CANDY|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|6a9196a6144d9eecc013cbc799aef187c334eb57|2.0|2015-02-24 16:52:00|80.779636304526477|2|2840019079|122|35.397000260101713|0|17|201|-80.764523|31|35.341927|POTATO CHIPS|0.0|1|CHESTERS HOT FRIES|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|35.392509581117899|00028400190787|SNACKS|G1 GROCERY|-80.782849|80.78285603145379|220|1
35.372142|25f99936d705ebf0a3e20c62d10ea6073eff3bcb|4.49|2015-03-03 18:41:00|1.4102725052409182|2|5200012125|122|0.617360341382972|0|1|171|-80.782849|20|35.372142|ISOTONIC DRINKS|0.71|1|GATORADE ASTAR ORANGE 6PK|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00052000129359|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|0d31f63d92b83051c4aea9d6cebebc6d466bba27|1.79|2015-01-31 12:59:00|1.4102725052409182|2|5100005977|122|0.617360341382972|0|1|212|-80.782849|33|35.372142|CONDENSED SOUP|0.0|1|CAMP HLTHY REQ CREAM OF CELERY|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00051000065698|SOUP|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|a484e6b50293570638f74ab78ec224158c3015b1|2.0|2014-12-31 19:06:00|1.4102725052409182|2|4300000953|122|0.617360341382972|0|1|272|-80.782849|307|35.372142|TOPPINGS FROZEN|1.01|5|COOL WHIP LITE WHIPPED TOPPING|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00043000009505|DESSERTS FROZEN|FROZEN|-80.782849|1.4099266941914086|122|1
35.372142|db2c2e46a4fbbcfc23234eb56c3f1f46fcd6c2bc|5.16|2014-10-09 15:45:00|1.4102725052409182|2|1657191030|122|0.617360341382972|0|1|30|-80.782849|4|35.372142|CARBONATED WATER|1.16|1|SPARKLING ICE KIWI STRAWBERRY|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00016571910327|BOTTLED WATER|G1 GROCERY|-80.782849|1.4099266941914086|122|4
35.372142|023b38ea17dfb22eb7c829c7eb8404c71c6149a8|1.29|2015-01-02 19:48:00|1.4102725052409182|2|2200000899|122|0.617360341382972|0|1|48|-80.782849|7|35.372142|REGISTER GUM|0.0|1|EXTRA SPEARMINT|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00022000008992|CANDY|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|8f9a266a6487a11f97a3d212e17a4d8f2cfaeea0|3.15|2015-01-06 08:02:00|1.4102725052409182|2|7225003706|122|0.617360341382972|0|1|1026|-80.782849|162|35.372142|WHEAT|0.0|7|NATOWN HONEYWHEAT BRD|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00072250037068|SLICED BREAD|COMMERCIAL BAKERY|-80.782849|1.4099266941914086|122|1
35.372142|1f426d4f52b8747995cf9208c5b232a02cb2e891|3.69|2015-02-27 10:01:00|80.779636304526477|2|2500005542|122|35.397000260101713|0|17|335|-80.764523|56|35.341927|ORANGE JUICE-REGRIGERATED|0.69|3|SIMPLY ORANGE CALCIUM|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|35.392509581117899|00025000055430|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.782849|80.78285603145379|220|1
35.372142|064a7c393c076345ee2255683b4046f51b036d76|2.39|2014-12-10 11:36:00|1.4102725052409182|2|31254662159|122|0.617360341382972|0|1|4207|-80.782849|1200|35.372142|COUGH DROP-ADULT|1.2|17|HALLS SF BREEZERS COOL BERRY|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00312546632233|COUGH/COLD/SINUS|HBC|-80.782849|1.4099266941914086|122|1
35.372142|8435e7e0a3d3b7eb425d56d8015716fd83badd6f|6.99|2015-01-24 20:15:00|1.4102725052409182|2|35058053404|122|0.617360341382972|0|1|4189|-80.782849|1200|35.372142|ALLERGY REMEDY-CHILDREN|0.0|17|BENADRYL CHILD ALLRGY CHRY LQ|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00350580534045|COUGH/COLD/SINUS|HBC|-80.782849|1.4099266941914086|122|1
35.372142|68b4de894fc4d7f0c97317ff2c280bfd20245372|15.99|2014-10-24 18:32:00|1.4102725052409182|2|18195400004|122|0.617360341382972|0|1|459|-80.782849|83|35.372142|IMPORT BEER|0.0|16|PERONI 12PK|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00181954000046|IMPORT BEER|BEER|-80.782849|1.4099266941914086|122|1
35.372142|ff222165c4e3969da6c85cba37f8221cf7a403ca|3.49|2014-10-13 22:02:00|80.779636304526477|2|2840023981|122|35.397000260101713|0|17|203|-80.764523|31|35.341927|CHEESE SNACKS|1.75|1|CHEETOS CRUNCHY HOT LIMON|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|35.392509581117899|00028400239851|SNACKS|G1 GROCERY|-80.782849|80.78285603145379|220|1
35.372142|18174de5a40ccc784173ec14d6a83bc37fdf977d|1.0|2014-11-30 21:48:00|1.4102725052409182|2|3400000031|122|0.617360341382972|0|1|47|-80.782849|7|35.372142|REGISTER BARS|0.25|1|HERSHEY KIT KAT BAR|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00034000002467|CANDY|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|6034fdabc488e134a54dfa68201ba91a745dc735|0.99|2014-10-06 19:52:00|1.4102725052409182|2|3400000031|122|0.617360341382972|0|1|47|-80.782849|7|35.372142|REGISTER BARS|0.5|1|HERSHEY ALMOND BAR|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00034000002412|CANDY|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|fd0f211ebef5c44d8e394f301e2c9a4cd00a00dc|1.0|2015-01-02 20:47:00|80.779636304526477|2|3400000031|122|35.397000260101713|0|17|47|-80.764523|7|35.341927|REGISTER BARS|0.0|1|HERSHEY ALMOND BAR|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|35.392509581117899|00034000002412|CANDY|G1 GROCERY|-80.782849|80.78285603145379|220|1
35.372142|3d0f0323d901ae2ddd1bf1c1a1df8191497dc8d0|4.29|2015-02-27 10:03:00|80.779636304526477|2|2100060085|122|35.397000260101713|0|17|316|-80.764523|52|35.341927|CREAM CHEESE|0.0|3|PHILLY SOFT CREAM CHEESE|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|35.392509581117899|00021000616886|CHEESE|DAIRY|-80.782849|80.78285603145379|220|1
35.372142|c358b7fa7e15bac5f50a4db3fb7e90cc43be960a|8.55|2014-11-29 18:15:00|80.779636304526477|2|3600038559|122|35.397000260101713|0|17|427|-80.764523|72|35.341927|NFS-TOILET TISSUE|0.0|1|COTTONELLE GENT CARE ALOE 12RL|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|35.392509581117899|00036000360943|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.782849|80.78285603145379|220|1
35.372142|20db8555f5ab8219b50f77f2ed074eef7d082187|4.58|2015-02-25 15:32:00|1.4102725052409182|2|7800023046|122|0.617360341382972|0|1|55|-80.782849|8|35.372142|REGULAR|0.79|23|CANADA DRY GINGER ALE NR 2LTR|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00078000152463|CARBONATED BEVERAGES|BEVERAGE|-80.782849|1.4099266941914086|122|2
35.372142|4cf673def4ff121bfebfac3d66daf7def052a895|8.99|2014-09-19 19:18:00|1.4102725052409182|2|87126011085|122|0.617360341382972|0|1|740|-80.782849|87|35.372142|NFS-ROSE BQT|0.0|9|BUNCH- 10 CONSUMER ROSE|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00871260110859|FLORAL|FLORAL|-80.782849|1.4099266941914086|122|1
35.372142|4f8792efbee30bfaf61e41f17aaa87b1ee55b074|1.19|2015-01-04 11:11:00|1.4102725052409182|2|7046209850|122|0.617360341382972|0|1|47|-80.782849|7|35.372142|REGISTER BARS|0.0|1|SOUR PATCH KIDS 2 OZ|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00070462098501|CANDY|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|775d3d762b8eab740c5c07d322108f9d2e0b0236|1.0|2015-01-18 14:50:00|80.779636304526477|2|3400000031|122|35.397000260101713|0|17|47|-80.764523|7|35.341927|REGISTER BARS|0.25|1|HERSHEY MILK CHOC BAR|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|35.392509581117899|00034000002405|CANDY|G1 GROCERY|-80.782849|80.78285603145379|220|1
35.372142|747807ca668f70366e30845c77ff7ee8e567d666|1.0|2015-02-06 22:20:00|1.4102725052409182|2|3400000031|122|0.617360341382972|0|1|47|-80.782849|7|35.372142|REGISTER BARS|0.0|1|HERSHEY MILK CHOC BAR|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00034000002405|CANDY|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|e213ff82a6cfd0b4c4e27ebe15998f3a7557d91b|0.99|2014-10-16 21:33:00|1.4102725052409182|2|3400000031|122|0.617360341382972|0|1|47|-80.782849|7|35.372142|REGISTER BARS|0.0|1|HERSHEY MILK CHOC BAR|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00034000002405|CANDY|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|9ff9317a10032c28c0cd602f9cfaa585fb00a57b|1.0|2014-10-23 20:05:00|1.4102725052409182|2|3400000031|122|0.617360341382972|0|1|47|-80.782849|7|35.372142|REGISTER BARS|0.0|1|HERSHEY MILK CHOC BAR|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00034000002405|CANDY|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|3e3bc6065be12713831a48a4a51ea3f48476fffe|1.0|2014-11-03 21:35:00|1.4102725052409182|2|3400000031|122|0.617360341382972|0|1|47|-80.782849|7|35.372142|REGISTER BARS|0.0|1|HERSHEY MILK CHOC BAR|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00034000002405|CANDY|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|32abf5e27187d3d37efca2c70d535e0a8d684c33|1.0|2015-01-30 22:22:00|1.4102725052409182|2|3400000031|122|0.617360341382972|0|1|47|-80.782849|7|35.372142|REGISTER BARS|0.25|1|HERSHEY MILK CHOC BAR|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00034000002405|CANDY|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|36fe6b6e328e986fe74f1d0fee4377ea02666191|1.0|2014-10-28 19:18:00|1.4102725052409182|2|3400000031|122|0.617360341382972|0|1|47|-80.782849|7|35.372142|REGISTER BARS|0.0|1|HERSHEY MILK CHOC BAR|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00034000002405|CANDY|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|103f9de53660126586f837f769fb5d7f2fd93bcd|1.0|2014-10-26 20:02:00|1.4102725052409182|2|3400000031|122|0.617360341382972|0|1|47|-80.782849|7|35.372142|REGISTER BARS|0.0|1|HERSHEY MILK CHOC BAR|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00034000002405|CANDY|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|30b64549aa87207c3fc6b3382a6e04f96d3e768b|1.0|2015-01-10 17:35:00|1.4102725052409182|2|3400000031|122|0.617360341382972|0|1|47|-80.782849|7|35.372142|REGISTER BARS|0.25|1|HERSHEY MILK CHOC BAR|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00034000002405|CANDY|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|da3ffa168a9a2ec8a74293059d4db3f0e4934479|11.15|2015-01-03 15:16:00|1.4102725052409182|2|3600040766|122|0.617360341382972|0|1|1205|-80.782849|67|35.372142|NFS-JUMBO DIAPERS|2.16|1|HUGGIES SLIP ON JUMBO 4|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00036000258097|DISPOSABLE DIAPERS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|8cfbb5da6ae86853072f652ec6118de79e6bf3ab|11.15|2014-12-28 09:15:00|1.4102725052409182|2|3600040766|122|0.617360341382972|0|1|1205|-80.782849|67|35.372142|NFS-JUMBO DIAPERS|2.16|1|HUGGIES SLIP ON JUMBO 4|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00036000258097|DISPOSABLE DIAPERS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|a7219d35bbbfc7ff41f955d03265003e4a3fbc92|4.99|2014-11-01 19:05:00|1.4102725052409182|2|2840008313|122|0.617360341382972|0|1|204|-80.782849|31|35.372142|TORTILLA CHIPS|1.0|1|TOSTITOS SCOOPS|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00028400083140|SNACKS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|ccd70c4a1448d2994299e61f10fce721b245631c|3.99|2015-01-21 19:07:00|1.4102725052409182|2|7433610006|122|0.617360341382972|0|1|342|-80.782849|57|35.372142|FRESH MILK|0.0|3|HUNTER 2%  MILK GALLON|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00074336100222|MILK|DAIRY|-80.782849|1.4099266941914086|122|1
35.372142|5111312b94659b804ae47033b771d9014fa93442|2.19|2014-12-11 17:58:00|1.4102725052409182|2|67293571020|122|0.617360341382972|0|1|4046|-80.782849|1080|35.372142|TOOTH BRUSH-CHILD|0.0|17|PEANUTS TBRUSH 4PK|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00672935710202|ORAL HYGIENE|HBC|-80.782849|1.4099266941914086|122|1
35.372142|0d0572d3ea8c7d16ba2a13deaae9ebcbf7e5e4c8|17.99|2015-02-23 19:37:00|1.4102725052409182|2|60240661584|122|0.617360341382972|0|1|5488|-80.782849|1502|35.372142|VILLAGE CANDLES|8.0|18|VCDECOR 18OZ TROPICAL GETAWAY|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00602406611455|CANDLES|GM|-80.782849|1.4099266941914086|122|1
35.372142|0b0e5a2177676c0bba393ac62f5cf1badba72f00|2.49|2014-11-20 21:31:00|1.4102725052409182|2|3400000312|122|0.617360341382972|0|1|1146|-80.782849|229|35.372142|SYRUPS|0.0|1|HERSHEY CHOCOLATE SYRUP|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00034000003129|COCOAS CREAMERS SYRUPS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|0cf3b747f9ed7e4c014a3bdfdb622d730ea18ef7|3.99|2014-10-21 16:52:00|1.4102725052409182|2|7203663995|122|0.617360341382972|0|1|342|-80.782849|57|35.372142|FRESH MILK|0.0|3|HARRIS TEETER 2% MILK|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00072036639981|MILK|DAIRY|-80.782849|1.4099266941914086|122|1
35.372142|12b4ff846caf835cccac2a483b57c58a88f08eed|3.65|2014-09-29 08:57:00|80.779636304526477|2|3800059663|122|35.397000260101713|0|17|61|-80.764523|9|35.341927|RTE CEREAL ADULT|0.0|1|KELLOGG RAISIN BRAN CRUNCH|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|35.392509581117899|00038000870101|CEREAL|G1 GROCERY|-80.782849|80.78285603145379|220|1
35.372142|4f2327cd0a8daf2a7b5fd124712f4bef572c9cc9|2.99|2014-12-28 15:25:00|1.4102725052409182|2|7203663217|122|0.617360341382972|0|1|330|-80.782849|55|35.372142|EGGS|0.0|3|HT GRADE A LARGE EGGS 18 CT|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00072036632173|EGGS FRESH|DAIRY|-80.782849|1.4099266941914086|122|1
35.372142|bae5fdba28eeb1334edeed3392fa918e4c07bb21|1.49|2015-01-04 19:13:00|1.4102725052409182|2|2840002819|122|0.617360341382972|0|1|206|-80.782849|31|35.372142|FRONT END SNACKS|0.0|1|CHEETOS CRUNCHY|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00028400028165|SNACKS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|689dd28912b2b205204f8e213df833fa2ac86a81|4.75|2014-11-02 17:07:00|1.4102725052409182|2|5170077050|122|0.617360341382972|0|1|388|-80.782849|66|35.372142|NFS-DISHWASH PWDR/LIQUID|0.0|1|FINISH POWER&FREE QUANT12CT|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00051700897124|DETERGENTS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|d8804153f65a3c62a2fa5b8310980a1f9492f7a0|1.0|2015-01-31 14:52:00|1.4102725052409182|2|4000000435|122|0.617360341382972|0|1|47|-80.782849|7|35.372142|REGISTER BARS|0.5|1|(FE)M&M PLAIN CANDY|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00040000000310|CANDY|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|3311e07d7efa90f4cdf31b00d64e2a63724049e8|1.0|2014-10-26 19:07:00|1.4102725052409182|2|4000000435|122|0.617360341382972|0|1|47|-80.782849|7|35.372142|REGISTER BARS|0.0|1|(FE)M&M PLAIN CANDY|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00040000000310|CANDY|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|35adc29ef2dd4980e91c8d6840b08a502343aad5|1.0|2014-12-22 16:57:00|1.4102725052409182|2|4000000435|122|0.617360341382972|0|1|47|-80.782849|7|35.372142|REGISTER BARS|0.2|1|(FE)M&M PLAIN CANDY|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00040000000310|CANDY|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.372142|22b2d368da155cd37c9543257e0db29b530fe6b7|2.39|2015-02-22 16:10:00|1.4102725052409182|2|1300000124|122|0.617360341382972|0|1|70|-80.782849|11|35.372142|KETCHUP|0.0|1|HEINZ KETCHUP 14 OZ|ebe254364f369079d1feff4ed47bbf9506faec4f|1.7176457881533291|0.61833652052202714|00013000001243|CONDIMENTS|G1 GROCERY|-80.782849|1.4099266941914086|122|1
35.04711|42823dc9177647b88db27b6f05528405fde9c7ef|4.29|2014-12-18 22:50:00|1.4091206135396188|1|2840016014|129|0.6116874628086298|0|47|201|-80.64817|31|35.04711|POTATO CHIPS|2.15|1|LAYS SALT & VINEGAR|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00028400160186|SNACKS|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|32bb265b4a3eb344a8e3ac5794a75f286beb5732|1.94|2014-11-01 12:38:00|1.4091206135396188|1|3100010903|129|0.6116874628086298|0|47|1279|-80.64817|48|35.04711|SINGLE SERVE FLAVOR|0.0|5|BANQUET TURKEY MEAL|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00031000109035|FROZEN MEALS|FROZEN|-80.64817|1.407576102208115|129|2
35.04711|07dd50a58e9af4cfe0e44a26be3ccb094bd233b2|2.58|2014-12-23 16:33:00|1.4091206135396188|1|2620011700|129|0.6116874628086298|0|47|206|-80.64817|31|35.04711|FRONT END SNACKS|0.58|1|SLIM JIM ORIGINAL GIANT|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00026200117003|SNACKS|G1 GROCERY|-80.64817|1.407576102208115|129|2
35.04711|eb02ac873a38017f426bad8a5cea25ec91b3648c|2.58|2014-12-08 21:25:00|1.4091206135396188|1|2620011700|129|0.6116874628086298|0|47|206|-80.64817|31|35.04711|FRONT END SNACKS|0.0|1|SLIM JIM ORIGINAL GIANT|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00026200117003|SNACKS|G1 GROCERY|-80.64817|1.407576102208115|129|2
35.04711|55445c4dfc8aea2346ccc7c49b22d4e4c1af6ae6|2.58|2015-02-21 19:57:00|1.4091206135396188|1|2620011700|129|0.6116874628086298|0|47|206|-80.64817|31|35.04711|FRONT END SNACKS|0.0|1|SLIM JIM ORIGINAL GIANT|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00026200117003|SNACKS|G1 GROCERY|-80.64817|1.407576102208115|129|2
35.04711|c4d639179206fea54d765824d54e7f5549e2f279|3.87|2015-01-03 16:37:00|1.4091206135396188|1|2620011700|129|0.6116874628086298|0|47|206|-80.64817|31|35.04711|FRONT END SNACKS|0.0|1|SLIM JIM ORIGINAL GIANT|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00026200117003|SNACKS|G1 GROCERY|-80.64817|1.407576102208115|129|3
35.04711|c0104536ebd5b2d0b5a3fbb6d662d5df5d6e6426|3.19|2015-02-27 19:37:00|1.4091206135396188|1|2733100032|129|0.6116874628086298|0|47|495|-80.64817|108|35.04711|NON REFRIGERATED|0.0|19|LA BANDERITA FLOUR TORTILLAS|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00027331000325|TORTILLAS|CASE READY MEATS|-80.64817|1.407576102208115|129|1
35.04711|b204ba4247f446d6232c0aee3a944fd501deeb63|1.29|2015-02-04 16:56:00|1.4091206135396188|1|2620011700|129|0.6116874628086298|0|47|206|-80.64817|31|35.04711|FRONT END SNACKS|0.0|1|SLIM JIM ORIGINAL GIANT|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00026200117003|SNACKS|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|eb04b77c31c062550be7c50e07bd0cc0b349699d|2.58|2014-11-22 20:14:00|1.4091206135396188|1|2620011700|129|0.6116874628086298|0|47|206|-80.64817|31|35.04711|FRONT END SNACKS|0.58|1|SLIM JIM ORIGINAL GIANT|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00026200117003|SNACKS|G1 GROCERY|-80.64817|1.407576102208115|129|2
35.04711|190818d183874d49302959f95ca0fb6404b2c60f|23.26|2015-01-21 19:34:00|1.4091206135396188|1|20140400000|129|0.6116874628086298|0|47|296|-80.64817|49|35.04711|RANCHER BEEF|9.7|2|BEEF LOIN NY STRIP STEAK BNLS|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00201404000003|BEEF|MEAT|-80.64817|1.407576102208115|129|1
35.04711|fffbbd9873f054af137a05da9ef9307a8776e0cd|2.58|2014-10-22 12:19:00|1.4091206135396188|1|5100002524|129|0.6116874628086298|0|47|179|-80.64817|27|35.04711|CANNED PASTA|0.58|1|SPAGHETTIOS PLUS CALCIUM|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00051000138194|PREPARED FOODS-RTS|G1 GROCERY|-80.64817|1.407576102208115|129|2
35.04711|327cc86f18a28f9717769b7f592cd8f6d99834a0|2.57|2015-01-04 18:26:00|1.4091206135396188|1|5150055003|129|0.6116874628086298|0|47|228|-80.64817|36|35.04711|TABLE SYRUP|1.26|1|HUNGRY JACK LITE PANCAKE SYRUP|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00051500550045|TABLE SYRUPS|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|e2112841b35063f80044583b1eb08ed304fedd67|2.97|2014-09-26 22:07:00|1.4091206135396188|1|5210009860|129|0.6116874628086298|0|47|75|-80.64817|34|35.04711|GRAVY MIXES|0.0|1|BROWN GRAVY LESS SODIUM|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00052100762494|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.64817|1.407576102208115|129|3
35.04711|672575ff8a6e5d155078729bae6e8d187ef1a8e9|0.97|2014-12-14 18:40:00|1.4091206135396188|1|7203697849|129|0.6116874628086298|0|47|1251|-80.64817|12|35.04711|WHOLESOME COOKIES|0.0|1|HT FIG BARS|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036978493|COOKIES|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|1da7bc2b0880fba93afda014ee80a73547293a2d|3.25|2015-01-01 18:36:00|1.4091206135396188|1|7203656080|129|0.6116874628086298|0|47|318|-80.64817|52|35.04711|SHREDDED/GRATED CHEESE|0.0|3|HT FANCY SHRED SHARP CHED CHE|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036550262|CHEESE|DAIRY|-80.64817|1.407576102208115|129|1
35.04711|e5400d04f3f80e178183abf1473c01769076fb27|6.98|2015-02-15 20:59:00|1.4091206135396188|1|7203660027|129|0.6116874628086298|0|47|361|-80.64817|105|35.04711|BREAKFAST SAUSAGE|0.99|19|HT BREAKFAST LINKS MAPLE|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036600301|BREAKFAST SAUSAGE|CASE READY MEATS|-80.64817|1.407576102208115|129|2
35.04711|ba61c0d136b5fa25d3fff0b2860061ffb436a428|6.5|2015-03-08 16:08:00|1.4091206135396188|1|7203656080|129|0.6116874628086298|0|47|318|-80.64817|52|35.04711|SHREDDED/GRATED CHEESE|0.0|3|HT FANCY SHRED SHARP CHED CHE|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036550262|CHEESE|DAIRY|-80.64817|1.407576102208115|129|2
35.04711|d5714bd3dc6278b858a5560aa70f625c52262faa|5.29|2014-11-06 18:30:00|1.4091206135396188|1|7203632028|129|0.6116874628086298|0|47|195|-80.64817|30|35.04711|SALAD & COOKING OIL|0.0|1|HT VEGETABLE OIL|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036320285|SHORTENING/OIL|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|9e860c5b5de6d382d7e469f8803a1f9c492c1e0d|2.85|2014-10-16 17:02:00|1.4091206135396188|1|7203604237|129|0.6116874628086298|0|47|41|-80.64817|6|35.04711|BREAKFAST BARS|1.19|1|HT BAR CEREAL BLUEBERRY|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036042392|BREAKFAST FOODS|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|24378388775a8df951088b768d2be802ac15f878|2.85|2015-01-22 18:43:00|1.4091206135396188|1|7203604237|129|0.6116874628086298|0|47|41|-80.64817|6|35.04711|BREAKFAST BARS|0.88|1|HT BAR CEREAL BLUEBERRY|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036042392|BREAKFAST FOODS|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|7d1be1d8b7cb8085d2c479cf214e73197696c6db|2.85|2015-01-28 12:19:00|1.4091206135396188|1|7203604237|129|0.6116874628086298|0|47|41|-80.64817|6|35.04711|BREAKFAST BARS|0.88|1|HT BAR CEREAL BLUEBERRY|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036042392|BREAKFAST FOODS|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|13c4ebee0cead113ce163b7334141e3d193bbbac|5.11|2014-10-15 18:33:00|1.4091206135396188|1|20165500000|129|0.6116874628086298|0|47|297|-80.64817|49|35.04711|GROUND BEEF|0.64|2|HT PREMIUM GRND BEEF 80% LEAN|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00201655000005|BEEF|MEAT|-80.64817|1.407576102208115|129|1
35.04711|5404951857801a88abd1de56085522bd5d89d416|6.26|2014-10-24 18:28:00|1.4091206135396188|1|20165500000|129|0.6116874628086298|0|47|297|-80.64817|49|35.04711|GROUND BEEF|0.47|2|HT PREMIUM GRND BEEF 80% LEAN|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00201655000005|BEEF|MEAT|-80.64817|1.407576102208115|129|1
35.04711|3e5461895d20d628a13859b259a3878c5f23eae0|7.0|2014-10-23 18:24:00|1.4091206135396188|1|7203698425|129|0.6116874628086298|0|47|254|-80.64817|892|35.04711|PREMIUM PIZZA|0.0|5|HT THIN CRUST PEPP/SAUS PIZZA|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036984265|FROZEN PIZZA|FROZEN|-80.64817|1.407576102208115|129|2
35.04711|57e8ffc0c2df04a3cf467f3d40d6957c9b409cb4|12.99|2015-02-07 18:52:00|1.4091206135396188|1|7203698519|129|0.6116874628086298|0|47|426|-80.64817|72|35.04711|NFS-PAPER TOWELS|3.0|1|YH ULT TOWEL 8RL SS WHITE|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036985200|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|531623ab765a7ecd6ac61d145e99a882cce05c67|3.14|2015-01-13 21:09:00|1.4091206135396188|1|7203697658|129|0.6116874628086298|0|47|44|-80.64817|6|35.04711|TOASTER PASTRIES-SHELF STABLE|0.0|1|HT TSTR PASTRY CHOC FUDGE|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036982230|BREAKFAST FOODS|G1 GROCERY|-80.64817|1.407576102208115|129|2
35.04711|56839891dc2843defcdae6ff4350064da7e36aac|2.59|2014-11-18 18:39:00|1.4091206135396188|1|7203695278|129|0.6116874628086298|0|47|1654|-80.64817|381|35.04711|DESSERT CAKES|0.0|14|DOUBLE FUDGE CAKE SLICE|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036952783|CAKES|BAKERY|-80.64817|1.407576102208115|129|1
35.04711|37169bfa411c54b1039da140dc5e6a664bc73527|7.49|2014-11-26 17:26:00|1.4091206135396188|1|7203695788|129|0.6116874628086298|0|47|1403|-80.64817|389|35.04711|THAW AND SELL PIES|2.5|14|"8"" PECAN PIE"|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036957887|PIES|BAKERY|-80.64817|1.407576102208115|129|1
35.04711|1b2bc9f8cf1d9cfd1124899a97fafc103e63d529|11.29|2015-02-23 20:43:00|1.4091206135396188|1|3600041241|129|0.6116874628086298|0|47|392|-80.64817|67|35.04711|NFS-DIAPER TRAINING PANT|1.8|1|GOODNITE BOY SMALL-MED JM 14CT|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00036000413137|DISPOSABLE DIAPERS|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|57627273298cf24893a2fa6606c41bc48ca23299|13.99|2015-01-10 22:00:00|1.4091206135396188|1|3410000342|129|0.6116874628086298|0|47|461|-80.64817|84|35.04711|FLAVORED MALT BEVERAGE|0.0|16|REDD'S WICKED ALE 12PK 10OZ CN|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00034100003425|SPECIALTY|BEER|-80.64817|1.407576102208115|129|1
35.04711|51837af9292ee5b4b60d0861022f227c9090c86c|11.29|2014-10-01 18:27:00|1.4091206135396188|1|3600041241|129|0.6116874628086298|0|47|392|-80.64817|67|35.04711|NFS-DIAPER TRAINING PANT|2.3|1|GOODNITE BOY SMALL-MED JM 14CT|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00036000413137|DISPOSABLE DIAPERS|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|48ea6391bbfa0980d06ead9c8a1fe7f5c987d03b|11.29|2014-10-08 18:55:00|1.4091206135396188|1|3600041241|129|0.6116874628086298|0|47|392|-80.64817|67|35.04711|NFS-DIAPER TRAINING PANT|2.3|1|GOODNITE BOY SMALL-MED JM 14CT|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00036000413137|DISPOSABLE DIAPERS|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|57e8b7266bb2e227da740dfc78243f362809c8a0|11.29|2014-09-26 18:23:00|1.4091206135396188|1|3600041241|129|0.6116874628086298|0|47|392|-80.64817|67|35.04711|NFS-DIAPER TRAINING PANT|2.3|1|GOODNITE BOY SMALL-MED JM 14CT|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00036000413137|DISPOSABLE DIAPERS|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|e80be54e40f7d041aac9f9dcc7ecfe10f90357d9|9.95|2015-02-06 20:25:00|1.4091206135396188|1|3114626257|129|0.6116874628086298|0|47|1217|-80.64817|273|35.04711|ASIAN MEAL KITS/MW|4.95|1|NONG SHIM BOWL PICANTE|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00031146250103|ASIAN PREP. FOODS|G1 GROCERY|-80.64817|1.407576102208115|129|5
35.04711|77e96945921eb88d31be0311a64faf6b12397960|11.29|2015-01-17 19:00:00|1.4091206135396188|1|3600041241|129|0.6116874628086298|0|47|392|-80.64817|67|35.04711|NFS-DIAPER TRAINING PANT|1.3|1|GOODNITE BOY SMALL-MED JM 14CT|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00036000413137|DISPOSABLE DIAPERS|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|876576fad02468bbee9b139f847ac5989560eb41|5.99|2014-11-05 18:41:00|1.4091206135396188|1|2100002492|129|0.6116874628086298|0|47|315|-80.64817|52|35.04711|CHEESE-PROCESSED-SLICED|2.02|3|KRAFT 2% AMERICAN SINGLE|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00021000024926|CHEESE|DAIRY|-80.64817|1.407576102208115|129|1
35.04711|98123a193cc93b7c63cb7ba345f37f63e41b14c9|1.58|2014-10-29 18:36:00|1.4091206135396188|1||129|0.6116874628086298|0|47|532|-80.64817|64|35.04711|FRESH CUCUMBERS|0.0|4|COO CUCUMBERS S/S|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00204062000002|FRESH PRODUCE|PRODUCE|-80.64817|1.407576102208115|129|2
35.04711|e7f93c3bde06194265234afbf26ffc1a0693aebc|7.59|2014-09-17 18:30:00|1.4091206135396188|1|1111112425|129|0.6116874628086298|0|47|726|-80.64817|73|35.04711|NFS-BODY WASHES|0.0|1|DOVE SHEA BUTTER BODYWASH|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00011111115224|PERSONAL SOAP/BATH ADDITIVES|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|839b8815269e9f9d3eb95dfb2e0943840aab24ee|1.67|2015-02-16 18:02:00|1.4091206135396188|1|7203697766|129|0.6116874628086298|0|47|325|-80.64817|54|35.04711|BISCUITS-REFRIGERATED|0.0|3|HT JUMBO BUTTERMILK BISC|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036977649|DOUGH PRODUCTS|DAIRY|-80.64817|1.407576102208115|129|1
35.04711|8e47facae02747fa550a4c5345216931c0d4cd1e|10.99|2015-02-09 18:51:00|1.4091206135396188|1|7203683001|129|0.6116874628086298|0|47|352|-80.64817|110|35.04711|IQF CHICKEN|2.21|19|HT 2.5 LB CHICKEN TENDR BRST|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036830029|FROZEN CASE MEAT|CASE READY MEATS|-80.64817|1.407576102208115|129|1
35.04711|3b4971177ec4b08544c6d28e0abbb3b955d8a3b2|1.2|2014-11-16 18:22:00|1.4091206135396188|1|3663203732|129|0.6116874628086298|0|47|685|-80.64817|61|35.04711|GREEK|0.2|3|DANNON LNF GREEK CHOC CHERRY|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00036632037503|YOGURT|DAIRY|-80.64817|1.407576102208115|129|1
35.04711|11fb3d3aba98a5b2c481bb237f82732b26f480c2|4.99|2014-10-26 18:02:00|1.4091206135396188|1|4260847021|129|0.6116874628086298|0|47|139|-80.64817|20|35.04711|REMAINING SHELF STABLE JUICES|0.0|1|LAKEWOOD HH POMEGRANT W/BLUBRY|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00042608470212|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|74a5fe05fbd79ce48e7110f9066c5cd06a9c75c5|3.97|2014-09-10 18:24:00|1.4091206135396188|1|7203658035|129|0.6116874628086298|0|47|358|-80.64817|100|35.04711|REGULAR BACON|0.97|19|HT REGULAR SLICED BACON|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036580351|BACON|CASE READY MEATS|-80.64817|1.407576102208115|129|1
35.04711|85d4818b323eca3084102b33fe35684e9f0d237a|5.99|2014-12-31 19:07:00|1.4091206135396188|1|7203658015|129|0.6116874628086298|0|47|1489|-80.64817|100|35.04711|STACK PACK BACON|0.0|19|HT MARKET STYLE THICK BACON|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036580153|BACON|CASE READY MEATS|-80.64817|1.407576102208115|129|1
35.04711|0a376342b76bf867724cdd488a56f7440b35bcbb|2.49|2015-01-28 18:34:00|1.4091206135396188|1|61126999100|129|0.6116874628086298|0|47|97|-80.64817|8|35.04711|ENERGY DRINKS|0.49|23|CB RED BULL ENERGY DRINK|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00611269991000|CARBONATED BEVERAGES|BEVERAGE|-80.64817|1.407576102208115|129|1
35.04711|e732d553198b2f6d7d3848b3c940d764c2e498aa|2.19|2014-09-19 20:55:00|1.4091206135396188|1|1200000496|129|0.6116874628086298|0|47|54|-80.64817|8|35.04711|DIET|0.69|23|DIET PEPSI 2 LTR NR|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00012000002311|CARBONATED BEVERAGES|BEVERAGE|-80.64817|1.407576102208115|129|1
35.04711|78aab89b71e90f8e651a06b8994a9034637b8fdd|2.89|2014-10-11 18:48:00|1.4091206135396188|1|7225004919|129|0.6116874628086298|0|47|1025|-80.64817|162|35.04711|WHITE|0.0|7|NATOWN BUTTERBREAD|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072250049191|SLICED BREAD|COMMERCIAL BAKERY|-80.64817|1.407576102208115|129|1
35.04711|582d89d02c780939dd73a843fa383016d7f0b557|2.89|2014-10-03 18:16:00|1.4091206135396188|1|7225004919|129|0.6116874628086298|0|47|1025|-80.64817|162|35.04711|WHITE|0.0|7|NATOWN BUTTERBREAD|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072250049191|SLICED BREAD|COMMERCIAL BAKERY|-80.64817|1.407576102208115|129|1
35.04711|b0d8c886feac0017cbfd3ba5abaa6a29358dcb59|5.32|2014-10-28 19:09:00|1.4091206135396188|1|20229600000|129|0.6116874628086298|0|47|299|-80.64817|49|35.04711|ANGUS BEEF|0.41|2|ANGUS BEEF EYE OF ROUND STEAK|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00202296000003|BEEF|MEAT|-80.64817|1.407576102208115|129|1
35.04711|fbfcd19c6102324292330e25033ba8efe556c496|1.25|2014-09-12 18:40:00|1.4091206135396188|1||129|0.6116874628086298|0|47|502|-80.64817|64|35.04711|FRESH BANANAS|0.0|4|BANANAS, YELLOW|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00204011000008|FRESH PRODUCE|PRODUCE|-80.64817|1.407576102208115|129|1
35.04711|f38a50d67da27db335863f8d217dca2fbfcc3e6a|1.47|2014-11-19 18:44:00|1.4091206135396188|1||129|0.6116874628086298|0|47|502|-80.64817|64|35.04711|FRESH BANANAS|0.0|4|BANANAS, YELLOW|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00204011000008|FRESH PRODUCE|PRODUCE|-80.64817|1.407576102208115|129|1
35.04711|b5e2ad2a8c8560beb64fc0e5f31806ad8ca4115d|1.49|2014-09-18 18:23:00|1.4091206135396188|1|20406100000|129|0.6116874628086298|0|47|525|-80.64817|64|35.04711|FRESH LETTUCE|0.0|4|ICEBERG LETTUCE|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00033383650203|FRESH PRODUCE|PRODUCE|-80.64817|1.407576102208115|129|1
35.04711|aaa21033fac3992e000a65a98e3775a05187cae7|8.59|2014-12-10 17:44:00|1.4091206135396188|1|7431207580|129|0.6116874628086298|0|47|4582|-80.64817|1215|35.04711|SPLMNT-WOMENS|0.0|17|NB HAIR SKIN AND NAILS|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00074312075803|VITAMINS & SUPPLEMENTS|HBC|-80.64817|1.407576102208115|129|1
35.04711|ca9e7c7321b2787ebda071feec859f2d52e624a2|7.39|2015-01-24 12:06:00|80.632521683083056|1|7527895005|129|35.21801023446762|0|39|1277|-80.699686|279|35.000049|FROZEN SNACKS|0.0|5|FSTR FRM MINI CRN DOGS 40-44CT|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|35.177497916598789|00075278950388|FROZEN SANDWICH AND SNACKS|FROZEN|-80.64817|80.648321474061262|249|1
35.04711|2336474c6175bc7dba58acd0977e466e7e049476|8.99|2014-11-12 18:41:00|1.4091206135396188|1|7199009511|129|0.6116874628086298|0|47|458|-80.64817|82|35.04711|CRAFT BEER|0.0|16|BLUE MOON BELGIAN WHT ALE 6PK|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00071990095116|DOMESTIC BEER|BEER|-80.64817|1.407576102208115|129|1
35.04711|10ce5eedc5861cfb604e5de05b1769b47f686204|5.99|2015-01-16 19:47:00|1.4091206135396188|1|7756725423|129|0.6116874628086298|0|47|252|-80.64817|45|35.04711|PREMIUM ICE CREAM|3.0|5|BREYERS MINT CHOC CHIP I/C|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00077567254245|ICE CREAM|FROZEN|-80.64817|1.407576102208115|129|1
35.04711|584b05af58b2c99d83b5fd5653946e4d1e1001a6|2.55|2014-09-29 18:30:00|1.4091206135396188|1|7535511228|129|0.6116874628086298|0|47|130|-80.64817|20|35.04711|CRANBERRY JUICE/DRINKS-SHELF|0.55|1|HEALTHY BALANCE POM/CRNBRY|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00075355111749|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|181ba91f0ca918c530b389d49ec650b22d917383|2.29|2015-01-20 18:52:00|1.4091206135396188|1|7800023046|129|0.6116874628086298|0|47|55|-80.64817|8|35.04711|REGULAR|0.79|23|CHEERWINE 2 LTR NR|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00070925000300|CARBONATED BEVERAGES|BEVERAGE|-80.64817|1.407576102208115|129|1
35.04711|6584419f5e97946f258407ca556d4da9bdc1562f|2.29|2014-12-06 19:56:00|1.4091206135396188|1|7800023046|129|0.6116874628086298|0|47|55|-80.64817|8|35.04711|REGULAR|1.29|23|CHEERWINE 2 LTR NR|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00070925000300|CARBONATED BEVERAGES|BEVERAGE|-80.64817|1.407576102208115|129|1
35.04711|5dfa89102361bcd5a38c82acc4ca2d23e53c59ce|3.79|2015-01-09 16:36:00|1.4091206135396188|1|7774529186|129|0.6116874628086298|0|47|555|-80.64817|64|35.04711|PACKAGED SALADS|0.3|4|R.P. BISTRO CRANBERRY WALNUT|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00077745294131|FRESH PRODUCE|PRODUCE|-80.64817|1.407576102208115|129|1
35.04711|ba3ac8354ca62f4f4fbbe12a65aee3a0f05b30c5|7.99|2015-02-01 18:16:00|1.4091206135396188|1|1820022979|129|0.6116874628086298|0|47|463|-80.64817|84|35.04711|HARD CIDER|0.0|16|JOHNNY APPLESEED 6PK|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00018200229794|SPECIALTY|BEER|-80.64817|1.407576102208115|129|1
35.04711|f934991be15f4e802cfb3ee244686e2cec9f83ed|1.34|2015-02-13 22:09:00|1.4091206135396188|1|7203660058|129|0.6116874628086298|0|47|325|-80.64817|54|35.04711|BISCUITS-REFRIGERATED|0.0|3|HT TEXAS STYLE BUTTER BISCUITS|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036600585|DOUGH PRODUCTS|DAIRY|-80.64817|1.407576102208115|129|1
35.04711|036115cd7b94d3e35b5560e6560e9a411457f8db|11.99|2014-12-02 18:40:00|1.4091206135396188|1|7203663048|129|0.6116874628086298|0|47|297|-80.64817|49|35.04711|GROUND BEEF|1.0|2|93% LEAN GROUND BEEF 2 LB|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036630483|BEEF|MEAT|-80.64817|1.407576102208115|129|1
35.04711|3cdf4ace43dbccb5d90bc1dc72b973f266488cb6|4.39|2014-10-05 18:48:00|1.4091206135396188|1|7433610006|129|0.6116874628086298|0|47|342|-80.64817|57|35.04711|FRESH MILK|0.0|3|HUNTER 2%  MILK GALLON|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00074336100222|MILK|DAIRY|-80.64817|1.407576102208115|129|1
35.04711|e634d1df052bbbb00298b672c64ed78e724a95e9|5.99|2015-01-26 18:39:00|1.4091206135396188|1|8500001707|129|0.6116874628086298|0|47|9939|-80.64817|885|35.04711|NFS POP PINOT NOIR|0.0|13|BAREFOOT PINOT NOIR|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00085000017074|POPULAR (4-$7.99)|WINE|-80.64817|1.407576102208115|129|1
35.04711|de5cfa9f63fed24b7a10bbaae3c7f33af01eeded|7.98|2014-11-25 16:05:00|1.4091206135396188|1|7218063244|129|0.6116874628086298|0|47|254|-80.64817|892|35.04711|PREMIUM PIZZA|0.0|5|RED BARON FRENCH BREAD PEP|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072180632449|FROZEN PIZZA|FROZEN|-80.64817|1.407576102208115|129|2
35.04711|c97797a5280c0c57433e9ce11af7fa70777f4f54|7.98|2014-11-05 18:35:00|1.4091206135396188|1|7218063244|129|0.6116874628086298|0|47|254|-80.64817|892|35.04711|PREMIUM PIZZA|0.0|5|RED BARON FRENCH BREAD PEP|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072180632449|FROZEN PIZZA|FROZEN|-80.64817|1.407576102208115|129|2
35.04711|3f8809ee26752896febd42e5be12f051928d0848|8.99|2015-03-02 21:12:00|1.4091206135396188|1|85337000208|129|0.6116874628086298|0|47|458|-80.64817|82|35.04711|CRAFT BEER|0.0|16|LONERIDER SWEET JOSIE 24/12|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00853370002088|DOMESTIC BEER|BEER|-80.64817|1.407576102208115|129|1
35.04711|b9534e153a658ce711ac94032aa39551ae68428a|7.99|2014-12-08 18:42:00|1.4091206135396188|1|1497450009|129|0.6116874628086298|0|47|463|-80.64817|84|35.04711|HARD CIDER|0.0|16|WOODCHUCK AMBER 6PK|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00014974500091|SPECIALTY|BEER|-80.64817|1.407576102208115|129|1
35.04711|d72b20f002174a365e61ea5977342e06d0b93225|8.99|2015-01-29 18:36:00|1.4091206135396188|1|1497450009|129|0.6116874628086298|0|47|463|-80.64817|84|35.04711|HARD CIDER|0.0|16|WOODCHUCK AMBER 6PK|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00014974500091|SPECIALTY|BEER|-80.64817|1.407576102208115|129|1
35.04711|a669c8384a0445cedd99508af8ca358e441ba2b6|8.99|2015-02-25 15:29:00|1.4091206135396188|1|1497450009|129|0.6116874628086298|0|47|463|-80.64817|84|35.04711|HARD CIDER|0.0|16|WOODCHUCK AMBER 6PK|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00014974500091|SPECIALTY|BEER|-80.64817|1.407576102208115|129|1
35.04711|8789a7b53279a925dab2f1b4a62b6430021c087f|6.89|2015-02-20 18:34:00|1.4091206135396188|1|7192196239|129|0.6116874628086298|0|47|284|-80.64817|892|35.04711|SUPER PREMIUM PIZZA|0.0|5|DIGIORNO 12in TC PEPPERONI|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00071921006594|FROZEN PIZZA|FROZEN|-80.64817|1.407576102208115|129|1
35.04711|58a25125eb10d7b11e4f45e4393537995ca0b05d|13.98|2015-03-04 18:46:00|1.4091206135396188|1|2500005838|129|0.6116874628086298|0|47|54|-80.64817|8|35.04711|DIET|3.5|23|MM L'ADE LIGHT 12OZ 12PK FP CN|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00025000058998|CARBONATED BEVERAGES|BEVERAGE|-80.64817|1.407576102208115|129|2
35.04711|5cb0d50cc40acdef45cd82aa127c552913a5b428|10.99|2015-02-17 21:19:00|1.4091206135396188|1|1834115101|129|0.6116874628086298|0|47|9935|-80.64817|885|35.04711|NFS POP CAB SAUV|0.0|13|BAREFOOT CAB SAUV 1.5L|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00018341151015|POPULAR (4-$7.99)|WINE|-80.64817|1.407576102208115|129|1
35.04711|6a6e81595cd226118d008c7f4a01de74d6c21b39|10.99|2015-02-10 20:49:00|1.4091206135396188|1|1834115101|129|0.6116874628086298|0|47|9935|-80.64817|885|35.04711|NFS POP CAB SAUV|0.0|13|BAREFOOT CAB SAUV 1.5L|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00018341151015|POPULAR (4-$7.99)|WINE|-80.64817|1.407576102208115|129|1
35.04711|b891882dc64404dd78a36dafa3cfa30d36b18825|9.38|2015-01-14 18:27:00|1.4091206135396188|1|7047046158|129|0.6116874628086298|0|47|685|-80.64817|61|35.04711|GREEK|0.0|3|YOPLAIT GRK STRAWBRY BLEND 4PK|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00070470461564|YOGURT|DAIRY|-80.64817|1.407576102208115|129|2
35.04711|69702492ff9c2b2d63b55d28e92661e78a9337c9|4.59|2015-02-18 18:33:00|1.4091206135396188|1|2740026499|129|0.6116874628086298|0|47|313|-80.64817|51|35.04711|MARGARINE|0.0|3|COUNTRY CROCK PLUS CALCIUM|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00027400264955|BUTTER & MARGARINE|DAIRY|-80.64817|1.407576102208115|129|1
35.04711|b0c2e6e62c51544d296e085f023d0268b299e1d9|8.39|2014-09-13 17:15:00|1.4091206135396188|1|3600016792|129|0.6116874628086298|0|47|1207|-80.64817|67|35.04711|NFS-WIPES|2.4|1|HUG WIP OD SCENT 3X REFILL 184|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00036000167924|DISPOSABLE DIAPERS|G1 GROCERY|-80.64817|1.407576102208115|129|1
35.04711|6ca181af7d6070044203d68dbd5676c7449b13e7|4.99|2014-10-05 12:22:00|80.632521683083056|1|7244010400|129|35.218010271732581|0|39|6787|-80.825175|1568|35.152722|MAGAZINES MONTHLY|0.0|18|SOUTHERN LIVING|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|35.177497916598789|00072440104006|MAGAZINES|GM|-80.64817|80.648232453931328|160|1
35.04711|8e3f1ab686e928e18c3d44ef02849ee0e7b142f4|9.3|2015-01-27 18:35:00|1.4091206135396188|1|7218063473|129|0.6116874628086298|0|47|254|-80.64817|892|35.04711|PREMIUM PIZZA|2.63|5|RED BARON THN CRUST PEPPERONI|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072180633224|FROZEN PIZZA|FROZEN|-80.64817|1.407576102208115|129|2
35.04711|3d98038f4e8d91eef1e6a7dc825026a4dc83e673|7.98|2014-09-22 18:28:00|1.4091206135396188|1|7203663995|129|0.6116874628086298|0|47|342|-80.64817|57|35.04711|FRESH MILK|0.0|3|HARRIS TEETER 2% MILK|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036639981|MILK|DAIRY|-80.64817|1.407576102208115|129|2
35.04711|b8a3b3d8a396d863bc74d2dc4d327c809943ff55|6.98|2015-02-03 18:34:00|1.4091206135396188|1|7203663995|129|0.6116874628086298|0|47|342|-80.64817|57|35.04711|FRESH MILK|0.0|3|HARRIS TEETER 2% MILK|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036639981|MILK|DAIRY|-80.64817|1.407576102208115|129|2
35.04711|9a752e0c0494d6fc839abdf89d27f7df10e72cc2|7.98|2014-10-19 18:46:00|1.4091206135396188|1|7203663995|129|0.6116874628086298|0|47|342|-80.64817|57|35.04711|FRESH MILK|0.0|3|HARRIS TEETER 2% MILK|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036639981|MILK|DAIRY|-80.64817|1.407576102208115|129|2
35.04711|e7f4dd890180797188f3db3ee7fde105273c2474|5.61|2014-10-20 20:22:00|1.4091206135396188|1|7203670901|129|0.6116874628086298|0|47|214|-80.64817|33|35.04711|BROTH|0.0|1|HT REDUC SOD CHICKN BROTH 32OZ|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036709028|SOUP|G1 GROCERY|-80.64817|1.407576102208115|129|3
35.04711|2a577f3ce6db700befe4bcedea4dc3c35b4ec54b|15.19|2014-10-23 22:09:00|1.4091206135396188|1|33160414271|129|0.6116874628086298|0|47|4579|-80.64817|1215|35.04711|SPLMNT-URINARY DSCMFRT|0.0|17|NM CRANBERRY SUP-STR SFTGEL|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00331604142712|VITAMINS & SUPPLEMENTS|HBC|-80.64817|1.407576102208115|129|1
35.04711|edf95b75da8e4babba1474121a514d4ed8175805|7.98|2014-09-15 18:38:00|1.4091206135396188|1|7203663995|129|0.6116874628086298|0|47|342|-80.64817|57|35.04711|FRESH MILK|0.0|3|HARRIS TEETER 2% MILK|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036639981|MILK|DAIRY|-80.64817|1.407576102208115|129|2
35.04711|c5500a201583425302dae50afa7a0adc3cb8691e|7.98|2014-12-22 18:34:00|1.4091206135396188|1|7203663995|129|0.6116874628086298|0|47|342|-80.64817|57|35.04711|FRESH MILK|0.0|3|HARRIS TEETER 2% MILK|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036639981|MILK|DAIRY|-80.64817|1.407576102208115|129|2
35.04711|bfff90655dbe882c898907d1ac616763e0204bc1|10.99|2014-10-25 18:57:00|1.4091206135396188|1|8500001736|129|0.6116874628086298|0|47|9939|-80.64817|885|35.04711|NFS POP PINOT NOIR|0.0|13|BAREFOOT PINOT NOIR 1.5L|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00085000017364|POPULAR (4-$7.99)|WINE|-80.64817|1.407576102208115|129|1
35.04711|4631f9386edd9090c712fa03ce98dd4f8db382ce|21.98|2015-02-11 19:54:00|1.4091206135396188|1|8500001736|129|0.6116874628086298|0|47|9939|-80.64817|885|35.04711|NFS POP PINOT NOIR|0.0|13|BAREFOOT PINOT NOIR 1.5L|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00085000017364|POPULAR (4-$7.99)|WINE|-80.64817|1.407576102208115|129|2
35.04711|ede240905a26306ee3185b6d9b4c7eb45cc560cf|9.99|2015-01-14 18:24:00|1.4091206135396188|1|8500001736|129|0.6116874628086298|0|47|9939|-80.64817|885|35.04711|NFS POP PINOT NOIR|0.0|13|BAREFOOT PINOT NOIR 1.5L|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00085000017364|POPULAR (4-$7.99)|WINE|-80.64817|1.407576102208115|129|1
35.04711|7f295ce723b27b15936ca9604e6a3145de911842|10.99|2015-02-14 22:07:00|1.4091206135396188|1|8500001736|129|0.6116874628086298|0|47|9939|-80.64817|885|35.04711|NFS POP PINOT NOIR|0.0|13|BAREFOOT PINOT NOIR 1.5L|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00085000017364|POPULAR (4-$7.99)|WINE|-80.64817|1.407576102208115|129|1
35.04711|c5f9d87ad822f9de66673aa158effae35623b8bf|10.99|2014-10-09 18:22:00|1.4091206135396188|1|8500001736|129|0.6116874628086298|0|47|9939|-80.64817|885|35.04711|NFS POP PINOT NOIR|0.0|13|BAREFOOT PINOT NOIR 1.5L|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00085000017364|POPULAR (4-$7.99)|WINE|-80.64817|1.407576102208115|129|1
35.04711|f5bcc4d3350dad5177297a7935de7eff2ee8981d|2.29|2014-09-25 20:52:00|1.4091206135396188|1|7800023046|129|0.6116874628086298|0|47|55|-80.64817|8|35.04711|REGULAR|0.79|23|CANADA DRY GINGER ALE NR 2LTR|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00078000152463|CARBONATED BEVERAGES|BEVERAGE|-80.64817|1.407576102208115|129|1
35.04711|1c17698e185e4ef01bc823c5610083d7838b9490|5.99|2015-01-23 21:11:00|1.4091206135396188|1|7704360805|129|0.6116874628086298|0|47|3196|-80.64817|1015|35.04711|HAND & BODY EVERYDAY|0.0|17|ST. IVES RENEW COLLAGEN BDY LT|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00077043608029|HAND & BODY LOTION/SUN CARE|HBC|-80.64817|1.407576102208115|129|1
35.04711|2871b14b8667563f7c2f6df52553109fac52b8de|1.37|2015-03-07 18:22:00|1.4091206135396188|1|7203690021|129|0.6116874628086298|0|47|1033|-80.64817|163|35.04711|HAMBURGER|0.0|7|H T HAMBURGER BUNS|f1bcfc21f6ca45c03e98fbcb2004b7ca29dbe15b|11.80879659472532|0.61242566243833529|00072036900210|BUNS/ROLLS|COMMERCIAL BAKERY|-80.64817|1.407576102208115|129|1
35.667941|12abac6e5827231e1b361b2b2dd616521164c4b8|9.7|2014-11-22 14:01:00|1.4057311447477159|4|3450015136|178|0.6225230078570788|0|52|312|-80.497332|51|35.667941|BUTTER|2.7|3|L O L BUTTER QUARTERS|f223520292e44026b47a591dd6be4c4a811e1854|3.7224787569137314|0.6209993146566879|00034500151368|BUTTER & MARGARINE|DAIRY|-80.497332|1.4049434824709919|178|2
35.667941|8a57317a7bff987e4bfdc6f4bce5536cb858ad98|18.98|2014-10-14 12:09:00|1.4057311447477159|4|5400011971|178|0.6225230078570788|0|52|427|-80.497332|72|35.667941|NFS-TOILET TISSUE|5.0|1|SCOTT 1000 WHITE 8 ROLL|f223520292e44026b47a591dd6be4c4a811e1854|3.7224787569137314|0.6209993146566879|00054000119712|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.497332|1.4049434824709919|178|2
35.667941|f5187abb83e7eeea3d70122e0151fdda498996cf|5.0|2014-11-26 16:58:00|1.4057311447477159|4|812|178|0.6225230078570788|0|52|1639|-80.497332|377|35.667941|BULK (DONUTS)|0.0|14|NEW BULK DONUT CODE|f223520292e44026b47a591dd6be4c4a811e1854|3.7224787569137314|0.6209993146566879|00000000008120|DONUTS|BAKERY|-80.497332|1.4049434824709919|178|5
34.95459|bc4281ae0787b11ad0925dbaebcb60c70360efe2|13.29|2014-12-10 07:53:00|1.4091206135396188|4|3700013882|182|0.6100726841846847|0|47|389|-80.758228|66|34.95459|NFS-LAUNDRY DETERGENTS|0.0|1|TIDE HE ORIGINAL 64 LD|fa32b88e325c47cb81b86f34bebcd1463acb840c|2.9422155896675766|0.61242566243833529|00037000088868|DETERGENTS|G1 GROCERY|-80.758228|1.4094969766762753|182|1
34.95459|8bff947ab45184a0566e2ce8830deabb473c8f74|3.99|2014-12-22 16:03:00|1.4091206135396188|4|70935189147|182|0.6100726841846847|0|47|556|-80.758228|64|34.95459|PACKAGED VEGETABLES|0.0|4|APIO GINGER BOK CHOY SALAD|fa32b88e325c47cb81b86f34bebcd1463acb840c|2.9422155896675766|0.61242566243833529|00709351891472|FRESH PRODUCE|PRODUCE|-80.758228|1.4094969766762753|182|1
34.95459|490ee7b41ac29380e423cda033d2347ae2db88d1|3.99|2014-10-08 13:41:00|80.758271881003409|4|70935189147|182|34.997170578676815|0|28|556|-80.837892|64|34.937113|PACKAGED VEGETABLES|0.0|4|APIO GINGER BOK CHOY SALAD|fa32b88e325c47cb81b86f34bebcd1463acb840c|2.9422155896675766|34.992988447249964|00709351891472|FRESH PRODUCE|PRODUCE|-80.758228|80.758256144608112|372|1
34.95459|af303dc49592d7e407b8cc8f7c09dea20149aa8c|3.99|2014-10-17 11:08:00|1.4091206135396188|4|70935189147|182|0.6100726841846847|0|47|556|-80.758228|64|34.95459|PACKAGED VEGETABLES|0.0|4|APIO GINGER BOK CHOY SALAD|fa32b88e325c47cb81b86f34bebcd1463acb840c|2.9422155896675766|0.61242566243833529|00709351891472|FRESH PRODUCE|PRODUCE|-80.758228|1.4094969766762753|182|1
34.95459|2b93147f34af54bfbe6a7ff5b52af3c7caa276a9|4.39|2014-09-13 19:00:00|1.4091206135396188|4|81857000851|182|0.6100726841846847|0|47|722|-80.758228|73|34.95459|NFS-HAND SOAPS|0.4|1|WATKINS LEMON LIQ SOAP|fa32b88e325c47cb81b86f34bebcd1463acb840c|2.9422155896675766|0.61242566243833529|00818570008520|PERSONAL SOAP/BATH ADDITIVES|G1 GROCERY|-80.758228|1.4094969766762753|182|1
34.95459|89a369fb98dd08085dad985e293795ff817c20bb|3.38|2014-10-03 12:46:00|1.4091206135396188|4|2100065897|182|0.6100726841846847|0|47|1441|-80.758228|274|34.95459|MAC AND CHEESE|1.38|1|KRAFT MAC CHEESE NINJA TURTLE|fa32b88e325c47cb81b86f34bebcd1463acb840c|2.9422155896675766|0.61242566243833529|00021000031542|PREP FOODS DINNERS|G1 GROCERY|-80.758228|1.4094969766762753|182|2
34.95459|1ebdc2dcb4114e4d65e74da70ae60441b2f23d23|4.99|2015-01-29 17:11:00|1.4091206135396188|4|78142152480|182|0.6100726841846847|0|47|1601|-80.758228|371|34.95459|BRANDED BREAD|2.0|14|LA BREA THREE CHEESE SEMOLINA|fa32b88e325c47cb81b86f34bebcd1463acb840c|2.9422155896675766|0.61242566243833529|00781421524800|BREAD|BAKERY|-80.758228|1.4094969766762753|182|1
34.95459|2a4310cfd8986203304abee5a86e0102c30fe085|3.95|2015-01-31 17:58:00|80.758271881003409|4|95546|182|34.997170578676815|0|28|1582|-80.837892|369|34.937113|NFS BEVERAGE TEA|0.0|22|CHAI TEA LATTE GRANDE|fa32b88e325c47cb81b86f34bebcd1463acb840c|2.9422155896675766|34.992988447249964|00000000955460|NFS STARBUCKS|COFFEE SHOP|-80.758228|80.758256144608112|372|1
34.95459|186197ad2870387ff67bedf6d8ca5228d301c430|2.85|2015-02-25 13:03:00|1.4091206135396188|4||182|0.6100726841846847|0|47|500|-80.758228|64|34.95459|FRESH APPLES|0.0|4|GOLD DEL APPLE, WA 56|fa32b88e325c47cb81b86f34bebcd1463acb840c|2.9422155896675766|0.61242566243833529|00233285000001|FRESH PRODUCE|PRODUCE|-80.758228|1.4094969766762753|182|1
34.95459|ac5f4718f59a959824c9b08bb1a3a0b547b10383|2.49|2015-01-31 17:56:00|80.758271881003409|4|3400019045|182|34.997170578676815|0|28|46|-80.837892|7|34.937113|PKG CHOC|0.0|1|HSY MILK CHOC GIANT BAR|fa32b88e325c47cb81b86f34bebcd1463acb840c|2.9422155896675766|34.992988447249964|00034000190454|CANDY|G1 GROCERY|-80.758228|80.758256144608112|372|1
34.95459|6c701c7aa06bfb3e5740a17fc8445cf55952e462|4.99|2015-01-31 11:21:00|1.4091206135396188|4|2301290130|182|0.6100726841846847|0|47|1477|-80.758228|485|34.95459|SUSHI HYBRID|0.0|6|CALIFORNIA ROLL SP|fa32b88e325c47cb81b86f34bebcd1463acb840c|2.9422155896675766|0.61242566243833529|00023012901301|SUSHI|DELI|-80.758228|1.4094969766762753|182|1
34.95459|e764e81e52ac8c6bb520a3d6354dd8e74d2e6c14|1.19|2015-02-01 11:26:00|1.4091206135396188|4|5210004606|182|0.6100726841846847|0|47|734|-80.758228|3|34.95459|NFS-CANDLES/BIRTHDAY SUP|0.0|1|MC POLKA DOT CANDLES|fa32b88e325c47cb81b86f34bebcd1463acb840c|2.9422155896675766|0.61242566243833529|00052100047126|BAKING SUPPLIES|G1 GROCERY|-80.758228|1.4094969766762753|182|1
34.95459|3cd917cb634b3b688bf7b7bf0745109ac0c97105|2.5|2015-02-05 18:55:00|80.758271881003409|4|7203695815|182|34.997170576682173|0|28|1687|-80.848528|385|35.053394|THAW & SELL (SWEET GOODS)|0.0|14|Bulk Pastry No Tax Each|fa32b88e325c47cb81b86f34bebcd1463acb840c|2.9422155896675766|34.992988447249964|00072036958150|SWEET GOODS|BAKERY|-80.758228|80.758260328301802|11|1
34.95459|2847fffbc0f4952fe7cddf76f7e23741eb91dda9|3.99|2014-09-21 12:46:00|1.4091206135396188|4|70935189142|182|0.6100726841846847|0|47|556|-80.758228|64|34.95459|PACKAGED VEGETABLES|0.0|4|APIO KALE SALAD KIT|fa32b88e325c47cb81b86f34bebcd1463acb840c|2.9422155896675766|0.61242566243833529|00709351891427|FRESH PRODUCE|PRODUCE|-80.758228|1.4094969766762753|182|1
35.082768|f3f900167baa31363904e201718994d92d778a83|7.75|2014-11-09 17:16:00|1.4091206135396188|1|1258760034|147|0.6123098123133061|0|47|443|-80.732725|76|35.082768|NFS-GARBAGE BAGS|0.0|1|GLAD TALL KIT DRAWSTRING 45 CT|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00012587783627|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.732725|1.409051865357139|147|1
35.082768|737861af60fb9a96978ee57ed0502f117224f899|9.99|2015-02-13 18:18:00|1.4091206135396188|1|85768000107|147|0.6123098123133061|0|47|9969|-80.732725|887|35.082768|NFS-S/PREM-OTHER RED|0.0|13|SHANNON RIDGE WRANGLER RED|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00857680001076|SUPER PREMIUM ($11-$14.99)|WINE|-80.732725|1.409051865357139|147|1
35.082768|e6ad9d5ec8735a174f5580396dbaa557212ab186|3.29|2014-12-15 09:04:00|1.4091206135396188|1|1600048772|147|0.6123098123133061|0|47|74|-80.732725|9|35.082768|RTE CEREAL ALL FAMILY|0.0|1|GM CHEERIOS 12 OZ|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00016000487727|CEREAL|G1 GROCERY|-80.732725|1.409051865357139|147|1
35.082768|f54ea38f89991c1cb80662849c8b7c30fb95b7f8|2.99|2015-02-28 17:27:00|80.732732175546019|1||147|35.099021295261316|0|35|542|-80.78468|64|35.096737|FRESH VEGETABLES REMAIN|0.0|4|COO ARTICHOKES, JBO (RPC)|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00204084000004|FRESH PRODUCE|PRODUCE|-80.732725|80.732726780676799|30|1
35.082768|b4894c8adf502dcd6ef7b02852c14548b3e79467|7.99|2014-12-09 21:05:00|1.4091206135396188|1||147|0.6123098123133061|0|47|506|-80.732725|64|35.082768|FRESH MELONS|0.0|4|WATERMELON, BIN|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00204032000001|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|1
35.082768|1a4c02e9862552f0bbe9ab0c5421741aec573910|2.49|2014-10-06 13:10:00|1.4091206135396188|1|7047044346|147|0.6123098123133061|0|47|682|-80.732725|61|35.082768|KIDS|0.49|3|TRIX STRAWBERRY PUNCH 4CT|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00070470443461|YOGURT|DAIRY|-80.732725|1.409051865357139|147|1
35.082768|c79b6f10aeb95082bc96fbb4de123915db9cce1a|2.49|2014-11-03 17:55:00|1.4091206135396188|1|7047044346|147|0.6123098123133061|0|47|682|-80.732725|61|35.082768|KIDS|0.0|3|TRIX STRAWBERRY PUNCH 4CT|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00070470443461|YOGURT|DAIRY|-80.732725|1.409051865357139|147|1
35.082768|180b1a064aa07a1a9c1cae70a663a8b4835480e7|2.49|2015-01-11 13:14:00|1.4091206135396188|1|7047044346|147|0.6123098123133061|0|47|682|-80.732725|61|35.082768|KIDS|0.49|3|TRIX STRAWBERRY PUNCH 4CT|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00070470443461|YOGURT|DAIRY|-80.732725|1.409051865357139|147|1
35.082768|e8c1e3aad062b98e3d536039c509b1d4e9123ac4|2.49|2014-12-24 14:34:00|1.4091206135396188|1|7047044346|147|0.6123098123133061|0|47|682|-80.732725|61|35.082768|KIDS|0.0|3|TRIX STRAWBERRY PUNCH 4CT|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00070470443461|YOGURT|DAIRY|-80.732725|1.409051865357139|147|1
35.082768|2b7092548de59b89403ef4d67e25e32fa9cb8418|2.49|2014-11-24 18:14:00|80.732732175546019|1|7047044346|147|35.099021295261316|0|35|682|-80.78468|61|35.096737|KIDS|0.0|3|TRIX STRAWBERRY PUNCH 4CT|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00070470443461|YOGURT|DAIRY|-80.732725|80.732726780676799|30|1
35.082768|079b4cd3b7a6f50b6132b39208122494ea783ecb|2.49|2014-12-05 18:00:00|80.732732175546019|1|7047044346|147|35.099021295261316|0|35|682|-80.78468|61|35.096737|KIDS|0.0|3|TRIX STRAWBERRY PUNCH 4CT|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00070470443461|YOGURT|DAIRY|-80.732725|80.732726780676799|30|1
35.082768|e3f45b119b01252ec79cd4a26271f4f1ca673260|9.98|2015-01-08 13:49:00|1.4091206135396188|1|5150014192|147|0.6123098123133061|0|47|104|-80.732725|16|35.082768|APPLESAUCE-CUPS|2.5|1|SMKR FRUITFULLS APPLE 4PK|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00051500141786|FRUIT-CAN/JAR|G1 GROCERY|-80.732725|1.409051865357139|147|2
35.082768|2e3c144a7498c806673798bc3550361e5ed9c393|3.39|2015-01-22 17:56:00|1.4091206135396188|1|5260305445|147|0.6123098123133061|0|47|214|-80.732725|33|35.082768|BROTH|0.0|1|PACIFIC ORG LS FR CHICKN BROTH|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00052603054454|SOUP|G1 GROCERY|-80.732725|1.409051865357139|147|1
35.082768|0866e74d884feeddc9a6bbb7010dfec577cf1480|6.78|2015-02-16 11:42:00|80.732732175546019|1|5260305445|147|35.099021295261316|0|35|214|-80.78468|33|35.096737|BROTH|0.0|1|PACIFIC ORG LS FR CHICKN BROTH|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00052603054454|SOUP|G1 GROCERY|-80.732725|80.732726780676799|30|2
35.082768|ce9c105f304206d9899a13aeeef910b416fa579c|6.78|2014-12-31 12:28:00|1.4091206135396188|1|5260305445|147|0.6123098123133061|0|47|214|-80.732725|33|35.082768|BROTH|0.0|1|PACIFIC ORG LS FR CHICKN BROTH|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00052603054454|SOUP|G1 GROCERY|-80.732725|1.409051865357139|147|2
35.082768|bc7556a93654bed62a612a7c9ba5803cb68a1327|5.99|2015-02-08 17:36:00|80.732732175546019|1|7485108639|147|35.099021295261316|0|35|6790|-80.78468|1568|35.096737|MAGAZINES SEMI ANNUAL|0.0|18|08639 PP FAV XWD DISP|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00074851086391|MAGAZINES|GM|-80.732725|80.732726780676799|30|1
35.082768|e4d9df3d770848023f2de6ec3d8ab176c1d65edc|13.99|2014-10-25 17:18:00|80.732732175546019|1|8382012368|147|35.099021295261316|0|35|459|-80.78468|83|35.096737|IMPORT BEER|0.0|16|GUINNESS CN|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00083820123685|IMPORT BEER|BEER|-80.732725|80.732726780676799|30|1
35.082768|7bab2edc75b1c794a0a9a046ef7f13c60316f27f|9.99|2014-10-11 19:20:00|1.4091206135396188|1|8224252043|147|0.6123098123133061|0|47|9948|-80.732725|886|35.082768|NFS-PREM-CAB SAUVIGNON|0.0|13|HANDCRAFT CABERNET|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00082242520430|PREMIUM ($8-$10.99)|WINE|-80.732725|1.409051865357139|147|1
35.082768|a06303165aff62a3e3cb679dea905f9f69746606|13.99|2014-12-19 16:53:00|80.732732175546019|1|8382012368|147|35.099021295261316|0|35|459|-80.78468|83|35.096737|IMPORT BEER|0.0|16|GUINNESS CN|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00083820123685|IMPORT BEER|BEER|-80.732725|80.732726780676799|30|1
35.082768|23ec1244af146f0a0630165a237f8e346f4e18e5|9.99|2015-02-06 13:34:00|1.4091206135396188|1|8224252043|147|0.6123098123133061|0|47|9948|-80.732725|886|35.082768|NFS-PREM-CAB SAUVIGNON|0.0|13|HANDCRAFT CABERNET|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00082242520430|PREMIUM ($8-$10.99)|WINE|-80.732725|1.409051865357139|147|1
35.082768|c5587e1c5272e2d0d2daaa2672fbd37aedb72281|15.99|2014-09-19 18:00:00|80.732732175546019|1|8382012368|147|35.099021295261316|0|35|459|-80.78468|83|35.096737|IMPORT BEER|0.0|16|GUINNESS CN|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00083820123685|IMPORT BEER|BEER|-80.732725|80.732726780676799|30|1
35.082768|66210e7cabf55c1729a753a5e09ec1b7b303d462|15.99|2014-10-03 17:42:00|1.4091206135396188|1|8382012368|147|0.6123098123133061|0|47|459|-80.732725|83|35.082768|IMPORT BEER|0.0|16|GUINNESS CN|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00083820123685|IMPORT BEER|BEER|-80.732725|1.409051865357139|147|1
35.082768|08c9b1d9b445c8005c2e9eb0094a1df4eac8303e|5.78|2015-01-04 14:53:00|1.4091206135396188|1|3800040260|147|0.6123098123133061|0|47|1269|-80.732725|41|35.082768|BREAKFAST SYRUP CARRIER|0.78|5|EGGO HOMESTYLE WAFFLES|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00038000402609|BREAKFAST FOODS FROZEN|FROZEN|-80.732725|1.409051865357139|147|2
35.082768|49f88cf74f690b6608fed84db8e7a0d60583f707|2.89|2014-11-30 16:28:00|1.4091206135396188|1|3800040260|147|0.6123098123133061|0|47|1269|-80.732725|41|35.082768|BREAKFAST SYRUP CARRIER|0.0|5|EGGO HOMESTYLE WAFFLES|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00038000402609|BREAKFAST FOODS FROZEN|FROZEN|-80.732725|1.409051865357139|147|1
35.082768|03c9972793ac06d76468bcd2cf01dceeb18e6e2e|3.25|2014-11-16 17:31:00|1.4091206135396188|1|3620022302|147|0.6123098123133061|0|47|1219|-80.732725|275|35.082768|PASTA SC CORE|0.0|1|BERTOLLI SC ORG TOMATO BASIL|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00036200222843|PASTA SAUCES|G1 GROCERY|-80.732725|1.409051865357139|147|1
35.082768|23eb93e1694e40fc8e0faccc20461f7775be0aaa|7.98|2014-09-29 19:17:00|1.4091206135396188|1|3338324028|147|0.6123098123133061|0|47|504|-80.732725|64|35.082768|FRESH BERRIES|4.64|4|BLACKBERRIES 5.6 OZ|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00033383240268|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|2
35.082768|9659fde257d16a0d15851e5b89cb3ce1074a0b22|2.85|2015-01-27 17:46:00|80.732732175546019|1|3800040260|147|35.099021295261316|0|35|1269|-80.78468|41|35.096737|BREAKFAST SYRUP CARRIER|0.0|5|EGGO HOMESTYLE WAFFLES|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00038000402609|BREAKFAST FOODS FROZEN|FROZEN|-80.732725|80.732726780676799|30|1
35.082768|56d732e5dbd032e8d4757d471f08ea60e963f342|8.55|2015-03-06 18:06:00|80.732732175546019|1|3800040260|147|35.099021295261316|0|35|1269|-80.78468|41|35.096737|BREAKFAST SYRUP CARRIER|0.85|5|EGGO HOMESTYLE WAFFLES|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00038000402609|BREAKFAST FOODS FROZEN|FROZEN|-80.732725|80.732726780676799|30|3
35.082768|945bbd896c99e71cc070fe8aa24d61c5b49e8938|5.99|2014-09-15 12:52:00|1.4091206135396188|1|3338311008|147|0.6123098123133061|0|47|507|-80.732725|64|35.082768|FRESH ORANGES|0.0|4|NAVEL ORANGE FL 8LB BAG|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00033383146218|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|1
35.082768|853f734fa0e7fefe0e3527cd84cac54e5823830b|5.99|2014-10-12 17:16:00|1.4091206135396188|1|3338311008|147|0.6123098123133061|0|47|507|-80.732725|64|35.082768|FRESH ORANGES|0.0|4|NAVEL ORANGE FL 8LB BAG|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00033383146218|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|1
35.082768|86acda90e427d9a8dff437482f1b27d3a28fb748|13.98|2015-01-09 18:11:00|1.4091206135396188|1|3338324000|147|0.6123098123133061|0|47|504|-80.732725|64|35.082768|FRESH BERRIES|6.0|4|BLACKBERRIES 12 OZ|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00033383240015|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|2
35.082768|d821b7912b15a06401a1ffc2cb94f38b05e4bd2b|1.58|2014-10-31 15:11:00|80.732732175546019|1||147|35.099021295261316|0|35|532|-80.78468|64|35.096737|FRESH CUCUMBERS|0.0|4|COO CUCUMBERS S/S|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00204062000002|FRESH PRODUCE|PRODUCE|-80.732725|80.732726780676799|30|2
35.082768|0588c63be7de31246691750e2ade3fd081adaa79|2.67|2015-01-17 17:43:00|1.4091206135396188|1||147|0.6123098123133061|0|47|532|-80.732725|64|35.082768|FRESH CUCUMBERS|0.0|4|COO CUCUMBERS S/S|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00204062000002|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|3
35.082768|f10bfa22952bcfd79316d9082fbcd8953af12832|1.58|2015-03-01 17:35:00|1.4091206135396188|1||147|0.6123098123133061|0|47|532|-80.732725|64|35.082768|FRESH CUCUMBERS|0.0|4|COO CUCUMBERS S/S|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00204062000002|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|2
35.082768|4ec86a45dd00bd0e2a03a32b0a546afe45011d3b|1.58|2015-02-22 16:11:00|1.4091206135396188|1||147|0.6123098123133061|0|47|532|-80.732725|64|35.082768|FRESH CUCUMBERS|0.0|4|COO CUCUMBERS S/S|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00204062000002|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|2
35.082768|86d4dce50fbd4fd94e592a7123793a2388846909|2.37|2015-01-25 17:53:00|1.4091206135396188|1||147|0.6123098123133061|0|47|532|-80.732725|64|35.082768|FRESH CUCUMBERS|0.0|4|COO CUCUMBERS S/S|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00204062000002|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|3
35.082768|02df97a13a8d56cf67b58ddf0b0db1d038546fee|2.37|2014-12-07 15:23:00|1.4091206135396188|1||147|0.6123098123133061|0|47|532|-80.732725|64|35.082768|FRESH CUCUMBERS|0.0|4|COO CUCUMBERS S/S|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00204062000002|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|3
35.082768|3cb9808a526982b1e3918c1b3c9bcc580a4666b2|2.19|2014-12-12 08:27:00|1.4091206135396188|1|64420941200|147|0.6123098123133061|0|47|10|-80.732725|2|35.082768|LAYER CAKE MIX|0.94|1|D HINES FRENCH VANILLA CAKE|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00644209412808|BAKING MIXES|G1 GROCERY|-80.732725|1.409051865357139|147|1
35.082768|7f2da929c60d9106c45e6be4107f78747f0748c6|7.99|2014-11-05 17:27:00|1.4091206135396188|1|20639400000|147|0.6123098123133061|0|47|1654|-80.732725|381|35.082768|DESSERT CAKES|0.0|14|WHITE PATTI CAKE 2 LAYERS|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00206394000002|CAKES|BAKERY|-80.732725|1.409051865357139|147|1
35.082768|5c1a038b59658f6361a281846cec80a4936c6ce0|3.99|2015-02-17 19:44:00|1.4091206135396188|1|4114305160|147|0.6123098123133061|0|47|119|-80.732725|17|35.082768|RAISINS|0.0|1|SUN MAID GOLDEN RAISINS|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00041143051603|FRUIT-DRIED|G1 GROCERY|-80.732725|1.409051865357139|147|1
35.082768|ae33626ae723b681a6ae9190cbf02a709770e43c|11.25|2014-12-27 16:37:00|1.4091206135396188|1|4610000084|147|0.6123098123133061|0|47|318|-80.732725|52|35.082768|SHREDDED/GRATED CHEESE|0.0|3|SARGENTO REDUCED FAT MOZZ|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00046100000823|CHEESE|DAIRY|-80.732725|1.409051865357139|147|3
35.082768|abfae7061ae3cec9b4c7ebf6a2e46e2db1b6648b|7.3|2014-11-08 17:20:00|1.4091206135396188|1|4610000084|147|0.6123098123133061|0|47|318|-80.732725|52|35.082768|SHREDDED/GRATED CHEESE|2.3|3|SARGENTO REDUCED FAT MOZZ|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00046100000823|CHEESE|DAIRY|-80.732725|1.409051865357139|147|2
35.082768|bcfa32ab4871dc0bb4038f48d80ad25614ec24a6|7.9|2014-10-03 13:32:00|1.4091206135396188|1|4610000084|147|0.6123098123133061|0|47|318|-80.732725|52|35.082768|SHREDDED/GRATED CHEESE|1.98|3|SARGENTO REDUCED FAT MOZZ|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00046100000823|CHEESE|DAIRY|-80.732725|1.409051865357139|147|2
35.082768|ddd5d9d52b8b97e1a61ceeb9d1c96f6e7d823ee6|3.49|2014-10-17 14:18:00|1.4091206135396188|1|4610000084|147|0.6123098123133061|0|47|318|-80.732725|52|35.082768|SHREDDED/GRATED CHEESE|0.0|3|SARGENTO REDUCED FAT MOZZ|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00046100000823|CHEESE|DAIRY|-80.732725|1.409051865357139|147|1
35.082768|4f2cb4777d9404ce27d7d82a1a194f31943d352f|3.65|2014-11-14 14:53:00|1.4091206135396188|1|4610000084|147|0.6123098123133061|0|47|318|-80.732725|52|35.082768|SHREDDED/GRATED CHEESE|0.0|3|SARGENTO REDUCED FAT MOZZ|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00046100000823|CHEESE|DAIRY|-80.732725|1.409051865357139|147|1
35.082768|f8294f840f60645121b63fa16195f19ef42213eb|3.99|2014-10-20 20:33:00|1.4091206135396188|1|5210000647|147|0.6123098123133061|0|47|1245|-80.732725|34|35.082768|SINGLE SPICES|0.0|1|MC ONION POWDER|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00052100006475|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.732725|1.409051865357139|147|1
35.082768|57bccfe6397adb426176a63e0fd7ce273162158f|4.49|2015-02-01 12:00:00|1.4091206135396188|1|7203695649|147|0.6123098123133061|0|47|1699|-80.732725|387|35.082768|EVERYDAY (COOKIES)|0.0|14|HT YELLOW SOFT SUGAR COOKIES|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00072036956507|COOKIES|BAKERY|-80.732725|1.409051865357139|147|1
35.082768|b0974a8f9a17386ed8eb08b3b9103d95c9f7b3ec|4.49|2014-11-15 10:08:00|80.732732175546019|1|7203695649|147|35.099021285953221|0|35|1699|-80.810056|387|35.219587|EVERYDAY (COOKIES)|0.0|14|HT YELLOW SOFT SUGAR COOKIES|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00072036956507|COOKIES|BAKERY|-80.732725|80.732746333056937|401|1
35.082768|6d519323d9af87806ec67fd225ca456153ffadcb|1.29|2014-10-27 18:20:00|80.732732175546019|1|7203678692|147|35.099021295261316|0|35|1208|-80.78468|23|35.096737|WHSE PASTA VALUE ADD|0.0|1|HTO WW SPAGHETTI|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00072036786920|PASTA|G1 GROCERY|-80.732725|80.732726780676799|30|1
35.082768|a9234f828899b538f3836233bf0d119cd6987ade|0.97|2015-01-19 18:18:00|1.4091206135396188|1|7203688002|147|0.6123098123133061|0|47|527|-80.732725|64|35.082768|FRESH CARROTS|0.0|4|HT WHOLE CARROTS 2LB BAG|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00072036880024|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|1
35.082768|f9d3538171d0ec65f04c70fcc0a41560f0ab7143|0.97|2015-01-11 15:51:00|1.4091206135396188|1|7203688002|147|0.6123098123133061|0|47|527|-80.732725|64|35.082768|FRESH CARROTS|0.0|4|HT WHOLE CARROTS 2LB BAG|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00072036880024|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|1
35.082768|b93fae937f492efcbef818eac9c5ac2d461f9863|3.99|2015-01-07 18:08:00|1.4091206135396188|1|75166677005|147|0.6123098123133061|0|47|522|-80.732725|64|35.082768|FRESH TOMATOES|0.0|4|NATURESWEET CHERUBS 10.5 OZ|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00751666770058|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|1
35.082768|1d85e3cf9e4a8f2d2a0495396945e5490037415f|3.99|2014-12-23 17:41:00|1.4091206135396188|1|75166677005|147|0.6123098123133061|0|47|522|-80.732725|64|35.082768|FRESH TOMATOES|0.0|4|NATURESWEET CHERUBS 10.5 OZ|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00751666770058|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|1
35.082768|8dbab5215d590d4c80e8a81bd788c731b26a0f3f|3.99|2015-02-11 09:00:00|80.732732175546019|1|75166677005|147|35.099021295261316|0|35|522|-80.78468|64|35.096737|FRESH TOMATOES|0.0|4|NATURESWEET CHERUBS 10.5 OZ|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00751666770058|FRESH PRODUCE|PRODUCE|-80.732725|80.732726780676799|30|1
35.082768|1b1ecf5755dd9dc06d44d7632eda391e301864e5|3.99|2015-01-19 17:39:00|1.4091206135396188|1|75166677005|147|0.6123098123133061|0|47|522|-80.732725|64|35.082768|FRESH TOMATOES|0.0|4|NATURESWEET CHERUBS 10.5 OZ|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00751666770058|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|1
35.082768|321a6b36e19a445e78ef4d0b055ba06ab5845a8d|3.99|2015-02-07 18:12:00|1.4091206135396188|1|75166677005|147|0.6123098123133061|0|47|522|-80.732725|64|35.082768|FRESH TOMATOES|0.0|4|NATURESWEET CHERUBS 10.5 OZ|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00751666770058|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|1
35.082768|3538418f8ea4ceb348c18839ce34345954ef219f|3.99|2015-01-30 14:08:00|1.4091206135396188|1|75166677005|147|0.6123098123133061|0|47|522|-80.732725|64|35.082768|FRESH TOMATOES|0.0|4|NATURESWEET CHERUBS 10.5 OZ|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00751666770058|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|1
35.082768|d47deb00f2eb764994e10ea6f280fc70eeac204d|3.99|2014-09-22 15:07:00|1.4091206135396188|1|75166677005|147|0.6123098123133061|0|47|522|-80.732725|64|35.082768|FRESH TOMATOES|1.49|4|NATURESWEET CHERUBS 10.5 OZ|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00751666770058|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|1
35.082768|d9a62172f8b8041d64d40203d5cd2ea75db87e06|18.99|2014-12-06 15:39:00|80.732732175546019|1|7270010500|147|35.099021295261316|0|35|796|-80.78468|219|35.096737|KOSHER, DAILY USE-SPEC|3.0|1|MANISCH CHANUKAH DECO KIT|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00072700105002|SPECIALTY-ETHNIC FOODS|G1 GROCERY|-80.732725|80.732726780676799|30|1
35.082768|2fecc6c7e8eb21c59192e8d2e2f9cd6b8f454045|3.99|2015-01-15 21:03:00|1.4091206135396188|1|2791891223|147|0.6123098123133061|0|47|525|-80.732725|64|35.082768|FRESH LETTUCE|0.0|4|ARTISAN LETTUCE-CLAMSHELL|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00027918912232|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|1
35.082768|008a15653790a33fc9b5db214802cea802daab05|7.98|2014-09-12 17:59:00|1.4091206135396188|1|2791891223|147|0.6123098123133061|0|47|525|-80.732725|64|35.082768|FRESH LETTUCE|0.0|4|ARTISAN LETTUCE-CLAMSHELL|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00027918912232|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|2
35.082768|132b457cdfacb19e00d4535816706791ee28aea7|4.99|2014-11-12 18:04:00|80.732732175546019|1|2840003400|147|35.099021295261316|0|35|201|-80.78468|31|35.096737|POTATO CHIPS|1.0|1|RUFFLES ORIGINAL|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00028400034005|SNACKS|G1 GROCERY|-80.732725|80.732726780676799|30|1
35.082768|7a81d22d6c4169ba2483185a875c02da05939686|4.15|2014-11-17 18:07:00|80.732732175546019|1|4400000488|147|35.099021295261316|0|35|89|-80.78468|12|35.096737|GRAHAM CRACKERS|0.0|1|HONEYMAID GRAHAMS|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00044000004637|COOKIES|G1 GROCERY|-80.732725|80.732726780676799|30|1
35.082768|52d2742802921fd1da2ab5ce98acec3901b37479|5.39|2014-09-28 14:41:00|1.4091206135396188|1|5210007107|147|0.6123098123133061|0|47|217|-80.732725|34|35.082768|EXTRACTS FOOD COLORING|0.0|1|MC ASSORTED FOOD COLORS|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00052100071077|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.732725|1.409051865357139|147|1
35.082768|6289ba96e95d16acdc325fa18c74ac37e0259337|1.45|2015-01-24 16:54:00|1.4091206135396188|1||147|0.6123098123133061|0|47|502|-80.732725|64|35.082768|FRESH BANANAS|0.0|4|BANANAS, YELLOW|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00204011000008|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|1
35.082768|35337fc07da4b694ebb8c6de039aa3c003c4920a|4.99|2015-02-25 17:25:00|80.732732175546019|1|1111018700|147|35.099021291635339|0|35|1647|-80.80146|379|35.17739|PACKAGED MUFFINS|2.0|14|FFM 4 CT BLUEBERRY MUFFIN|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00011110187000|MUFFINS|BAKERY|-80.732725|80.732738387318278|208|1
35.082768|164b665b22e8e8c09963c587f689ca7d24b4ee57|4.69|2015-01-23 18:15:00|1.4091206135396188|1|81829001308|147|0.6123098123133061|0|47|685|-80.732725|61|35.082768|GREEK|0.0|3|CHOBANI 100 STRAWBERRY 4 PK|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00818290013071|YOGURT|DAIRY|-80.732725|1.409051865357139|147|1
35.082768|17e06a5989c972ac8c99e75d2e5e02f2229f6cfa|9.99|2015-02-20 14:30:00|1.4091206135396188|1|85768000101|147|0.6123098123133061|0|47|9960|-80.732725|887|35.082768|NFS-S/PREM-CAB SAUVIGNON|0.0|13|SHANNON RIDGE CABERNET SAUVIGN|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00857680001014|SUPER PREMIUM ($11-$14.99)|WINE|-80.732725|1.409051865357139|147|1
35.082768|f1efdb346248e2c9a0e4e39958698b10736fb114|1.5|2015-02-02 14:20:00|80.732732175546019|1||147|35.099021295261316|0|35|1617|-80.78468|373|35.096737|ROLLS BULK|0.0|14|BULK ROLLS|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00072036955555|ROLLS|BAKERY|-80.732725|80.732726780676799|30|2
35.082768|b60417f7b4b8f2b0d95e5182030daa0164f3935a|1.5|2014-12-03 09:07:00|80.732732175546019|1||147|35.099021295261316|0|35|1617|-80.78468|373|35.096737|ROLLS BULK|0.0|14|BULK ROLLS|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00072036955555|ROLLS|BAKERY|-80.732725|80.732726780676799|30|2
35.082768|70b25a017882d1777a626abf17f7338d636b740e|1.5|2014-09-17 18:33:00|1.4091206135396188|1||147|0.6123098123133061|0|47|1617|-80.732725|373|35.082768|ROLLS BULK|0.0|14|BULK ROLLS|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00072036955555|ROLLS|BAKERY|-80.732725|1.409051865357139|147|2
35.082768|80496c5491e9a4841ae5afd0a4e3c083cab907b3|14.669999999999998|2014-10-24 13:58:00|80.732732175546019|1|74236526435|147|35.099021295261316|0|35|345|-80.78468|57|35.096737|ORGANIC MILK|0.0|3|HORIZON ORGANIC FF DHA|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00742365003295|MILK|DAIRY|-80.732725|80.732726780676799|30|3
35.082768|d90a3031d033f3b5d5ce28d5f21a0645dd1128f0|10.12|2015-01-28 13:45:00|1.4091206135396188|1||147|0.6123098123133061|0|47|503|-80.732725|64|35.082768|FRESH GRAPES|1.45|4|RED GRAPES,SEEDLESS 12/16|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00204023000003|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|1
35.082768|4f03fee3239348a2de639161956bc4d66e609143|6.78|2014-09-27 18:54:00|1.4091206135396188|1|3800012158|147|0.6123098123133061|0|47|41|-80.732725|6|35.082768|BREAKFAST BARS|1.78|1|SPECIAL K BAR CHOC PRETZEL|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00038000466205|BREAKFAST FOODS|G1 GROCERY|-80.732725|1.409051865357139|147|2
35.082768|a14308e2f081fa0981a494f8888f6fe008571f84|10.98|2014-09-26 18:52:00|80.732732175546019|1|1410009589|147|35.099021295261316|0|35|1255|-80.78468|13|35.096737|LUNCH BOX CRACKERS|0.0|1|PP PF MULTIPACK GOLDFISH COLOR|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00014100096597|CRACKERS|G1 GROCERY|-80.732725|80.732726780676799|30|2
35.082768|cb68d8e34e46c8f5e1763596fa9d12714b3e4736|16.99|2015-02-14 18:56:00|1.4091206135396188|1|8500001163|147|0.6123098123133061|0|47|9972|-80.732725|888|35.082768|NFS-U/PREM-CAB SAUVIGNON|0.0|13|LOUIS MARTINI CAB SAUV SONOMA|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00085000011638|ULTRA PREMIUM ($15-$19.99)|WINE|-80.732725|1.409051865357139|147|1
35.082768|d33d1dd5bb8d544fe4a12dde9e64e06c1c5c1f34|9.99|2014-10-22 17:37:00|1.4091206135396188|1|7023666021|147|0.6123098123133061|0|47|751|-80.732725|87|35.082768|NFS-BOUQUETS|0.0|9|LOVE IN BLOOM|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00070236660217|FLORAL|FLORAL|-80.732725|1.409051865357139|147|1
35.082768|8df5f5d5648a7ab8c9ef613157f6baf3c8456f49|7.18|2014-12-02 18:11:00|1.4091206135396188|1||147|0.6123098123133061|0|47|500|-80.732725|64|35.082768|FRESH APPLES|0.0|4|CORTLAND APPLES|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00204106000005|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|1
35.082768|1f1d478f1fcfdce0a6910957f0b121da44045bc6|2.07|2014-10-04 11:14:00|1.4091206135396188|1||147|0.6123098123133061|0|47|500|-80.732725|64|35.082768|FRESH APPLES|0.0|4|CORTLAND APPLES|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00204106000005|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|1
35.082768|b8ba12971c3c3260b09617b652156aa4eb67bafd|2.78|2015-02-04 09:06:00|80.732732175546019|1|7675324990|147|35.099021295261316|0|35|5903|-80.78468|1538|35.096737|STRAWS|0.0|18|(JHK)(PPL) GDCK STRAWS JUMBO|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00076753249904|KITCHEN GADGETS|GM|-80.732725|80.732726780676799|30|2
35.082768|f52ff51c74f7fe779fbb02172b50b8520aef2dd7|8.98|2015-01-31 19:04:00|1.4091206135396188|1|70897191772|147|0.6123098123133061|0|47|1703|-80.732725|387|35.082768|SEASONAL COOKIES|2.0|14|VALENTINE PINK FRSTD SGR COOK|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00708971917722|COOKIES|BAKERY|-80.732725|1.409051865357139|147|2
35.082768|09e9e378459fb0cb7068b2c2def369d783add264|13.98|2014-10-09 18:02:00|1.4091206135396188|1|7203663045|147|0.6123098123133061|0|47|974|-80.732725|201|35.082768|FRESH TURKEY|2.0|2|HT 99% LEAN GRND TURKEY BREAST|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00072036630452|POULTRY|MEAT|-80.732725|1.409051865357139|147|2
35.082768|e34097cec2e193ca33c6c5956c7793228a81f727|3.99|2014-10-09 08:11:00|1.4091206135396188|1|4850002013|147|0.6123098123133061|0|47|335|-80.732725|56|35.082768|ORANGE JUICE-REGRIGERATED|0.99|3|TROPICANA PP ORIGINAL|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00048500301029|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.732725|1.409051865357139|147|1
35.082768|502b5ce4652b6d212a9eedfbf3197b942c3b2ee7|1.49|2014-10-17 13:29:00|80.732732175546019|1|1254600523|147|35.099021294357676|0|35|48|-80.771677|7|35.066546|REGISTER GUM|0.0|1|(FE)SOUR PATCH REDBERRY GUM|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00012546005234|CANDY|G1 GROCERY|-80.732725|80.732731858897139|45|1
35.082768|aa5cf56dd32db75e0f78e5f4f410a0df248c16a1|7.49|2014-09-28 14:52:00|1.4091206135396188|1|7675314987|147|0.6123098123133061|0|47|5879|-80.732725|1538|35.082768|FOOD PREPARATION|0.0|18|FUNNEL, CLPSBL|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00076753149877|KITCHEN GADGETS|GM|-80.732725|1.409051865357139|147|1
35.082768|e845327961ae71d9a8a00bbc5c1c9928ad3419fa|2.29|2014-10-10 19:13:00|1.4091206135396188|1|7203695739|147|0.6123098123133061|0|47|1976|-80.732725|475|35.082768|COLD PIZZA OTHER|0.0|6|WHITE PIZZA DOUGH BALLS|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00072036957399|PIZZA|DELI|-80.732725|1.409051865357139|147|1
35.082768|bf6c59729c139f585e51c18d0d9a6e8e9b71f392|7.98|2014-11-11 13:12:00|1.4091206135396188|1|20405400000|147|0.6123098123133061|0|47|504|-80.732725|64|35.082768|FRESH BERRIES|4.98|4|RED RASPBERRIES 6 OZ|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00715756100019|FRESH PRODUCE|PRODUCE|-80.732725|1.409051865357139|147|2
35.082768|75c38c8a4bfc4472571b67a68db7aa66889ccda7|4.99|2014-12-06 15:41:00|80.732732175546019|1|8817722767|147|35.099021295261316|0|35|79|-80.78468|273|35.096737|ASIAN SAUCES/SEASONINGS|0.0|1|SOY VAY ISLAND TERIYAKI|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00088177227642|ASIAN PREP. FOODS|G1 GROCERY|-80.732725|80.732726780676799|30|1
35.082768|53c36b5b62088ea596257eaccfa283d1774b4963|7.42|2014-10-10 18:54:00|80.732732175546019|1||147|35.099021295261316|0|35|503|-80.78468|64|35.096737|FRESH GRAPES|3.72|4|RED GRAPES,SEEDLESS 12/16|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00204023000003|FRESH PRODUCE|PRODUCE|-80.732725|80.732726780676799|30|1
35.082768|1d9695bc5550a76d43ead2232c5197f4bc53be0b|3.29|2014-09-25 19:08:00|80.732732175546019|1|1410008786|147|35.099021295261316|0|35|1034|-80.78468|163|35.096737|HOT DOG|0.3|7|PEP FRANKFURTER ROLLS PP|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|35.101032182271901|00014100070948|BUNS/ROLLS|COMMERCIAL BAKERY|-80.732725|80.732726780676799|30|1
35.082768|b4e45c0149e8520bbc44c70abe3a7c2d0e850d73|6.39|2014-11-24 21:50:00|1.4091206135396188|1|5150072001|147|0.6123098123133061|0|47|125|-80.732725|19|35.082768|PEANUT BUTTER|0.0|1|JIF CREAMY PEANUT BUTTER|faf99929d3673626b2b0fd5967bd524409556b57|1.1230634567663924|0.61242566243833529|00051500720011|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.732725|1.409051865357139|147|1
35.341927|640ba8b12561491ece7286abfae2f9909a9bf565|1.5|2015-01-16 11:03:00|80.780380710856576|4||220|35.367798795946413|0|48|1617|-80.66939|373|35.28326|ROLLS BULK|0.0|14|BULK ROLLS|fb9852d1cae58bd121b721d9e0aca9feae8e72e6|1.7876786498451105|35.351085445956379|00072036955555|ROLLS|BAKERY|-80.764523|80.764528624319681|46|2
35.341927|c77a1247f5f659855d4b211e455e4ffc00045eb0|4.79|2014-12-15 14:28:00|80.780380710856576|4|20165500000|220|35.367798795946413|0|48|297|-80.66939|49|35.28326|GROUND BEEF|0.0|2|HT PREMIUM GRND BEEF 80% LEAN|fb9852d1cae58bd121b721d9e0aca9feae8e72e6|1.7876786498451105|35.351085445956379|00201655000005|BEEF|MEAT|-80.764523|80.764528624319681|46|1
35.341927|72951bad98c843440515006be9db2e8467bc42a1|1.61|2014-09-26 16:51:00|80.780380710856576|4||220|35.367798795946413|0|48|505|-80.66939|64|35.28326|FRESH SOFT FRUIT|0.27|4|BLACK PLUMS|fb9852d1cae58bd121b721d9e0aca9feae8e72e6|1.7876786498451105|35.351085445956379|00204040000000|FRESH PRODUCE|PRODUCE|-80.764523|80.764528624319681|46|1
35.341927|e4717525bcb38ae6b429aeabe24670d2893cd17b|2.19|2014-11-26 14:55:00|80.780380710856576|4|1200000230|220|35.367798795946413|0|48|55|-80.66939|8|35.28326|REGULAR|0.94|23|SIERRA MIST NATURAL 2 LITER|fb9852d1cae58bd121b721d9e0aca9feae8e72e6|1.7876786498451105|35.351085445956379|00012000158056|CARBONATED BEVERAGES|BEVERAGE|-80.764523|80.764528624319681|46|1
35.341927|8800b59ab7bb4d49d8436543e41ceb742abde6b4|2.19|2015-01-06 14:52:00|80.780380710856576|4|1200000230|220|35.367798795946413|0|48|55|-80.66939|8|35.28326|REGULAR|0.94|23|SIERRA MIST NATURAL 2 LITER|fb9852d1cae58bd121b721d9e0aca9feae8e72e6|1.7876786498451105|35.351085445956379|00012000158056|CARBONATED BEVERAGES|BEVERAGE|-80.764523|80.764528624319681|46|1
35.341927|8ef96c35810e7f0217c555e8d2ce3707420540a6|8.34|2014-09-24 15:07:00|80.780380710856576|4||220|35.367798795946413|0|48|542|-80.66939|64|35.28326|FRESH VEGETABLES REMAIN|0.0|4|COO RHUBARB|fb9852d1cae58bd121b721d9e0aca9feae8e72e6|1.7876786498451105|35.351085445956379|00204745000008|FRESH PRODUCE|PRODUCE|-80.764523|80.764528624319681|46|1
35.341927|23bb292bea63566e12b687f4bda719bb2d83457e|3.85|2014-12-01 15:20:00|80.780380710856576|4|2100060464|220|35.367798795946413|0|48|315|-80.66939|52|35.28326|CHEESE-PROCESSED-SLICED|0.0|3|KRAFT WHITE AMERICAN|fb9852d1cae58bd121b721d9e0aca9feae8e72e6|1.7876786498451105|35.351085445956379|00021000604654|CHEESE|DAIRY|-80.764523|80.764528624319681|46|1
35.372142|1619a65c19f37d5cc79def26805eeca6c6e62a30|4.99|2015-02-06 14:40:00|80.779636304526477|3|1111018700|122|35.407683132507167|0|17|1647|-80.814133|379|35.333742|PACKAGED MUFFINS|2.5|14|FFM 4 CT LEMON POPPY MUFFIN|fc1c2b38011658417d4b6b4e8592ef5fadf4e629|2.4558067871319182|35.392509581117899|00011110187048|MUFFINS|BAKERY|-80.782849|80.7828725943764|472|1
35.372142|cfa5583f084c35e5d082080d999bf4dd6221ef81|4.99|2015-01-08 10:50:00|80.779636304526477|3|1111018700|122|35.407683132507167|0|17|1647|-80.814133|379|35.333742|PACKAGED MUFFINS|2.5|14|FFM 4 CT LEMON POPPY MUFFIN|fc1c2b38011658417d4b6b4e8592ef5fadf4e629|2.4558067871319182|35.392509581117899|00011110187048|MUFFINS|BAKERY|-80.782849|80.7828725943764|472|1
35.372142|9eb97f0e8a2fc0ce13832832b7141cf9dbe4a3ef|3.99|2014-11-04 13:13:00|80.779636304526477|3|1906301228|122|35.407683132507167|0|17|31|-80.814133|4|35.333742|NON CARBONATED WATER|1.0|1|VYFINE FRUIT 2 O NAT STRW 6PK|fc1c2b38011658417d4b6b4e8592ef5fadf4e629|2.4558067871319182|35.392509581117899|00019063232341|BOTTLED WATER|G1 GROCERY|-80.782849|80.7828725943764|472|1
35.372142|039194530830cb8b038b1e85e886ae2bffb62645|3.99|2014-11-12 18:46:00|80.779636304526477|3|1906301228|122|35.407683132507167|0|17|31|-80.814133|4|35.333742|NON CARBONATED WATER|0.49|1|VYFINE FRUIT 2 O NAT STRW 6PK|fc1c2b38011658417d4b6b4e8592ef5fadf4e629|2.4558067871319182|35.392509581117899|00019063232341|BOTTLED WATER|G1 GROCERY|-80.782849|80.7828725943764|472|1
35.372142|bc19379b66cc9e2c5f1d8b501afb5887293aeec8|3.99|2014-09-19 10:34:00|80.779636304526477|3|1906301228|122|35.407683132507167|0|17|31|-80.814133|4|35.333742|NON CARBONATED WATER|2.0|1|VYFINE FRUIT 2 O NAT STRW 6PK|fc1c2b38011658417d4b6b4e8592ef5fadf4e629|2.4558067871319182|35.392509581117899|00019063232341|BOTTLED WATER|G1 GROCERY|-80.782849|80.7828725943764|472|1
35.372142|bc9fa5d6c281defa84a3d618a9c7e965931748b7|7.98|2015-03-02 16:56:00|80.779636304526477|3|1906301228|122|35.407683132507167|0|17|31|-80.814133|4|35.333742|NON CARBONATED WATER|1.99|1|VYFINE FRUIT 2 O NAT STRW 6PK|fc1c2b38011658417d4b6b4e8592ef5fadf4e629|2.4558067871319182|35.392509581117899|00019063232341|BOTTLED WATER|G1 GROCERY|-80.782849|80.7828725943764|472|2
35.372142|fb192604c1b3a0ec4ef0ba6054214df596202e53|3.99|2015-02-01 17:19:00|80.779636304526477|3|1906301228|122|35.407683132507167|0|17|31|-80.814133|4|35.333742|NON CARBONATED WATER|1.0|1|VYFINE FRUIT 2 O NAT STRW 6PK|fc1c2b38011658417d4b6b4e8592ef5fadf4e629|2.4558067871319182|35.392509581117899|00019063232341|BOTTLED WATER|G1 GROCERY|-80.782849|80.7828725943764|472|1
35.372142|13098b5ff535604ccf75182d02a20f5868312887|2.58|2014-11-25 11:54:00|80.779636304526477|3|5100002524|122|35.407683136766913|0|17|179|-80.764523|27|35.341927|CANNED PASTA|0.58|1|SPAGHETTIOS PLUS CALCIUM|fc1c2b38011658417d4b6b4e8592ef5fadf4e629|2.4558067871319182|35.392509581117899|00051000138194|PREPARED FOODS-RTS|G1 GROCERY|-80.782849|80.78285905456417|220|2
35.372142|d865d7ffb34bb1db73213b3bdb8549fa50492a55|3.99|2014-10-01 15:10:00|80.779636304526477|3|4650072048|122|35.40768313246425|0|17|393|-80.780702|68|35.318911|NFS-AIR FRESHENERS|0.0|1|GLADE DECOR GLASS LINEN|fc1c2b38011658417d4b6b4e8592ef5fadf4e629|2.4558067871319182|35.392509581117899|00046500720482|FRESHENERS/DEODORIZERS|G1 GROCERY|-80.782849|80.782872691456504|167|1
35.372142|85a137531a0064ff189ddc39437218e668b117f2|6.79|2015-03-06 11:11:00|80.779636304526477|3|30085075605|122|35.40768313246425|0|17|4243|-80.780702|1200|35.318911|NASAL PRODUCT-ADULT|1.8|17|AFRIN NASAL SPRAY 15ML-75605|fc1c2b38011658417d4b6b4e8592ef5fadf4e629|2.4558067871319182|35.392509581117899|00300850756059|COUGH/COLD/SINUS|HBC|-80.782849|80.782872691456504|167|1
35.372142|f22009868c24a824a27ddd242c6b63ffedcfe8cd|1.2|2014-12-22 18:54:00|80.779636304526477|3|7047000100|122|35.407683132507167|0|17|687|-80.814133|61|35.333742|BLENDED|0.0|3|YOPLAIT VANILLA CUSTARD|fc1c2b38011658417d4b6b4e8592ef5fadf4e629|2.4558067871319182|35.392509581117899|00070470001128|YOGURT|DAIRY|-80.782849|80.7828725943764|472|2
35.372142|b63238bfc35ef36d7c93976c6bdcda1153d8e036|2.4|2014-10-24 12:19:00|80.779636304526477|3|7047000100|122|35.407683132507167|0|17|687|-80.814133|61|35.333742|BLENDED|0.0|3|YOPLAIT VANILLA CUSTARD|fc1c2b38011658417d4b6b4e8592ef5fadf4e629|2.4558067871319182|35.392509581117899|00070470001128|YOGURT|DAIRY|-80.782849|80.7828725943764|472|4
35.372142|db9ace19750a58444903572ad6a7c88c3d03b5e8|2.79|2015-02-20 15:50:00|80.779636304526477|3|4300004209|122|35.407683132507167|0|17|343|-80.814133|59|35.333742|PUDDINGS|0.79|3|JELL-O SF VANILLA|fc1c2b38011658417d4b6b4e8592ef5fadf4e629|2.4558067871319182|35.392509581117899|00043000042007|SNACKS/SPREADS/DIPS-DAIRY|DAIRY|-80.782849|80.7828725943764|472|1
35.372142|b9e16c40cb7dd33dbdfc966850774bf61bbcd45c|4.99|2014-11-19 17:43:00|80.779636304526477|3|1111018700|122|35.407683132507167|0|17|1647|-80.814133|379|35.333742|PACKAGED MUFFINS|1.02|14|FFM 4 CT BLUEBERRY MUFFIN|fc1c2b38011658417d4b6b4e8592ef5fadf4e629|2.4558067871319182|35.392509581117899|00011110187000|MUFFINS|BAKERY|-80.782849|80.7828725943764|472|1
35.372142|26900a83d128d4f3128380dd1d264cc2ded932da|3.25|2014-12-12 13:56:00|80.779636304526477|3|7203656080|122|35.407683132507167|0|17|318|-80.814133|52|35.333742|SHREDDED/GRATED CHEESE|0.0|3|HT FANCY SHRED SHARP CHED CHE|fc1c2b38011658417d4b6b4e8592ef5fadf4e629|2.4558067871319182|35.392509581117899|00072036550262|CHEESE|DAIRY|-80.782849|80.7828725943764|472|1
35.372142|83794a97c8e9449650e474243c79224be75d7996|4.69|2015-01-22 14:01:00|80.779636304526477|3|5200050632|122|35.407683132507167|0|17|30|-80.814133|4|35.333742|CARBONATED WATER|2.34|1|PROPEL BERRY 6PK|fc1c2b38011658417d4b6b4e8592ef5fadf4e629|2.4558067871319182|35.392509581117899|00052000506334|BOTTLED WATER|G1 GROCERY|-80.782849|80.7828725943764|472|1
35.372142|960072b14f3ef225d811beff7a874839b4d4efc1|5.79|2015-01-14 16:24:00|80.779636304526477|3|7203001108|122|35.407683132507167|0|17|1685|-80.814133|385|35.333742|ENTENMANNS (SWEET GOODS)|0.0|14|ENT SOFTEE VARIETY DNTS PP|fc1c2b38011658417d4b6b4e8592ef5fadf4e629|2.4558067871319182|35.392509581117899|00072030011080|SWEET GOODS|BAKERY|-80.782849|80.7828725943764|472|1
35.372142|e65c6ec2689a1d8c3c0b3d3832138b31b647cb65|2.75|2014-12-24 11:41:00|80.779636304526477|3|5150025537|122|35.407683132507167|0|17|125|-80.814133|19|35.333742|PEANUT BUTTER|0.0|1|JIF CREAMY PEANUT BUTTER|fc1c2b38011658417d4b6b4e8592ef5fadf4e629|2.4558067871319182|35.392509581117899|00051500255162|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.782849|80.7828725943764|472|1
35.43259|d538b0af9fe5e8cbfcdd6a80edcdb99e80136f49|7.99|2014-11-20 14:40:00|1.4057311447477159|4|3338314604|202|0.6184153580092175|0|52|509|-80.605588|64|35.43259|FRESH CITRUS-REMAINING|3.0|4|CLEMENTINES 5LB BOX|fee19bda19cf63d8dbe351e6d7a10e974101f2da|10.434887448795624|0.6209993146566879|00033383146041|FRESH PRODUCE|PRODUCE|-80.605588|1.406832906106031|202|1
35.066546|d4e74434e5fa8a80c835651d958a05a045e8b00c|3.99|2015-01-31 14:20:00|1.4091206135396188|1|9220900152|45|0.6120266850020475|0|47|559|-80.771677|64|35.066546|SPECIALTY-DRIED FRUIT & VEG.|0.0|4|DRIED NUTRA FIGS   9 OZ|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00097209001525|FRESH PRODUCE|PRODUCE|-80.771677|1.409731706007376|45|1
35.066546|5d8e51e012ba930b7fba456ab61539614d1fdb9f|9.99|2014-09-13 14:31:00|80.782094729586973|1|8500001222|45|35.085677203710837|0|27|9939|-80.770346|885|35.052812|NFS POP PINOT NOIR|0.0|13|REDWOOD CREEK PINOT NOIR 1.5L|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00085000012222|POPULAR (4-$7.99)|WINE|-80.771677|80.771680204378441|40|1
35.066546|3e11945c15bc99116ca7209385172b0eb3a70d65|9.99|2014-11-30 14:52:00|1.4091206135396188|1|8500001688|45|0.6120266850020475|0|47|9941|-80.771677|885|35.066546|NFS POP ZINFANDEL|0.0|13|REDWOOD CREEK RED MOSCATO 1.5L|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00085000016886|POPULAR (4-$7.99)|WINE|-80.771677|1.409731706007376|45|1
35.066546|af41b2f53934adcab0b66956222beade3cd02b5b|3.49|2014-11-10 17:45:00|80.782094729586973|1|8087800218|45|35.085677203265348|0|27|3536|-80.78468|1045|35.096737|SHAMPOO-PREMIUM|0.0|17|PANTENE SH FINE FLAT/VOLUME|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00080878042166|HAIR & SCALP CARE|HBC|-80.771677|80.771682976423307|30|1
35.066546|1b9462acab525ce82b0ff6e2945ed0c41f67891e|8.58|2014-09-21 13:49:00|1.4091206135396188|1|7341000305|45|0.6120266850020475|0|47|1026|-80.771677|162|35.066546|WHEAT|2.15|7|ARN CNTRY OATMEAL BREAD WP PP|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00073410003558|SLICED BREAD|COMMERCIAL BAKERY|-80.771677|1.409731706007376|45|2
35.066546|f40007b0cefd3db4f38779fa411f315e99ecc83c|2.99|2014-12-10 17:02:00|80.782094729586973|1|2484201121|45|35.085677203265348|0|27|1887|-80.78468|440|35.096737|PASTA CUTS|0.0|6|BUITONI FETTUCINE|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00024842011215|PASTA|DELI|-80.771677|80.771682976423307|30|1
35.066546|1ba839680c78ebc2389b7cea75f36578d6f77a1a|3.99|2014-12-20 13:21:00|1.4091206135396188|1|2791891223|45|0.6120266850020475|0|47|525|-80.771677|64|35.066546|FRESH LETTUCE|0.0|4|ARTISAN LETTUCE-CLAMSHELL|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00027918912232|FRESH PRODUCE|PRODUCE|-80.771677|1.409731706007376|45|1
35.066546|c352e246f0923343d52126da014b4e4d3e347181|2.99|2014-10-22 16:41:00|80.782094729586973|1|2484201151|45|35.085677203265348|0|27|1887|-80.78468|440|35.096737|PASTA CUTS|0.0|6|BUITONI ANGEL HAIR|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00024842011512|PASTA|DELI|-80.771677|80.771682976423307|30|1
35.066546|0af8810f2e174183b4014c30daf8eba60436d178|3.29|2015-01-29 17:38:00|80.782094729586973|1|2484201151|45|35.085677203265348|0|27|1887|-80.78468|440|35.096737|PASTA CUTS|0.0|6|BUITONI ANGEL HAIR|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00024842011512|PASTA|DELI|-80.771677|80.771682976423307|30|1
35.066546|84af90ef8e560840725a7a76baaf57183c224b53|2.99|2014-12-22 17:17:00|80.782094729586973|1|20424200000|45|35.085677203265348|0|27|512|-80.78468|64|35.096737|FRSH PROD FRSH FRUIT REM|0.99|4|CRANBERRIES 12 OZ|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00031200900043|FRESH PRODUCE|PRODUCE|-80.771677|80.771682976423307|30|1
35.066546|02fbf2a1687b0d0670148d547418cd13cf4243f4|7.99|2015-02-08 13:32:00|1.4091206135396188|1|2840000288|45|0.6120266850020475|0|47|205|-80.771677|31|35.066546|REMAINING SNACKS|1.0|1|SUNCHIPS & ROLD GOLD MIX|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00028400264983|SNACKS|G1 GROCERY|-80.771677|1.409731706007376|45|1
35.066546|42bb828e032aecef9c1b6600da90ae7e1b6687b1|1.99|2015-01-17 11:28:00|80.782094729586973|1|7203688096|45|35.085677196303678|0|27|526|-80.709466|64|35.124987|FRESH MUSHROOMS|0.2|4|HT SLICED WHITE MUSHROOMS|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00072036880963|FRESH PRODUCE|PRODUCE|-80.771677|80.771697818915101|157|1
35.066546|d8aa2918993ccf71792a98d934c0182f6c5ab03c|3.98|2015-02-28 14:23:00|1.4091206135396188|1|7203688096|45|0.6120266850020475|0|47|526|-80.771677|64|35.066546|FRESH MUSHROOMS|0.4|4|HT SLICED WHITE MUSHROOMS|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00072036880963|FRESH PRODUCE|PRODUCE|-80.771677|1.409731706007376|45|2
35.066546|34ce882382339ea8f250a6c73014a45331cf6310|1.99|2015-02-18 15:10:00|80.782094729586973|1|7203688096|45|35.085677203265348|0|27|526|-80.78468|64|35.096737|FRESH MUSHROOMS|0.0|4|HT SLICED WHITE MUSHROOMS|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00072036880963|FRESH PRODUCE|PRODUCE|-80.771677|80.771682976423307|30|1
35.066546|ff25e86afd494d48f6aa762f164563a11c4bb3c8|1.99|2015-01-11 13:22:00|1.4091206135396188|1|7203688096|45|0.6120266850020475|0|47|526|-80.771677|64|35.066546|FRESH MUSHROOMS|0.1|4|HT SLICED WHITE MUSHROOMS|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00072036880963|FRESH PRODUCE|PRODUCE|-80.771677|1.409731706007376|45|1
35.066546|2bde46f092579507fc50038a5cd1987a5df5fdc6|1.99|2014-12-07 12:03:00|1.4091206135396188|1|7203688096|45|0.6120266850020475|0|47|526|-80.771677|64|35.066546|FRESH MUSHROOMS|0.2|4|HT SLICED WHITE MUSHROOMS|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00072036880963|FRESH PRODUCE|PRODUCE|-80.771677|1.409731706007376|45|1
35.066546|4b1ee7ac26673d4a4037603cde229b0096cce384|1.99|2014-12-29 14:09:00|1.4091206135396188|1|7203688096|45|0.6120266850020475|0|47|526|-80.771677|64|35.066546|FRESH MUSHROOMS|0.0|4|HT SLICED WHITE MUSHROOMS|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00072036880963|FRESH PRODUCE|PRODUCE|-80.771677|1.409731706007376|45|1
35.066546|669a2ecffdd51bbb303d9034a3d264c11f91ddc0|1.99|2015-02-02 17:09:00|1.4091206135396188|1|7203688096|45|0.6120266850020475|0|47|526|-80.771677|64|35.066546|FRESH MUSHROOMS|0.2|4|HT SLICED WHITE MUSHROOMS|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00072036880963|FRESH PRODUCE|PRODUCE|-80.771677|1.409731706007376|45|1
35.066546|a7c38476f37a814dc17894aba688869ccc4763bc|1.99|2015-01-03 14:56:00|1.4091206135396188|1|7203688096|45|0.6120266850020475|0|47|526|-80.771677|64|35.066546|FRESH MUSHROOMS|0.0|4|HT SLICED WHITE MUSHROOMS|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00072036880963|FRESH PRODUCE|PRODUCE|-80.771677|1.409731706007376|45|1
35.066546|4302c2a7a4617f3b9c228ee250dc52d0991f22f8|1.99|2015-02-04 17:39:00|80.782094729586973|1|7203688096|45|35.085677203265348|0|27|526|-80.78468|64|35.096737|FRESH MUSHROOMS|0.0|4|HT SLICED WHITE MUSHROOMS|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00072036880963|FRESH PRODUCE|PRODUCE|-80.771677|80.771682976423307|30|1
35.066546|83c5608e2b8b938bc8e21c486d5da24ae4c84264|2.99|2014-10-03 18:04:00|80.782094729586973|1|89602800100|45|35.085677203265348|0|27|544|-80.78468|64|35.096737|FRESH PRODUCE FRSH HERBS|0.0|4|HYDROPONIC LIVING BASIL|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00895148002111|FRESH PRODUCE|PRODUCE|-80.771677|80.771682976423307|30|1
35.066546|786131002cdea309442a71d45262f926f6c7d669|3.29|2014-12-03 17:17:00|80.782094729586973|1|1410008786|45|35.085677203265348|0|27|1033|-80.78468|163|35.096737|HAMBURGER|0.0|7|PEP  WHEAT HAMBURGER BUNS PP|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00014100087861|BUNS/ROLLS|COMMERCIAL BAKERY|-80.771677|80.771682976423307|30|1
35.066546|3554e09c6e5c43833ffe23442149e8c5236cd2f4|29.58|2015-01-26 17:13:00|80.782094729586973|1|76211177857|45|35.085677203265348|0|27|36|-80.78468|10|35.096737|PREMIUM GROUND|5.6|1|STARBUCKS GRND BRKFST BLEND|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00762111778574|COFFEE|G1 GROCERY|-80.771677|80.771682976423307|30|2
35.066546|569d1505849689b5444f6fe43033d6fc187fa85d|2.99|2015-01-07 17:17:00|1.4091206135396188|1|3338365583|45|0.6120266850020475|0|47|522|-80.771677|64|35.066546|FRESH TOMATOES|0.2|4|SWEET GRAPE TOMATO (PINT)|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00814369011214|FRESH PRODUCE|PRODUCE|-80.771677|1.409731706007376|45|1
35.066546|ac59cee279425c01dc2ff4df324dfc3c7bf8bedc|2.99|2014-12-14 17:08:00|1.4091206135396188|1|3338365583|45|0.6120266850020475|0|47|522|-80.771677|64|35.066546|FRESH TOMATOES|0.49|4|SWEET GRAPE TOMATO (PINT)|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00814369011214|FRESH PRODUCE|PRODUCE|-80.771677|1.409731706007376|45|1
35.066546|eae6ad43f8ea5774d9d0615977993e9109cc39da|14.79|2015-02-23 16:35:00|80.782094729586973|1|76211177857|45|35.085677203265348|0|27|36|-80.78468|10|35.096737|PREMIUM GROUND|1.8|1|STARBUCKS GRND BRKFST BLEND|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00762111778574|COFFEE|G1 GROCERY|-80.771677|80.771682976423307|30|1
35.066546|c050a95fb9cf6a038a0fdf30ee592de9e7c39e96|14.79|2014-09-25 18:55:00|1.4091206135396188|1|76211177857|45|0.6120266850020475|0|47|36|-80.771677|10|35.066546|PREMIUM GROUND|0.0|1|STARBUCKS GRND BRKFST BLEND|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00762111778574|COFFEE|G1 GROCERY|-80.771677|1.409731706007376|45|1
35.066546|f9ef938c243c0946ec71ec2fd24b3ef627d39e64|14.79|2014-12-31 14:32:00|1.4091206135396188|1|76211177857|45|0.6120266850020475|0|47|36|-80.771677|10|35.066546|PREMIUM GROUND|0.0|1|STARBUCKS GRND BRKFST BLEND|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00762111778574|COFFEE|G1 GROCERY|-80.771677|1.409731706007376|45|1
35.066546|47554a9bd2cc52f8fd85a045fae8f2c78cbf44c8|14.79|2014-10-09 16:46:00|80.782094729586973|1|76211177857|45|35.085677203265348|0|27|36|-80.78468|10|35.096737|PREMIUM GROUND|0.0|1|STARBUCKS GRND BRKFST BLEND|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00762111778574|COFFEE|G1 GROCERY|-80.771677|80.771682976423307|30|1
35.066546|993c37681a31823424308cdcf1d5ca75e7f2b6e1|14.79|2014-10-26 14:41:00|1.4091206135396188|1|76211177857|45|0.6120266850020475|0|47|36|-80.771677|10|35.066546|PREMIUM GROUND|0.0|1|STARBUCKS GRND BRKFST BLEND|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00762111778574|COFFEE|G1 GROCERY|-80.771677|1.409731706007376|45|1
35.066546|484c61bc18da2c5edcad84a3d5d936e94daa2918|14.79|2015-02-13 17:15:00|1.4091206135396188|1|76211177857|45|0.6120266850020475|0|47|36|-80.771677|10|35.066546|PREMIUM GROUND|0.0|1|STARBUCKS GRND BRKFST BLEND|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00762111778574|COFFEE|G1 GROCERY|-80.771677|1.409731706007376|45|1
35.066546|ba97c6cbf462ba7eb8ae68005a9a55f1693e6cb2|2.99|2014-11-22 17:38:00|1.4091206135396188|1|3338365583|45|0.6120266850020475|0|47|522|-80.771677|64|35.066546|FRESH TOMATOES|0.2|4|SWEET GRAPE TOMATO (PINT)|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00814369011214|FRESH PRODUCE|PRODUCE|-80.771677|1.409731706007376|45|1
35.066546|b2495b6155c40e58c281da54f0c1a785ad5d93be|12.78|2014-12-13 11:07:00|1.4091206135396188|1|4154800385|45|0.6120266850020475|0|47|252|-80.771677|45|35.066546|PREMIUM ICE CREAM|6.4|5|EDY'S LIGHT VANILLA BEAN|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00041548003863|ICE CREAM|FROZEN|-80.771677|1.409731706007376|45|2
35.066546|206e4ba4fb3c93f48c7febe86a0a2b9df21c3218|6.39|2014-10-13 17:14:00|80.782094729586973|1|4154800385|45|35.085677203265348|0|27|252|-80.78468|45|35.096737|PREMIUM ICE CREAM|1.61|5|EDY'S SLOW CHURNED CARAMEL D|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00041548345864|ICE CREAM|FROZEN|-80.771677|80.771682976423307|30|1
35.066546|f396f78f02c206fde5c513d71d5e04543cdc3677|1.39|2014-12-23 14:53:00|1.4091206135396188|1|3710003578|45|0.6120266850020475|0|47|245|-80.771677|39|35.066546|VEGETABLES-CORE|0.2|1|LIBBY GRN BEANS CUT|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00037100033188|VEGETABLES-CAN/JAR|G1 GROCERY|-80.771677|1.409731706007376|45|1
35.066546|156ced756ba3e16b64aa8208927389c0a6fe25f5|2.79|2015-01-08 16:58:00|80.782094729586973|1|3800035900|45|35.085677203710837|0|27|41|-80.770346|6|35.052812|BREAKFAST BARS|0.29|1|KLGS NUTRI GRN BAR BLUEBERRY|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00038000357008|BREAKFAST FOODS|G1 GROCERY|-80.771677|80.771680204378441|40|1
35.066546|098dba45e9bb02f7fa5c649bdc36d98c394bf2ce|2.58|2015-01-20 17:07:00|1.4091206135396188|1|3940001810|45|0.6120266850020475|0|47|242|-80.771677|39|35.066546|CANNED BEANS|0.58|1|BUSH PEAS BLACKEYE|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00039400013686|VEGETABLES-CAN/JAR|G1 GROCERY|-80.771677|1.409731706007376|45|2
35.066546|d0a1f3f91a534de72d4158c8dfe8f8098b9d1cfb|3.59|2014-10-18 16:38:00|1.4091206135396188|1|3700007100|45|0.6120266850020475|0|47|393|-80.771677|68|35.066546|NFS-AIR FRESHENERS|0.6|1|FEBREZE AIR AFFECTS LINEN SKY|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00037000071006|FRESHENERS/DEODORIZERS|G1 GROCERY|-80.771677|1.409731706007376|45|1
35.066546|70d3b71257e510bcfa75f1dec6483849e6c4d78f|3.99|2015-02-16 13:45:00|1.4091206135396188|1|4129497325|45|0.6120266850020475|0|47|400|-80.771677|69|35.066546|NFS-LIQUID CLEANERS|0.0|1|PINE SOL LIQUID 40 OZ|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00041294973250|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.771677|1.409731706007376|45|1
35.066546|79795920855bc5c268abdd88b95ec18697c421f0|2.99|2015-03-03 16:39:00|80.782094729586973|1|3338365583|45|35.085677203265348|0|27|522|-80.78468|64|35.096737|FRESH TOMATOES|0.49|4|SWEET GRAPE TOMATO (PINT)|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00072036880284|FRESH PRODUCE|PRODUCE|-80.771677|80.771682976423307|30|1
35.066546|dd256400112f4acee4c87495a0f19fa5570a1a5c|4.98|2015-03-07 15:33:00|1.4091206135396188|1|7203688048|45|0.6120266850020475|0|47|526|-80.771677|64|35.066546|FRESH MUSHROOMS|0.98|4|HT SLICED BABY BELLAS|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00072036880482|FRESH PRODUCE|PRODUCE|-80.771677|1.409731706007376|45|2
35.066546|467900370b98ceee9ff4e7e68aa52cb2ef9e6ca7|3.99|2014-09-18 18:13:00|80.782094729586973|1|3400007610|45|35.085677203265348|0|27|727|-80.78468|7|35.096737|SEASONAL CANDY-SINGLE FAC|0.4|1|I/O(H15)KIT KAT HARVEST BAG|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00034000076109|CANDY|G1 GROCERY|-80.771677|80.771682976423307|30|1
35.066546|5190a532e0f86dfb993c11f8c3f62ca88cfc3ec1|3.39|2015-02-10 16:37:00|1.4091206135396188|1|5260305445|45|0.6120266850020475|0|47|214|-80.771677|33|35.066546|BROTH|0.0|1|PACIFIC ORG LS BEEF BROTH|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00052603054362|SOUP|G1 GROCERY|-80.771677|1.409731706007376|45|1
35.066546|474c11ad3c0b6afb1091b2791fb537341a54d226|2.38|2014-11-03 17:28:00|1.4091206135396188|1|7203600022|45|0.6120266850020475|0|47|6859|-80.771677|1581|35.066546|RE USEABLE EVERYDAY|0.4|18|HT REUSABLE GREEN TOTE|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00072036000224|SHOPPING BAGS|GM|-80.771677|1.409731706007376|45|2
35.066546|4061d2d8890e6a7c6b67fcb728af2c16115380ff|1.69|2015-02-25 16:50:00|80.782094729586973|1|7090050126|45|35.085677203265348|0|27|1221|-80.78468|275|35.096737|PASTA SC VALUE|0.0|1|DEI FRTLI PIZZA SAUCE|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00070900501266|PASTA SAUCES|G1 GROCERY|-80.771677|80.771682976423307|30|1
35.066546|8827937078d67fc2b2d3dec9294bf1f8e42c9bf1|4.99|2014-12-06 16:14:00|80.782094729586973|1|7144830025|45|35.085677203265348|0|27|2021|-80.78468|505|35.096737|FRESH CHEESE|0.0|6|ALOUETTE SPINACH & ARTICHOKE|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00071448300199|SPECIALTY CHEESE|DELI|-80.771677|80.771682976423307|30|1
35.066546|16d7751c0fc672b70c4d52558e6916257566e709|1.19|2014-11-14 16:43:00|80.782094729586973|1|7203600022|45|35.085677203265348|0|27|6859|-80.78468|1581|35.096737|RE USEABLE EVERYDAY|0.2|18|HT REUSABLE GREEN TOTE|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00072036000224|SHOPPING BAGS|GM|-80.771677|80.771682976423307|30|1
35.066546|a5f6298becb03782f4456e35d787b48efd3bcc9b|4.99|2015-01-13 17:19:00|80.782094729586973|1|7144830025|45|35.085677203265348|0|27|2021|-80.78468|505|35.096737|FRESH CHEESE|0.0|6|ALOUETTE SPINACH & ARTICHOKE|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00071448300199|SPECIALTY CHEESE|DELI|-80.771677|80.771682976423307|30|1
35.066546|3753984edcba01050886bc2bce3d187f8ef1cee6|1.59|2014-09-10 17:41:00|80.782094729586973|1|7090050126|45|35.085677203265348|0|27|1221|-80.78468|275|35.096737|PASTA SC VALUE|0.0|1|DEI FRTLI PIZZA SAUCE|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00070900501266|PASTA SAUCES|G1 GROCERY|-80.771677|80.771682976423307|30|1
35.066546|6f07d297c4215e74cff5d92ac341c5f6c0f7e0a1|9.99|2014-10-11 10:58:00|80.782094729586973|1|8500001870|45|35.085677203710837|0|27|9917|-80.770346|891|35.052812|NFS-OTHER WINE|0.0|13|REDWOOD CREEK RED BLEND 1.5L|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00085000018705|WINE REMAINING|WINE|-80.771677|80.771680204378441|40|1
35.066546|8ee2c36d324a951b36bad18c50ba3b59b9c7650c|19.98|2014-11-15 15:29:00|1.4091206135396188|1|8500001870|45|0.6120266850020475|0|47|9917|-80.771677|891|35.066546|NFS-OTHER WINE|0.0|13|REDWOOD CREEK RED BLEND 1.5L|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00085000018705|WINE REMAINING|WINE|-80.771677|1.409731706007376|45|2
35.066546|8acf7029f259eda781bdd5dcac96a8b9afded5b5|10.98|2014-12-17 16:41:00|80.782094729586973|1|8087806217|45|35.085677203265348|0|27|3592|-80.78468|1050|35.096737|HAIR STYLING HAIR SPRAY|2.0|17|PANTENE X STRONG HS NON AERO|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00080878062201|HAIR STYLING|HBC|-80.771677|80.771682976423307|30|2
35.066546|878737c9a04519b19f70120860010e27f43b8fa8|7.99|2014-09-16 16:55:00|80.782094729586973|1|4242150024|45|35.085677203265348|0|27|1839|-80.78468|420|35.096737|BH PRESLICED MEATS|0.0|6|BH PRE-SLICED HONEY SMK TURKEY|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00042421500240|PRESLICED MEAT|DELI|-80.771677|80.771682976423307|30|1
35.066546|ca37164ab3cf3f1e1f085b5f8d741e9471ebfc16|25.98|2014-11-19 16:08:00|80.782094729586973|1|3680014780|45|35.085677203265348|0|27|4379|-80.78468|1210|35.096737|ACID BLOCKER-SWALLOW|0.0|17|TC ACID REDUCER MAX STR|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00036800147805|STOMACH REMEDIES|HBC|-80.771677|80.771682976423307|30|2
35.066546|205957de547fc799bc8ef8becb5172811ec892f1|0.72|2014-09-29 17:35:00|80.782094729586973|1||45|35.085677203265348|0|27|502|-80.78468|64|35.096737|FRESH BANANAS|0.0|4|BANANAS, YELLOW|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00204011000008|FRESH PRODUCE|PRODUCE|-80.771677|80.771682976423307|30|1
35.066546|ed40041f7e814898c44a582cea387f5f64060714|0.77|2014-11-06 16:46:00|80.782094729586973|1||45|35.085677203265348|0|27|502|-80.78468|64|35.096737|FRESH BANANAS|0.0|4|BANANAS, YELLOW|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00204011000008|FRESH PRODUCE|PRODUCE|-80.771677|80.771682976423307|30|1
35.066546|e38c273dce1749dd93d6cee9b7923076c24a73f9|3.99|2014-12-24 18:25:00|80.782094729586973|1|2386509984|45|35.085677195695084|0|27|387|-80.739|65|35.141204|NFS-REMAIN CHAR/LOGS/ACC|0.0|1|FLATWOOD NATURAL FIRESTARTER|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00023865099842|CHARCOAL/LOGS/ACCESSORIES|G1 GROCERY|-80.771677|80.771698637821785|171|1
35.066546|fdf3389b5a134c57771e0944c747cea6af7ebd78|7.49|2014-11-25 06:39:00|80.782094729586973|1|2840000288|45|35.085677203265348|0|27|205|-80.78468|31|35.096737|REMAINING SNACKS|0.5|1|FRITOLAY FLAVOR 20 CTN|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00028400002899|SNACKS|G1 GROCERY|-80.771677|80.771682976423307|30|1
35.066546|64aa65638813a80f41d5de56a4edee5f297ad519|7.99|2015-02-27 06:51:00|80.782094729586973|1|2840000288|45|35.085677203265348|0|27|205|-80.78468|31|35.096737|REMAINING SNACKS|1.0|1|FRITOLAY CLASSIC 20 CTN|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00028400002882|SNACKS|G1 GROCERY|-80.771677|80.771682976423307|30|1
35.066546|33284850657e4c7057fcd03e439f4fb547074803|8.19|2014-10-02 17:22:00|80.782094729586973|1|2840000288|45|35.085677203265348|0|27|205|-80.78468|31|35.096737|REMAINING SNACKS|1.2|1|FRITOLAY CLASSIC 20 CTN|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00028400002882|SNACKS|G1 GROCERY|-80.771677|80.771682976423307|30|1
35.066546|6d77b8143241e72ceff91b88fc36cd0526830a85|7.99|2015-01-29 17:37:00|80.782094729586973|1|2840000288|45|35.085677203265348|0|27|205|-80.78468|31|35.096737|REMAINING SNACKS|0.0|1|FRITOLAY CLASSIC 20 CTN|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00028400002882|SNACKS|G1 GROCERY|-80.771677|80.771682976423307|30|1
35.066546|d87093815cbf3b78a63be90676f050721f277294|3.99|2015-02-20 17:20:00|80.782094729586973|1|3338365592|45|35.085677203265348|0|27|561|-80.78468|64|35.096737|FR PROD ORGANIC PRODUCE|0.0|4|ORG GRAPE TOMATOES|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00033383655925|FRESH PRODUCE|PRODUCE|-80.771677|80.771682976423307|30|1
35.066546|4c50a05a17e2a7bf1fcdf665f47aaf220b97310c|2.0|2014-10-02 17:24:00|80.782094729586973|1||45|35.085677203265348|0|27|511|-80.78468|64|35.096737|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00204770000004|FRESH PRODUCE|PRODUCE|-80.771677|80.771682976423307|30|1
35.066546|344f070f906847f5e8892335da6b94188de36746|6.49|2014-10-06 16:50:00|1.4091206135396188|1|4155453973|45|0.6120266850020475|0|47|3030|-80.771677|1000|35.066546|BRAND-MAYBELLINE|0.0|17|071290 MAY MASC GRT LSH DRK BR|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|0.61242566243833529|00041554532982|COSMETICS|HBC|-80.771677|1.409731706007376|45|1
35.066546|fba3dfb739601eddc614c1e0578e2f696e8484a5|3.99|2014-11-11 17:11:00|80.782094729586973|1|3338365548|45|35.085677203265348|0|27|522|-80.78468|64|35.096737|FRESH TOMATOES|0.0|4|ORANGE GLORY TMATOES 16 OZ|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00033383655482|FRESH PRODUCE|PRODUCE|-80.771677|80.771682976423307|30|1
35.066546|a4ee152b0d86dfdea6226b0ec75dd0a6582cb429|7.49|2014-11-06 16:45:00|80.782094729586973|1|2840000288|45|35.085677203265348|0|27|205|-80.78468|31|35.096737|REMAINING SNACKS|0.5|1|DORITOS & CHEETOS 20 CTN|0b7f70489e052674ca8d4a68d9efe4b6a7d67100|1.3219199886349495|35.102887530186244|00028400238243|SNACKS|G1 GROCERY|-80.771677|80.771682976423307|30|1
35.03469|2b6d8b4b4d57182a8223b44bf2681a419b37fb88|8.3|2014-09-21 16:37:00|1.4132775322775095|4|3800043381|82|0.6114706929155321|0|58|1256|-80.97058|13|35.03469|WHOLESOME CRACKERS|3.3|1|SPECIAL K MULTIGRAIN CRACKERS|0ba89b7185d2dc737c2155b17ebc7fe0ed00c72f|2.6054106043673597|0.61177642288969325|00038000433818|CRACKERS|G1 GROCERY|-80.97058|1.4132032182494703|82|2
35.03469|33bded26d9c7ede0edf65e10db5cf0b14a86f4f8|3.35|2015-02-13 17:06:00|1.4132775322775095|4|2529300098|82|0.6114706929155321|0|58|1265|-80.97058|57|35.03469|ALMOND MILK|0.0|3|SILK PURE ALMOND UNSWEETENED|0ba89b7185d2dc737c2155b17ebc7fe0ed00c72f|2.6054106043673597|0.61177642288969325|00025293001497|MILK|DAIRY|-80.97058|1.4132032182494703|82|1
35.03469|82884e24033d366d84c5f756ecaaf9509277ac2c|3.29|2014-11-08 17:37:00|1.4132775322775095|4|71514150349|82|0.6114706929155321|0|58|330|-80.97058|55|35.03469|EGGS|0.0|3|EGGLAND BEST GRADE A LARGE EGG|0ba89b7185d2dc737c2155b17ebc7fe0ed00c72f|2.6054106043673597|0.61177642288969325|00715141503494|EGGS FRESH|DAIRY|-80.97058|1.4132032182494703|82|1
35.103409|f7fbabc47411419a487f6900e7d19770295392b9|8.98|2015-02-28 09:31:00|80.992192682720116|2|75703751693|88|35.113590041033326|0|56|420|-80.97058|71|35.03469|NFS-SOIL/SPOT/STAIN REMO|3.98|1|OXI CLEAN LAUNDRY STAIN REMOVR|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00757037516935|LAUNDRY SUPPLIES|G1 GROCERY|-80.992182|80.992189682913178|82|2
35.103409|c1f2a92cb3f292e7741f1d7f7cc53c3f8f4e7811|9.38|2015-01-10 09:29:00|80.992192682720116|2|7261345111|88|35.113590041033326|0|56|417|-80.97058|71|35.03469|NFS-FABRIC SOFTENERS|3.38|1|SNUGGLE SPARKLE SHEETS 80CT|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00072613451111|LAUNDRY SUPPLIES|G1 GROCERY|-80.992182|80.992189682913178|82|2
35.103409|65f97917bf09efa56b8815476d1a93461029865c|2.79|2014-11-02 10:01:00|1.4132775322775095|2|1800000501|88|0.6126700657242101|0|58|327|-80.992182|54|35.103409|DINNER ROLLS-REFRIGERATED|0.0|3|PILLSBURY CINN CREAM CHS ROLLS|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00018000005123|DOUGH PRODUCTS|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|ca2020bf07db9971768dd0d89880718c7a5eb34c|1.29|2014-12-24 08:08:00|80.992192682720116|2|2700039014|88|35.113590041033326|0|56|257|-80.97058|39|35.03469|TOMATOES|0.29|1|HUNTS TOMATO SAUCE 15|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00027000390146|VEGETABLES-CAN/JAR|G1 GROCERY|-80.992182|80.992189682913178|82|1
35.103409|ed84a9f559ea3ca0c07e09043238ae3afed5054a|6.38|2015-02-14 08:49:00|80.992192682720116|2|2220094152|88|35.113590041033326|0|56|3876|-80.97058|1070|35.03469|SOLID-MALE|0.69|17|SPEED STICK AP/DEO REGULAR|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00022200941525|DEODORANT|HBC|-80.992182|80.992189682913178|82|2
35.103409|abde5ac982c48a14f1124496114492b59f0bb168|1.38|2014-12-20 08:26:00|80.992192682720116|2|3080000973|88|35.113590041033326|0|56|727|-80.97058|7|35.03469|SEASONAL CANDY-SINGLE FAC|0.34|1|I/O(C15)SPNGLR PPRMNT R&W|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00030800009736|CANDY|G1 GROCERY|-80.992182|80.992189682913178|82|2
35.103409|b68fd3617119870b31c04809aae829466035ce04|1.99|2015-01-03 08:43:00|80.992192682720116|2|3700035716|88|35.113590041033326|0|56|422|-80.97058|71|35.03469|NFS-REMAIN LAUNDRY SUPPL|0.0|1|E  DOWNY BALL DISPENSER|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00037000357162|LAUNDRY SUPPLIES|G1 GROCERY|-80.992182|80.992189682913178|82|1
35.103409|16748038ffabe212469cea664abe151d5278eaa3|4.99|2014-11-24 14:25:00|1.4132775322775095|2|7203688187|88|0.6126700657242101|0|58|561|-80.992182|64|35.103409|FR PROD ORGANIC PRODUCE|0.0|4|ORG HT BABY SPINACH 11 OZ|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00072036881878|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|1
35.103409|a64977087e3a380360d6b3ab77acb80f417c01e7|4.79|2014-10-18 09:37:00|80.992192682720116|2|7203676457|88|35.113590041033326|0|56|312|-80.97058|51|35.03469|BUTTER|0.0|3|HTO ORGANIC BUTTER SALTED|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00072036763419|BUTTER & MARGARINE|DAIRY|-80.992182|80.992189682913178|82|1
35.103409|0cf65f23f26e9a5a751ced9f9226bd3535d83f72|5.99|2014-10-29 18:29:00|80.992192682720116|2|8500001444|88|35.113590041966788|0|56|9938|-80.994596|885|35.061685|NFS POP PINOT GRS/GRIGIO|0.0|13|CB-BAREFOOT PINOT GRIGIO|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00085000014448|POPULAR (4-$7.99)|WINE|-80.992182|80.99218753400686|475|1
35.103409|b89f496e558e8564083bd9ec8bc08ab1917c1eb4|0.91|2015-02-14 14:57:00|1.4132775322775095|2||88|0.6126700657242101|0|58|527|-80.992182|64|35.103409|FRESH CARROTS|0.0|4|COO CARROTS, BULK|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00204562000007|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|1
35.103409|b19557846e83725ee9e7b41fa70ea094262264be|0.44|2015-03-08 13:44:00|80.992192682720116|2||88|35.113590041966788|0|56|522|-80.994596|64|35.061685|FRESH TOMATOES|0.0|4|COO RED ROMA TOMATOES|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00204087000001|FRESH PRODUCE|PRODUCE|-80.992182|80.99218753400686|475|1
35.103409|ae7386b80ce354cf70a3744e5d3dd562f0ba910a|17.33|2015-03-07 10:44:00|1.4132775322775095|2|20943700000|88|0.6126700657242101|0|58|664|-80.992182|145|35.103409|SHRIMP WILD CAUGHT|10.2|12|WC ARGENTINA PINK SHRIMP 16/20|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00209437000007|SHRIMP|SEAFOOD|-80.992182|1.413580244274486|88|1
35.103409|2488c23f7aec85a454d2ae4775d7116c3993c600|2.29|2015-01-11 11:02:00|80.992192682720116|2|31254662920|88|35.113590041966788|0|56|4207|-80.994596|1200|35.061685|COUGH DROP-ADULT|0.79|17|HALLS DEF VIT. C WMLN-63158|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00312546631588|COUGH/COLD/SINUS|HBC|-80.992182|80.99218753400686|475|1
35.103409|773be46328abb173251fb92ab443c04ac86ed2ec|2.6|2014-12-13 08:42:00|80.992192682720116|2||88|35.113590041033326|0|56|502|-80.97058|64|35.03469|FRESH BANANAS|0.0|4|BANANAS, YELLOW|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00204011000008|FRESH PRODUCE|PRODUCE|-80.992182|80.992189682913178|82|2
35.103409|7248292743602bbf4b6c1d9d4c73ad3892122876|1.25|2014-11-29 08:32:00|80.992192682720116|2||88|35.113590041033326|0|56|502|-80.97058|64|35.03469|FRESH BANANAS|0.0|4|BANANAS, YELLOW|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00204011000008|FRESH PRODUCE|PRODUCE|-80.992182|80.992189682913178|82|1
35.103409|6c4765334296c01802d6b6109aa7aa8536b61254|0.55|2015-02-21 09:51:00|1.4132775322775095|2||88|0.6126700657242101|0|58|502|-80.992182|64|35.103409|FRESH BANANAS|0.0|4|BANANAS, YELLOW|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00204011000008|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|1
35.103409|9631120e5765923314d29123f9250204e0fb733d|3.59|2014-11-26 12:07:00|1.4132775322775095|2|4850002013|88|0.6126700657242101|0|58|335|-80.992182|56|35.103409|ORANGE JUICE-REGRIGERATED|0.59|3|TROPICANA PP W/CALCIUM|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00048500305690|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|3b60d8e7029a48eb65a725a56c8386ff5d8fa486|19.49|2015-01-31 09:39:00|80.992192682720116|2|30259319282|88|35.113590041033326|0|56|4844|-80.97058|1235|35.03469|FIRST AID TREATMENT|0.0|17|MEDERMA CREAM W/SPF 30|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00302593192828|FIRST AID|HBC|-80.992182|80.992189682913178|82|1
35.103409|2e96c0b0e690cc21cb44e066023f2f17a8eeba23|6.39|2015-01-11 13:43:00|1.4132775322775095|2|4154800385|88|0.6126700657242101|0|58|252|-80.992182|45|35.103409|PREMIUM ICE CREAM|3.2|5|EDY'S SLOW CHURNED LIMITED E|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00041548451862|ICE CREAM|FROZEN|-80.992182|1.413580244274486|88|1
35.103409|3a0132af0f2686ba6cdd604a4f6b96847b46d2f9|3.19|2015-03-07 08:30:00|80.992192682720116|2|1600027532|88|35.113590041033326|0|56|81|-80.97058|9|35.03469|RTE CEREAL KIDS|1.6|1|GM TRIX|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00016000275324|CEREAL|G1 GROCERY|-80.992182|80.992189682913178|82|1
35.103409|e9c667997d40521c5bd2cbc4e8b9314a1cc79488|2.79|2014-09-13 09:10:00|80.992192682720116|2|1600042060|88|35.113590041033326|0|56|13|-80.97058|2|35.03469|ROLLS/BISCUIT MIXES|1.29|1|BC BISQUICK|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00016000420601|BAKING MIXES|G1 GROCERY|-80.992182|80.992189682913178|82|1
35.103409|77a5ae5c25eafabcc2d4b32d91ca19ebc136d08b|1.0|2014-10-07 07:46:00|80.992192682720116|2|812|88|35.113590041966788|0|56|1639|-80.994596|377|35.061685|BULK (DONUTS)|0.0|14|NEW BULK DONUT CODE|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00000000008120|DONUTS|BAKERY|-80.992182|80.99218753400686|475|1
35.103409|41aabfb843edb17647a92c4f7e0b857b4902292c|2.0|2015-01-17 08:26:00|80.992192682720116|2|812|88|35.113590041033326|0|56|1639|-80.97058|377|35.03469|BULK (DONUTS)|0.0|14|NEW BULK DONUT CODE|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00000000008120|DONUTS|BAKERY|-80.992182|80.992189682913178|82|2
35.103409|1c02620cf267f1966a441ff2f6f396e7b7e9b9fb|1.0|2014-10-07 07:44:00|80.992192682720116|2|812|88|35.113590041966788|0|56|1639|-80.994596|377|35.061685|BULK (DONUTS)|0.0|14|NEW BULK DONUT CODE|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00000000008120|DONUTS|BAKERY|-80.992182|80.99218753400686|475|1
35.103409|d71a82666cd263f1b4d79dbebfd463d002961583|3.49|2014-11-10 17:22:00|1.4132775322775095|2|4178000211|88|0.6126700657242101|0|58|202|-80.992182|31|35.103409|PRETZELS|0.7|1|UTZ HOLIDAY SHAPED PRETZELS|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00041780022882|SNACKS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|6dc606e93cd7ec89759e8abb2b051eed21b8b991|20.99|2014-11-01 13:15:00|80.992192682720116|2|7499904067|88|35.113590041966788|0|56|8068|-80.994596|1700|35.061685|HOUSEHOLD STEAM CLEANER|0.0|18|RUG DR PET FORMULA CARPET CLNR|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00074999040675|CARPET CLEANING/RENTAL|GM|-80.992182|80.99218753400686|475|1
35.103409|749a8491e88dfb65ee8bdd64d16ffe5eedae6795|9.99|2014-12-06 12:57:00|1.4132775322775095|2|7674007012|88|0.6126700657242101|0|58|62|-80.992182|7|35.103409|SPECIALTY BAR/BOX CHOCOLATE|3.0|1|WHITMAN SAMPLER BOX PP9.99|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00076740070122|CANDY|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|b6fa4340b4bdff85624cae13e85c400707b2687b|6.1|2014-10-11 13:43:00|1.4132775322775095|2||88|0.6126700657242101|0|58|503|-80.992182|64|35.103409|FRESH GRAPES|3.06|4|RED GRAPES, SEEDLESS|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00204635000002|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|1
35.103409|c35520c881e49ca1e2528188fbe7b413e8ad6295|6.95|2014-10-05 12:50:00|1.4132775322775095|2|20889700000|88|0.6126700657242101|0|58|660|-80.992182|154|35.103409|FISH FILLETS WILD CGHT|1.75|12|WC FROZ  SWORDFISH STKS (EC)|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00208897000008|FISH FILLETS/STEAKS|SEAFOOD|-80.992182|1.413580244274486|88|1
35.103409|9d8631eca56b3f7885ed650b25e083fee1371583|4.49|2014-12-19 18:46:00|1.4132775322775095|2|4198500007|88|0.6126700657242101|0|58|9924|-80.992182|882|35.103409|NFS-PREMIUM BOX|0.0|13|FOXHORN MERLOT 500ml|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00041985000074|PREMIUM BOX|WINE|-80.992182|1.413580244274486|88|1
35.103409|2558822984be7b21ac14beb0d482ac5cf56cad28|12.98|2014-12-22 18:35:00|1.4132775322775095|2|4000024908|88|0.6126700657242101|0|58|46|-80.992182|7|35.103409|PKG CHOC|3.24|1|M&M PEANUT LARGE BAG|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00040000249290|CANDY|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|f71bfd4231bf3aef23dd9bae317b140953b14aa5|2.99|2015-02-13 18:26:00|1.4132775322775095|2|4610001992|88|0.6126700657242101|0|58|317|-80.992182|52|35.103409|CHUNK AND BAR CHEESE|0.49|3|SARGENTO FIESTA PEPPER JACK|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00046100019931|CHEESE|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|87c7f95d2a998f7d136127559a5da09e900a4789|5.58|2015-01-13 07:58:00|1.4132775322775095|2|5200032669|88|0.6126700657242101|0|58|171|-80.992182|20|35.103409|ISOTONIC DRINKS|0.82|1|GATORADE G2 GRAPE|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00052000640014|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|527b904c5158f1c19ffdd7a067b140a5719aaeb9|2.79|2014-09-20 08:04:00|1.4132775322775095|2|5200032669|88|0.6126700657242101|0|58|171|-80.992182|20|35.103409|ISOTONIC DRINKS|0.29|1|GATORADE G2 GRAPE|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00052000640014|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|dd573a2db044cf33f30be7464465e37ed8fd4daf|2.79|2015-01-25 15:56:00|80.992192682720116|2|5200032669|88|35.113590041966788|0|56|171|-80.994596|20|35.061685|ISOTONIC DRINKS|0.41|1|GATORADE G2 GRAPE|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00052000640014|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.992182|80.99218753400686|475|1
35.103409|1e76f8de23003684833d163b50eb43d5d5389edf|2.79|2014-12-27 07:39:00|1.4132775322775095|2|5200032669|88|0.6126700657242101|0|58|171|-80.992182|20|35.103409|ISOTONIC DRINKS|0.41|1|GATORADE G2 GRAPE|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00052000640014|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|53443bc99b13805e0a696029b0250d87e8bb86d4|2.79|2015-01-31 07:43:00|1.4132775322775095|2|5200032669|88|0.6126700657242101|0|58|171|-80.992182|20|35.103409|ISOTONIC DRINKS|0.41|1|GATORADE G2 GRAPE|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00052000640014|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|8cd28adda0bed969820dfb23960dd8a408a7d03f|3.68|2015-01-17 16:15:00|1.4132775322775095|2|20557100000|88|0.6126700657242101|0|58|1820|-80.992182|410|35.103409|BH BEEF|0.0|6|BOARS HEAD LONDON BROIL|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00205571000002|BH MEAT|DELI|-80.992182|1.413580244274486|88|1
35.103409|84ef3d209f7116dc470d7c9e94a77619c1d43ef8|2.23|2014-10-04 13:20:00|1.4132775322775095|2||88|0.6126700657242101|0|58|561|-80.992182|64|35.103409|FR PROD ORGANIC PRODUCE|0.32|4|ORG TOMATOES|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00294064000001|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|1
35.103409|3223c33ac33694d822b0d6c93be93c651b639312|0.43|2015-02-08 14:29:00|80.992192682720116|2||88|35.113590041966788|0|56|522|-80.994596|64|35.061685|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00204664000004|FRESH PRODUCE|PRODUCE|-80.992182|80.99218753400686|475|1
35.103409|6fe6f07562aefa57becde813a167257f6dc043fd|0.42|2014-10-25 15:13:00|1.4132775322775095|2||88|0.6126700657242101|0|58|524|-80.992182|64|35.103409|FRESH PROD FRESH ONIONS|0.0|4|COO YELLOW ONIONS, LRG|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00204665000003|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|1
35.103409|0ce48c7270c98a90a0de6f79e3018e64f66ad31e|5.0|2015-01-31 15:51:00|80.992192682720116|2|8500001581|88|35.113590041966788|0|56|9943|-80.994596|885|35.061685|NFS POP RIESLING|0.0|13|BAREFOOT RIESLING|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00085000015810|POPULAR (4-$7.99)|WINE|-80.992182|80.99218753400686|475|1
35.103409|c082477815af58a493d0605a2bea41ef90e19012|6.99|2014-11-01 11:39:00|1.4132775322775095|2|7203695946|88|0.6126700657242101|0|58|1295|-80.992182|383|35.103409|PIES PASTRY CASE TAX|2.0|14|"9"" CHOCOLATE SILK PIE"|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00072036959461|PASTRY CASE|BAKERY|-80.992182|1.413580244274486|88|1
35.103409|bfed5b3b1c40a22817070f906a5c0792a16be439|3.29|2014-12-21 12:33:00|1.4132775322775095|2|2840004768|88|0.6126700657242101|0|58|202|-80.992182|31|35.103409|PRETZELS|0.29|1|ROLD GOLD CHEDDAR CHEESE PRETL|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00028400021869|SNACKS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|9f6b180ae3c2839e1be99ee1102eec5c0cec99cb|3.29|2015-01-18 14:08:00|80.992192682720116|2|2840004768|88|35.113590041033326|0|56|202|-80.97058|31|35.03469|PRETZELS|1.65|1|ROLD GOLD CHEDDAR CHEESE PRETL|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00028400021869|SNACKS|G1 GROCERY|-80.992182|80.992189682913178|82|1
35.103409|e9622c2803d293717d2e403d35480fcf78358334|2.99|2014-11-07 13:47:00|1.4132775322775095|2|20789900000|88|0.6126700657242101|0|58|1677|-80.992182|383|35.103409|INDIVIDUALS (PASTRY CASE)|0.0|14|MEGA CHARACTER CUPCAKE|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00207899000009|PASTRY CASE|BAKERY|-80.992182|1.413580244274486|88|1
35.103409|5d64de0bdfa99ee6df5524e06e0471c7175ba1fe|9.98|2015-01-23 17:51:00|1.4132775322775095|2|8500002254|88|0.6126700657242101|0|58|9943|-80.992182|885|35.103409|NFS POP RIESLING|0.0|13|GALLO FMLY VINEYARDS RIESLING|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00085000022542|POPULAR (4-$7.99)|WINE|-80.992182|1.413580244274486|88|2
35.103409|03512fd897478ebbada631e17d97d42491aadb90|9.98|2015-02-08 14:45:00|1.4132775322775095|2|8500002254|88|0.6126700657242101|0|58|9943|-80.992182|885|35.103409|NFS POP RIESLING|0.0|13|GALLO FMLY VINEYARDS RIESLING|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00085000022542|POPULAR (4-$7.99)|WINE|-80.992182|1.413580244274486|88|2
35.103409|4bd8da8d64cc4b8cf22e1179e821bd216edeabab|4.99|2015-01-18 12:31:00|1.4132775322775095|2|2840003400|88|0.6126700657242101|0|58|201|-80.992182|31|35.103409|POTATO CHIPS|1.0|1|RUFFLES ORIGINAL|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00028400034005|SNACKS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|9c95f316c0c5dcf698ca4805172d3c42f67739cf|5.97|2014-12-27 15:50:00|80.992192682720116|2|7203676359|88|35.113590041966788|0|56|345|-80.994596|57|35.061685|ORGANIC MILK|0.0|3|HTO ORGANIC 2% MILK GAL|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00072036763600|MILK|DAIRY|-80.992182|80.99218753400686|475|1
35.103409|c7e025419a7a7d2994a70f2c80d922edcdf3860e|1.68|2015-01-12 11:33:00|80.992192682720116|2|20579000000|88|35.113590041966788|0|56|1824|-80.994596|410|35.061685|BH LOAVES|0.42|6|BOARS HEAD LOWER SODIUM BOLGNA|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00205790000005|BH MEAT|DELI|-80.992182|80.99218753400686|475|1
35.103409|ad6c6d3e7a145ce7007734ffbb36a1b4dff45bf7|3.99|2014-12-06 09:05:00|80.992192682720116|2||88|35.113590041033326|0|56|512|-80.97058|64|35.03469|FRSH PROD FRSH FRUIT REM|0.0|4|POMEGRANATES  STACKER|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00233440000006|FRESH PRODUCE|PRODUCE|-80.992182|80.992189682913178|82|1
35.103409|3747a87d185df592eb87fbc2f800779e9aed4aaf|7.96|2014-11-15 08:51:00|80.992192682720116|2|3040080888|88|35.113590041033326|0|56|424|-80.97058|72|35.03469|NFS-FACIAL TISSUE|3.96|1|ANGEL SOFT FACIAL TISSUE 165CT|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00030400819100|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.992182|80.992189682913178|82|4
35.103409|7f757cdb2942ee816e78ab0ea4ac296cfb810704|4.29|2014-11-02 12:11:00|80.992192682720116|2|2840006399|88|35.113590041966788|0|56|204|-80.994596|31|35.061685|TORTILLA CHIPS|1.79|1|TOSTITOS FAJITAS SCOOPS|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00028400220538|SNACKS|G1 GROCERY|-80.992182|80.99218753400686|475|1
35.103409|7acd136c7a062a995f8d8bf8da852475fab03c40|4.29|2014-12-14 12:58:00|80.992192682720116|2|2840006399|88|35.113590041966788|0|56|204|-80.994596|31|35.061685|TORTILLA CHIPS|1.29|1|TOSTITOS FAJITAS SCOOPS|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00028400220538|SNACKS|G1 GROCERY|-80.992182|80.99218753400686|475|1
35.103409|313e654308292d9abf7c4225eb1b017439fb6d9a|3.58|2015-01-11 11:17:00|80.992192682720116|2|1700000300|88|35.113590041966788|0|56|429|-80.994596|73|35.061685|NFS-BAR SOAP|0.58|1|DIAL BASIC HYPOALLERGENIC 3BAR|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00017000003009|PERSONAL SOAP/BATH ADDITIVES|G1 GROCERY|-80.992182|80.99218753400686|475|2
35.103409|64bcb01a0101cb9c80c256a4c08f5ec2559be1e0|14.98|2015-01-03 11:11:00|1.4132775322775095|2|3040021526|88|0.6126700657242101|0|58|426|-80.992182|72|35.103409|NFS-PAPER TOWELS|3.0|1|SPARKLE 8 RL REGULAR PRINT|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00030400216503|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|75eb17f93f7c9c4af5ff146787e08ba645d8d923|1.67|2014-09-25 09:09:00|1.4132775322775095|2|1070002152|88|0.6126700657242101|0|58|53|-80.992182|7|35.103409|THEATER BOX|0.0|1|E  REESE PIECES BIG BOX|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00034000114702|CANDY|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|525a1d1076bade752a3c453372a238e853034b8d|13.79|2014-09-29 07:24:00|80.992192682720116|2|76394804293|88|35.113590041966788|0|56|4531|-80.994596|1215|35.061685|SPLMNT-DIGESTIVE AID|3.0|17|(JHK) ACIDOPHILUS PEARLS|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00763948042937|VITAMINS & SUPPLEMENTS|HBC|-80.992182|80.99218753400686|475|1
35.103409|aa0a6394368f3c23359ef5091964cdfa4726b390|2.59|2014-09-23 17:09:00|1.4132775322775095|2|7203695299|88|0.6126700657242101|0|58|1654|-80.992182|381|35.103409|DESSERT CAKES|0.0|14|TRIPLE COCONUT SLICE|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00072036952998|CAKES|BAKERY|-80.992182|1.413580244274486|88|1
35.103409|74a9a68cf186f6a4ed75af4f583f0e9ae343ef6c|11.98|2015-01-19 07:19:00|80.992192682720116|2|7203695041|88|35.113590041966788|0|56|1654|-80.994596|381|35.061685|DESSERT CAKES|0.0|14|2 CT. CHOC OVERLOAD TORTE|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00072036950413|CAKES|BAKERY|-80.992182|80.99218753400686|475|2
35.103409|80129caec2d78d2f0d16581b122864b9bc110bab|7.95|2014-12-24 08:09:00|80.992192682720116|2|76211160216|88|35.113590041033326|0|56|1595|-80.97058|370|35.03469|WHOLE BEANS|3.18|22|CHRISTMAS COFFEE WB 8 OZ|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00762111602169|STARBUCKS|COFFEE SHOP|-80.992182|80.992189682913178|82|1
35.103409|cf04a4c8c01e84e2aac8a8f3175b6158d9df170e|2.79|2014-12-17 09:13:00|1.4132775322775095|2|1130038110|88|0.6126700657242101|0|58|50|-80.992182|7|35.103409|PEG CANDY|0.0|1|BRACHS SPICE DROPS|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00011300741647|CANDY|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|97eaf74138299353cc07bd5e32e65dbb249dff0f|1.87|2014-12-17 15:04:00|1.4132775322775095|2|7203670210|88|0.6126700657242101|0|58|399|-80.992182|69|35.103409|NFS-DISINFECTANTS|0.0|1|YH DISINFECTING WIPES LEMON|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00072036702111|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|f580c8573eb094cec7d0f6ef045716c12d3b7ffc|1.87|2014-12-29 17:27:00|1.4132775322775095|2|7203670210|88|0.6126700657242101|0|58|399|-80.992182|69|35.103409|NFS-DISINFECTANTS|0.0|1|YH DISINFECTING WIPES LEMON|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00072036702111|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|ead11ca5114b29fa8b4ee88d023aa25d4158a24e|10.35|2015-02-14 08:57:00|80.992192682720116|2|4460030438|88|35.113590041033326|0|56|730|-80.97058|24|35.03469|NFS-CAT LITTER|5.18|1|FRESH STEP SCOOP MULTI CAT LIT|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00044600304380|PET FOOD/SUPPLIES|G1 GROCERY|-80.992182|80.992189682913178|82|1
35.103409|cc44f211bd99c7fb8f106dd64446024b9c221c6f|103.49999999999999|2015-02-12 17:26:00|1.4132775322775095|2|4460030438|88|0.6126700657242101|0|58|730|-80.992182|24|35.103409|NFS-CAT LITTER|5.18|1|FRESH STEP SCOOP MULTI CAT LIT|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00044600304380|PET FOOD/SUPPLIES|G1 GROCERY|-80.992182|1.413580244274486|88|10
35.103409|9fab6928e1739f6d920e6d62dfbb15d669282e29|103.49999999999999|2015-02-11 08:17:00|80.992192682720116|2|4460030438|88|35.113590041033326|0|56|730|-80.97058|24|35.03469|NFS-CAT LITTER|5.18|1|FRESH STEP SCOOP MULTI CAT LIT|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00044600304380|PET FOOD/SUPPLIES|G1 GROCERY|-80.992182|80.992189682913178|82|10
35.103409|2cc00880aa7fc709f35964881df2903092056290|41.4|2015-02-11 07:58:00|80.992192682720116|2|4460030438|88|35.113590041966788|0|56|730|-80.994596|24|35.061685|NFS-CAT LITTER|5.18|1|FRESH STEP SCOOP MULTI CAT LIT|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00044600304380|PET FOOD/SUPPLIES|G1 GROCERY|-80.992182|80.99218753400686|475|4
35.103409|75395f9d8cd1477807aafb9ccfefa08b702959ae|134.54999999999998|2015-02-14 08:30:00|1.4132775322775095|2|4460030438|88|0.6126700657242101|0|58|730|-80.992182|24|35.103409|NFS-CAT LITTER|0.0|1|FRESH STEP SCOOP MULTI CAT LIT|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00044600304380|PET FOOD/SUPPLIES|G1 GROCERY|-80.992182|1.413580244274486|88|13
35.103409|2e5c9f0dff79cd2dd343c7bb0c0ae25085a31c34|20.7|2015-02-13 15:29:00|80.992192682720116|2|4460030438|88|35.113590041966788|0|56|730|-80.994596|24|35.061685|NFS-CAT LITTER|5.17|1|FRESH STEP SCOOP MULTI CAT LIT|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00044600304380|PET FOOD/SUPPLIES|G1 GROCERY|-80.992182|80.99218753400686|475|2
35.103409|ae8d1943350011adccc3697ec8a24009f6725f71|1.35|2015-01-10 11:29:00|1.4132775322775095|2||88|0.6126700657242101|0|58|500|-80.992182|64|35.103409|FRESH APPLES|0.13|4|GALA APPLES|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00204135000007|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|1
35.103409|e2f0d0590529ead0fd214ba45ef8a9abab246c5a|2.0|2014-09-28 20:32:00|80.992192682720116|2|78352032108|88|35.113590041966788|0|56|8598|-80.994596|1792|35.061685|NEWSPAPERS|0.0|18|SUNDAY CHARLOTTE OBSERVER|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00783520321083|NEWSPAPERS|GM|-80.992182|80.99218753400686|475|1
35.103409|a5382d1f429715a878b566ba8c53b5f7b1b050d8|7.99|2015-02-07 12:48:00|1.4132775322775095|2|3700014389|88|0.6126700657242101|0|58|388|-80.992182|66|35.103409|NFS-DISHWASH PWDR/LIQUID|2.0|1|CASCADE DAWN FRESH SCENT 32CT|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00037000143895|DETERGENTS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|5493dafe6f6a9c3dfcfa7456651b28debe6c397d|2.31|2014-10-22 12:54:00|80.992192682720116|2|20037600000|88|35.113590041966788|0|56|1801|-80.994596|400|35.061685|FFM TURKEY|0.0|6|TURKEY BREAST|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00200376000004|FFM MEAT|DELI|-80.992182|80.99218753400686|475|1
35.103409|a8f588b3e9c908783ed807f598a038cee183dcb0|3.15|2014-11-14 12:35:00|80.992192682720116|2|20037600000|88|35.113590041966788|0|56|1801|-80.994596|400|35.061685|FFM TURKEY|0.0|6|TURKEY BREAST|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00200376000004|FFM MEAT|DELI|-80.992182|80.99218753400686|475|1
35.103409|a673b9963af3d4755e0f947e712c61ae66119dbf|3.15|2014-09-10 13:08:00|1.4132775322775095|2|20037600000|88|0.6126700657242101|0|58|1801|-80.992182|400|35.103409|FFM TURKEY|0.0|6|TURKEY BREAST|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00200376000004|FFM MEAT|DELI|-80.992182|1.413580244274486|88|1
35.103409|461952e3e0cd6c38f74b3e9a6cd843df6387b70f|1.75|2014-10-21 16:50:00|80.992192682720116|2|20037600000|88|35.113590041966788|0|56|1801|-80.994596|400|35.061685|FFM TURKEY|0.0|6|TURKEY BREAST|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00200376000004|FFM MEAT|DELI|-80.992182|80.99218753400686|475|1
35.103409|cce4f1b39131585e04bc4d5db65c80a2845320a6|2.45|2014-12-05 14:02:00|1.4132775322775095|2|20037600000|88|0.6126700657242101|0|58|1801|-80.992182|400|35.103409|FFM TURKEY|0.0|6|TURKEY BREAST|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00200376000004|FFM MEAT|DELI|-80.992182|1.413580244274486|88|1
35.103409|5459cc78c00320f3a25b717e8379c82380b79200|3.5|2014-10-03 13:47:00|1.4132775322775095|2|20037600000|88|0.6126700657242101|0|58|1801|-80.992182|400|35.103409|FFM TURKEY|0.0|6|TURKEY BREAST|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00200376000004|FFM MEAT|DELI|-80.992182|1.413580244274486|88|1
35.103409|35cbff9f68392bb6b2eeee1fc0b139c0ab40a3d0|21.98|2014-10-25 09:47:00|80.992192682720116|2|3040077569|88|35.113590041033326|0|56|427|-80.97058|72|35.03469|NFS-TOILET TISSUE|6.0|1|ANGEL SOFT SOFT/STRONG 16R|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00030400775697|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.992182|80.992189682913178|82|2
35.103409|758b9391a6a76128968a51cf58e0380a380444b5|0.75|2014-12-12 13:28:00|1.4132775322775095|2||88|0.6126700657242101|0|58|1617|-80.992182|373|35.103409|ROLLS BULK|0.0|14|BULK ROLLS|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00072036955555|ROLLS|BAKERY|-80.992182|1.413580244274486|88|1
35.103409|4153bf8186c3122ae5d315ce912e1630df7e0f60|1.99|2014-10-21 12:20:00|1.4132775322775095|2|1130082079|88|0.6126700657242101|0|58|727|-80.992182|7|35.103409|SEASONAL CANDY-SINGLE FAC|0.4|1|I/O(H15)BRACH AUTUMN MIX|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00011300820793|CANDY|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|b40dd3e1f71d25e0fc3f1dc55282979323a3744d|1.69|2014-10-27 12:28:00|1.4132775322775095|2|5200033875|88|0.6126700657242101|0|58|171|-80.992182|20|35.103409|ISOTONIC DRINKS|0.69|1|GATORADE G2 GRAPE|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|0.61177642288969325|00052000321999|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|b720b060aab60ece854d95a5f8da88eeea136c04|5.07|2014-11-03 06:30:00|80.992192682720116|2|5200033875|88|35.113590041966788|0|56|171|-80.994596|20|35.061685|ISOTONIC DRINKS|1.38|1|GATORADE G2 GRAPE|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00052000321999|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.992182|80.99218753400686|475|3
35.103409|ac0f130707189c4f51279103f4861473b4eb4f22|3.99|2014-10-31 17:50:00|80.992192682720116|2|7203663061|88|35.113590041966788|0|56|364|-80.994596|55|35.061685|ORGANIC AND CF EGGS|0.0|3|HTO ORGANIC GRD A LARGE EGG BR|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00072036630612|EGGS FRESH|DAIRY|-80.992182|80.99218753400686|475|1
35.103409|2b975246aad222a3de2cb54dfc073ff743fc89c6|10.19|2015-02-15 15:33:00|80.992192682720116|2|20839500000|88|35.113590041966788|0|56|660|-80.994596|154|35.061685|FISH FILLETS WILD CGHT|4.8|12|WC FROZ TUNA STKS (VT)|1250b3b110a203740fe9cf780bf356104429927b|0.7034854831191146|35.113093007298254|00208395000005|FISH FILLETS/STEAKS|SEAFOOD|-80.992182|80.99218753400686|475|1
34.977331|8c2dcef6b3fa56743fc44501e80d26e0809df003|7.99|2015-01-27 17:49:00|80.992238315890603|4|7100750742|149|35.235114700239841|0|22|1277|-80.992182|279|35.103409|FROZEN SNACKS|0.0|5|EL MONTEREY BEEF TAMALES|13188e51f8cbcdb0f4446979d52b31776501ed23|17.812250445069584|35.131650835559327|00071007507427|FROZEN SANDWICH AND SNACKS|FROZEN|-81.027334|81.027797670546974|88|1
34.977331|68c2879a6941d9060fc3e55bea6e3c69576b33c7|5.29|2014-12-20 15:12:00|80.992238315890603|4|7203695450|149|35.235114700239841|0|22|1603|-80.992182|371|35.103409|PRIVATE LABEL BREAD|1.8|14|BAND OF BAKERS HARVEST BREAD|13188e51f8cbcdb0f4446979d52b31776501ed23|17.812250445069584|35.131650835559327|00072036954503|BREAD|BAKERY|-81.027334|81.027797670546974|88|1
35.41832|359c0e7d70b4b3b2a1df45004a5675f0fe219e62|3.19|2014-09-20 16:37:00|80.749667378538092|2|3400014830|190|35.464876711042834|0|3|16|-80.662946|3|35.412407|BAKING CHOCOLATE/CHIPS/MORSELS|0.0|1|HEATH BITS O BRICKLE TOFFEE|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00034000061808|BAKING SUPPLIES|G1 GROCERY|-80.746334|80.746352221258178|68|1
35.41832|09f5326b6802e222e233e82ceeae304a3d6209a2|3.65|2015-03-07 14:43:00|80.749667378538092|2|3010001610|190|35.464876711042834|0|3|1254|-80.662946|12|35.412407|FUDGE ENROBED|0.0|1|FUDGE SHOPPE  COCONUT DREAMS|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00030100505617|COOKIES|G1 GROCERY|-80.746334|80.746352221258178|68|1
35.41832|e0474fb3f41e0600fa54d665a5bdf0ecc6edbc6c|1.99|2014-11-05 19:44:00|80.749667378538092|2|5100017520|190|35.464876580478958|0|3|1201|-80.8438|33|35.23102|RTS CANNED|0.49|1|CAM HOMESTYLE CHICKEN NOODLE|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00051000016591|SOUP|G1 GROCERY|-80.746334|80.746470557922436|205|1
35.41832|fa1305dc88df44a9a5f53e5882d658a423cf35c0|3.99|2015-03-07 17:05:00|80.749667378538092|2|3260190085|190|35.464876580478958|0|3|561|-80.8438|64|35.23102|FR PROD ORGANIC PRODUCE|0.0|4|EBF ORG BABY LETTUCE 5 OZ|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00032601900854|FRESH PRODUCE|PRODUCE|-80.746334|80.746470557922436|205|1
35.41832|6563bcd20262f3246dc28534ff79a1f73227eb5a|3.99|2015-02-16 18:00:00|80.749667378538092|2|3260190085|190|35.464876580478958|0|3|561|-80.8438|64|35.23102|FR PROD ORGANIC PRODUCE|0.0|4|EBF ORG BABY LETTUCE 5 OZ|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00032601900854|FRESH PRODUCE|PRODUCE|-80.746334|80.746470557922436|205|1
35.41832|858c9713e934f5e6804a7971acc1bb373e35b243|4.99|2014-12-18 18:18:00|80.749667378538092|2|3338390203|190|35.464876580478958|0|3|561|-80.8438|64|35.23102|FR PROD ORGANIC PRODUCE|0.0|4|ORG CARROTS 5LB BAG|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00033383902036|FRESH PRODUCE|PRODUCE|-80.746334|80.746470557922436|205|1
35.41832|c4a307a54bfbcd8212b1a365e34a72514af4b013|3.79|2015-01-16 17:52:00|80.749667378538092|2|4138700530|190|35.464876580478958|0|3|209|-80.8438|20|35.23102|POWDERED SOFT DRINKS|0.0|1|4C LEMONADE LIQ WTR ENHNCR|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00041387005325|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.746334|80.746470557922436|205|1
35.41832|c05aed2b5d8b978677b68f25b31a7488780b48e8|2.55|2015-01-04 11:22:00|80.749667378538092|2|4156514116|190|35.464876580478958|0|3|1211|-80.8438|272|35.23102|HISP SALSA/DIPS|0.55|1|PACE REST SALSA MED|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00041565193882|HISPANIC PREP. FOODS|G1 GROCERY|-80.746334|80.746470557922436|205|1
35.41832|b52dc6d531402ca1e72a0c591fe57cd4872bc0be|4.19|2015-02-22 16:51:00|80.749667378538092|2|81088201002|190|35.464876711042834|0|3|882|-80.662946|178|35.412407|FROZEN NATURAL/ORGANIC|0.5|5|KIDFRESH CHEESY PIZZA|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00810882010055|FROZEN NATURAL/ORGANIC|FROZEN|-80.746334|80.746352221258178|68|1
35.41832|8885b03342f38ce63b77807658194cefa469f31c|2.19|2014-09-23 17:02:00|80.749667378538092|2|76857300210|190|35.464876711042834|0|3|544|-80.662946|64|35.412407|FRESH PRODUCE FRSH HERBS|0.2|4|PKG FRESH BAY LEAVES|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00768573002905|FRESH PRODUCE|PRODUCE|-80.746334|80.746352221258178|68|1
35.41832|d5f53367aa6b91e7c8f73c74c3dc5057d4fed7e1|19.98|2014-12-23 16:16:00|80.749667378538092|2|89991100046|190|35.464876711042834|0|3|9958|-80.662946|886|35.412407|NFS-PREM-OTHER WHITE|0.0|13|NEW AGE WHITE|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00899911000465|PREMIUM ($8-$10.99)|WINE|-80.746334|80.746352221258178|68|2
35.41832|4eea01f5521d547b432915ad8a4246af68c44f21|2.99|2014-10-04 10:59:00|80.749667378538092|2|1620033128|190|35.464876711042834|0|3|226|-80.662946|35|35.412407|SUGAR-POWDERED|0.0|1|DIXIE CRYSTAL 10X SUGAR BAG|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00016200331288|SUGAR/SUBSTITUTES|G1 GROCERY|-80.746334|80.746352221258178|68|1
35.41832|e50caaefade360073febd1ec23cf2541c0acf934|3.99|2014-11-17 18:05:00|80.749667378538092|2|7835470843|190|35.464876547546233|0|3|317|-80.844274|52|35.204336|CHUNK AND BAR CHEESE|1.49|3|CABOT 50% LIGHT CHEDDAR|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00078354707289|CHEESE|DAIRY|-80.746334|80.746486538521197|61|1
35.41832|b398bc2eb87e756ca8c20d3408cdd3ac3e9758c4|4.59|2015-01-31 15:15:00|80.749667378538092|2|7318000002|190|35.464876711042834|0|3|208|-80.662946|32|35.412407|NFS-COCKTAIL ACCESSORIES|0.0|1|SOODHALTER KING SIZE PICK|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00073180000023|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.746334|80.746352221258178|68|1
35.41832|244060f8ba933bdc0c8cf2820107f7a92df03b42|4.99|2014-11-18 15:24:00|80.749667378538092|2|7274500143|190|35.464876711042834|0|3|1226|-80.662946|107|35.412407|HEAT & EAT ENTREES|0.0|19|PERDUE DINO CHICKEN NUGGETS|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00072745001079|HEAT & EAT|CASE READY MEATS|-80.746334|80.746352221258178|68|1
35.41832|5fe2171d3b1be03e330343a0144e573e4a772414|3.59|2015-02-18 18:41:00|80.749667378538092|2|7357000008|190|35.464876580478958|0|3|317|-80.8438|52|35.23102|CHUNK AND BAR CHEESE|1.8|3|HELUVA GOOD COLBY JACK|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00073570000183|CHEESE|DAIRY|-80.746334|80.746470557922436|205|1
35.41832|317dbc58b8584a3c311685ebb760e806cc60fec8|3.98|2014-10-29 12:19:00|80.749667378538092|2|7203688096|190|35.464876711042834|0|3|526|-80.662946|64|35.412407|FRESH MUSHROOMS|0.4|4|HT SLICED WHITE MUSHROOMS|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00072036880963|FRESH PRODUCE|PRODUCE|-80.746334|80.746352221258178|68|2
35.41832|99f1e589767f826568fe91b81b2511c42877e839|3.99|2015-01-20 20:22:00|80.749667378538092|2|7203676057|190|35.464876580478958|0|3|1220|-80.8438|275|35.23102|PASTA SC PREMIUM|1.49|1|HT TRADER SAUCE TOM BASIL|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00072036760579|PASTA SAUCES|G1 GROCERY|-80.746334|80.746470557922436|205|1
35.41832|672b66a16e336b33cb02a8767a50503d2e9b2616|2.95|2014-12-24 08:46:00|80.749667378538092|2|7203663125|190|35.464876711042834|0|3|1262|-80.662946|57|35.412407|HALF N HALF WHIPPING CREAM|0.45|3|HT HEAVY WHIPPING CREAM|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00072036630988|MILK|DAIRY|-80.746334|80.746352221258178|68|1
35.41832|964a33c2d70d528993f8aa4f635697d633722c8f|3.25|2015-03-01 15:42:00|80.749667378538092|2|7203655010|190|35.464876580478958|0|3|317|-80.8438|52|35.23102|CHUNK AND BAR CHEESE|0.0|3|HT COLBY JACK CHEESE|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00072036705105|CHEESE|DAIRY|-80.746334|80.746470557922436|205|1
35.41832|de5b6d3423b46bf4cc507c34bd76367de5e276b8|6.55|2014-09-23 08:57:00|80.749667378538092|2|7570616502|190|35.464876546244774|0|3|254|-80.826724|892|35.195689|PREMIUM PIZZA|0.57|5|PALERMOS HT MEAT LOVERS PZZA|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00075706148073|FROZEN PIZZA|FROZEN|-80.746334|80.746487135802653|412|1
35.41832|c34593113ecf656b03efa14e79eca0f3052dbdb7|2.39|2014-09-27 16:09:00|80.749667378538092|2|4127102562|190|35.464876711042834|0|3|341|-80.662946|57|35.412407|CREAMERS|0.0|3|ITNAT'L AMARETTO CREAM|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00041271019667|MILK|DAIRY|-80.746334|80.746352221258178|68|1
35.41832|baf210eb846bdaec567cbca22e78c1e926c3e796|6.39|2014-12-09 16:22:00|80.749667378538092|2|4154800385|190|35.464876711042834|0|3|252|-80.662946|45|35.412407|PREMIUM ICE CREAM|1.61|5|EDY'S SLOW CHURNED CARAMEL D|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00041548345864|ICE CREAM|FROZEN|-80.746334|80.746352221258178|68|1
35.41832|7b5755c42e0d242f406b7ccd4c1aa3135e9a4b4f|0.95|2014-10-11 16:30:00|80.749667378538092|2|5210002123|190|35.464876711042834|0|3|80|-80.662946|34|35.412407|SEASONING PACKETS|0.0|1|MC FAJITAS MARINADE|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00052100021218|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.746334|80.746352221258178|68|1
35.41832|7bd1132bd3c8c304b3b1afcda5af04a8a39835e3|8.79|2014-10-19 10:08:00|80.749667378538092|2|9955508520|190|35.464876711042834|0|3|37|-80.662946|10|35.412407|PODS/CUPS/SINGLES|0.0|1|TULLY'S BREAKFAST BLEND K-CUPS|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00099555088007|COFFEE|G1 GROCERY|-80.746334|80.746352221258178|68|1
35.41832|4becb1ed9d6d98d212917233071b57455c0e3683|9.97|2015-01-13 14:17:00|80.749667378538092|2|20253500000|190|35.464876711042834|0|3|299|-80.662946|49|35.412407|ANGUS BEEF|0.0|2|ANGUS BEEF SIRLOIN STIR FRY|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00202533000001|BEEF|MEAT|-80.746334|80.746352221258178|68|2
35.41832|7e70c4f7343802198730548055f84c63190a566a|0.79|2014-12-06 18:54:00|80.749667378538092|2||190|35.464876580478958|0|3|532|-80.8438|64|35.23102|FRESH CUCUMBERS|0.0|4|COO CUCUMBERS S/S|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00204062000002|FRESH PRODUCE|PRODUCE|-80.746334|80.746470557922436|205|1
35.41832|ba02bb1532b4618b72beaee76a8c2c8b9a73fa6c|4.8|2014-11-09 12:20:00|80.749667378538092|2|20602200000|190|35.464876546244774|0|3|2018|-80.826724|505|35.195689|PRESSED CHEESE|1.6|6|YANCEYS JALAPENO&PEPPADEW (FC)|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00206022000008|SPECIALTY CHEESE|DELI|-80.746334|80.746487135802653|412|1
35.41832|81353111dc5312fe3bf2f82e728c67cd7055e7ad|1.98|2014-12-11 14:02:00|80.749667378538092|2|7339000780|190|35.464876711042834|0|3|48|-80.662946|7|35.412407|REGISTER GUM|0.0|1|MENTOS MINT ROLL 15CT|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00073390000110|CANDY|G1 GROCERY|-80.746334|80.746352221258178|68|2
35.41832|b2c7f10ee3407c78b5e5fd390fef6bbcc1d1e5f6|5.78|2014-10-22 16:34:00|80.749667378538092|2|7203695917|190|35.464876711042834|0|3|1625|-80.662946|373|35.412407|FROZEN DOUGH (ROLLS)|2.8|14|FRESH CHICAGO ROLL|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00072036959171|ROLLS|BAKERY|-80.746334|80.746352221258178|68|2
35.41832|41d7208ce61d4ff8bfa8ad5cf273416006bbd388|3.89|2014-12-03 18:24:00|80.749667378538092|2|8411410812|190|35.464876580478958|0|3|201|-80.8438|31|35.23102|POTATO CHIPS|1.39|1|KETTLE JALAPENO CHIPS|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00084114116321|SNACKS|G1 GROCERY|-80.746334|80.746470557922436|205|1
35.41832|ff7d50bd54c5bf6cd15dca913c2b58471ed67ec3|19.99|2015-01-30 12:21:00|80.749667378538092|2|7203695592|190|35.464876711042834|0|3|1653|-80.662946|381|35.412407|CELEBRATION CAKES|0.0|14|1/4 SHT DL MARBLE CAK  W/BUTCR|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00072036955920|CAKES|BAKERY|-80.746334|80.746352221258178|68|1
35.41832|ab0929e75ef7c34d88ebd9d5aab89d688b7b31b5|3.89|2014-09-29 13:40:00|80.749667378538092|2|7203695502|190|35.464876711042834|0|3|1693|-80.662946|385|35.412407|CROISSANTS|0.0|14|ARTISAN BUTTER CROISSANTS|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00072036955029|SWEET GOODS|BAKERY|-80.746334|80.746352221258178|68|1
35.41832|507d096989576dcc66162ccd7d93496e0b0a6847|2.99|2015-02-09 19:11:00|80.749667378538092|2|3338365583|190|35.464876580478958|0|3|522|-80.8438|64|35.23102|FRESH TOMATOES|1.5|4|SWEET GRAPE TOMATO (PINT)|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00072036880284|FRESH PRODUCE|PRODUCE|-80.746334|80.746470557922436|205|1
35.41832|d723f4181fe53a159ffae893fe6cd0507dbe5385|1.69|2014-11-09 18:28:00|80.749667378538092|2|7203688003|190|35.464876580478958|0|3|527|-80.8438|64|35.23102|FRESH CARROTS|0.19|4|HT BABY CARROTS 1LB BAG|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00072036880031|FRESH PRODUCE|PRODUCE|-80.746334|80.746470557922436|205|1
35.41832|df900753f4bf94f18bcd162a6e6704a4833235fe|2.69|2015-02-06 16:58:00|80.749667378538092|2|3100019601|190|35.464876711042834|0|3|1279|-80.662946|48|35.412407|SINGLE SERVE FLAVOR|0.3|5|KID CUISINE FUN  NUGGETS|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00031000196240|FROZEN MEALS|FROZEN|-80.746334|80.746352221258178|68|1
35.41832|691871944401fb3947de8013371dd0930fde5550|7.38|2014-10-13 19:21:00|80.749667378538092|2|2113150124|190|35.464876711042834|0|3|1279|-80.662946|48|35.412407|SINGLE SERVE FLAVOR|2.38|5|M CALLENDER CHICKEN POT PIE|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00021131501242|FROZEN MEALS|FROZEN|-80.746334|80.746352221258178|68|2
35.41832|eb0c96db9bbf8753020a2e847bda5fffede17f90|2.49|2014-11-04 10:27:00|80.749667378538092|2|7279900861|190|35.46487650500918|0|3|50|-80.85013|7|35.175855|PEG CANDY|0.0|1|WERTHER'S ORIG. S/F CANDIES|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00072799831400|CANDY|G1 GROCERY|-80.746334|80.74650498322184|218|1
35.41832|8665f302d6849cba49de858b713a2be03aa6733d|9.99|2015-02-11 19:56:00|80.749667378538092|2|7274580558|190|35.464876580478958|0|3|353|-80.8438|110|35.23102|FROZEN CASE MEAT|0.0|19|PERDUE SIMPLY SMART GRLD STRIP|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00072745805868|FROZEN CASE MEAT|CASE READY MEATS|-80.746334|80.746470557922436|205|1
35.41832|726d8ff82ca5431cc3990aea92f10adb9e37f101|0.3|2014-12-16 19:19:00|80.749667378538092|2||190|35.464876580478958|0|3|527|-80.8438|64|35.23102|FRESH CARROTS|0.0|4|COO CARROTS, BULK|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00204562000007|FRESH PRODUCE|PRODUCE|-80.746334|80.746470557922436|205|1
35.41832|8d81381e15cccbabcad40f51483328a6df913c63|0.11|2014-11-29 17:38:00|80.749667378538092|2||190|35.464876580478958|0|3|527|-80.8438|64|35.23102|FRESH CARROTS|0.0|4|COO CARROTS, BULK|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00204562000007|FRESH PRODUCE|PRODUCE|-80.746334|80.746470557922436|205|1
35.41832|1e722271e723b093f29a5c76f17fc041408eaa90|10.06|2015-01-10 11:03:00|80.749667378538092|2|20039000000|190|35.464876547546233|0|3|1801|-80.844274|400|35.204336|FFM TURKEY|1.12|6|HONEY SMOKED TURKEY BREAST|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00200397000007|FFM MEAT|DELI|-80.746334|80.746486538521197|61|2
35.41832|8716a46fe146ed7fd31ca927c709e15f8aa0fcf7|0.47|2015-01-18 12:55:00|80.749667378538092|2|7203608133|190|35.464876711042834|0|3|82|-80.662946|11|35.412407|VINEGAR|0.0|1|HT VINEGAR WHITE DISTILLED 16|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00072036081339|CONDIMENTS|G1 GROCERY|-80.746334|80.746352221258178|68|1
35.41832|cd76fe196781066c5636f50fdd2ae67f48cd81de|5.49|2014-12-11 17:35:00|80.749667378538092|2|7254506262|190|35.464876580478958|0|3|353|-80.8438|110|35.23102|FROZEN CASE MEAT|0.0|19|STEAK UMM STEAKS 9 OZ|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00072545062621|FROZEN CASE MEAT|CASE READY MEATS|-80.746334|80.746470557922436|205|1
35.41832|fa039e50d4e91dd0b849c0d1062d0155629d61e5|13.99|2014-11-02 12:07:00|80.749667378538092|2|7199031600|190|35.464876711042834|0|3|455|-80.662946|82|35.412407|DOMESTIC PREMIUM 12PK&>|0.0|16|COORS LIGHT 24PK 12OZ CAN|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00071990316006|DOMESTIC BEER|BEER|-80.746334|80.746352221258178|68|1
35.41832|dee328140706b029b0ab8a42c0155cd6c975cea9|2.99|2015-01-11 16:34:00|80.749667378538092|2||190|35.464876580478958|0|3|504|-80.8438|64|35.23102|FRESH BERRIES|0.0|4|BLUEBERRIES PINT|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00033383222356|FRESH PRODUCE|PRODUCE|-80.746334|80.746470557922436|205|1
35.41832|3783bd36807c77cc179c3c34917c846ff77f06d7|8.84|2014-12-07 11:00:00|80.749667378538092|2|20894700000|190|35.464876711042834|0|3|977|-80.662946|201|35.412407|FRESH HT CHICKEN|0.0|2|HT WHOLE CHICKEN|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00208947000002|POULTRY|MEAT|-80.746334|80.746352221258178|68|1
35.41832|a6ea7090e82989d4cbdc397d7919084db61becb3|3.49|2014-10-24 16:43:00|80.749667378538092|2|7146426040|190|35.464876486833511|0|3|577|-80.825175|136|35.152722|OTHER MERCH FR MSC JUICE|0.0|4|BOLTHOUSE PROTEIN PLUS COFFEE|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00071464016272|OTHER MERCHANDISE|PRODUCE|-80.746334|80.746512283520943|160|1
35.41832|f6b561de8b62839d7ef74bc8bb31280d07543936|8.0|2015-01-03 13:30:00|80.749667378538092|2|84115200732|190|35.464876711042834|0|3|1165|-80.662946|87|35.412407|NFS-FRESH CONSUMER BUNCH|0.0|9|BUNCH- 3/$12 DAISY BUNCHES|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00841152007321|FLORAL|FLORAL|-80.746334|80.746352221258178|68|2
35.41832|8363e2b11511d7fe5419046ab6ec754290f01574|3.99|2014-12-23 19:15:00|80.749667378538092|2|7203676057|190|35.464876580478958|0|3|1220|-80.8438|275|35.23102|PASTA SC PREMIUM|1.49|1|HT TRADER SAUCE MARINARA|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00072036760586|PASTA SAUCES|G1 GROCERY|-80.746334|80.746470557922436|205|1
35.41832|f718aff36a4568dc1674dd5948976373ee8f0bf4|3.19|2014-12-29 17:43:00|80.749667378538092|2|7203655010|190|35.464876580478958|0|3|317|-80.8438|52|35.23102|CHUNK AND BAR CHEESE|1.52|3|HT MILD CHEDDAR CHEESE|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00072036550101|CHEESE|DAIRY|-80.746334|80.746470557922436|205|1
35.41832|69789f656499ef3c56efa697c8f1610d8c5d16f9|3.69|2015-01-18 19:09:00|80.749667378538092|2|2016922150|190|35.464876546244774|0|3|494|-80.826724|107|35.195689|HEAT & EAT SIDES|0.0|19|SIMPLY PARMESAN POTATOES|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00020169221801|HEAT & EAT|CASE READY MEATS|-80.746334|80.746487135802653|412|1
35.41832|a98fff01ebe495696ee60d0cb3bcaa6713aeea64|1.55|2014-10-22 21:17:00|80.749667378538092|2|78616201000|190|35.464876580478958|0|3|31|-80.8438|4|35.23102|NON CARBONATED WATER|0.55|1|VIT WATER ZERO XXX|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00786162002969|BOTTLED WATER|G1 GROCERY|-80.746334|80.746470557922436|205|1
35.41832|d129fa9075f36de4be83db51c145d4311f15f3b8|0.79|2014-10-12 12:32:00|80.749667378538092|2||190|35.464876711042834|0|3|524|-80.662946|64|35.412407|FRESH PROD FRESH ONIONS|0.2|4|COO GREEN ONIONS|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00204068000006|FRESH PRODUCE|PRODUCE|-80.746334|80.746352221258178|68|1
35.41832|149855247ad4b22e25bb62d5c6e433ec2e30036b|3.19|2015-01-25 18:13:00|80.749667378538092|2|2100000730|190|35.464876580478958|0|3|316|-80.8438|52|35.23102|CREAM CHEESE|1.19|3|PHILLY SOFT CREAM CHEESE|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00021000000142|CHEESE|DAIRY|-80.746334|80.746470557922436|205|1
35.41832|ccbcd615b4251aac1742d34ae8efb066928f240f|3.67|2014-11-12 20:08:00|80.749667378538092|2|7203698628|190|35.464876580478958|0|3|284|-80.8438|892|35.23102|SUPER PREMIUM PIZZA|0.33|5|HTT MARGHERITA FLATBRD PIZZA|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00072036986313|FROZEN PIZZA|FROZEN|-80.746334|80.746470557922436|205|1
35.41832|6c61b4958d80cef88f0fa6dbedb884432b822922|3.75|2014-10-30 10:46:00|80.749667378538092|2|7203698557|190|35.464876580478958|0|3|424|-80.8438|72|35.23102|NFS-FACIAL TISSUE|0.25|1|HT FACIAL TISSUE|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00072036985576|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.746334|80.746470557922436|205|3
35.41832|a352b0de5588b02642dd5c990a2dee6685af51bd|7.78|2015-01-14 18:50:00|80.749667378538092|2|7192100989|190|35.464876580478958|0|3|284|-80.8438|892|35.23102|SUPER PREMIUM PIZZA|0.78|5|DIG FOR 1 TTRADITION CRUST PEP|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00071921008291|FROZEN PIZZA|FROZEN|-80.746334|80.746470557922436|205|2
35.41832|9a2cd37c3af84048d325df601a15d047b96f6862|2.99|2015-02-03 20:14:00|80.749667378538092|2|2100000028|190|35.464876580478958|0|3|316|-80.8438|52|35.23102|CREAM CHEESE|0.99|3|PHILLY LIGHT SOFT CRM CHEESE|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00021000000289|CHEESE|DAIRY|-80.746334|80.746470557922436|205|1
35.41832|e802982205d119545090419f8a1d96d7c7557b99|5.99|2014-10-14 18:49:00|80.749667378538092|2|2858800340|190|35.464876711042834|0|3|5846|-80.662946|1538|35.412407|KITCHEN GADGETS BARWARE|1.2|18|(JHK) WAITERS CORKSCREW|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00028588003404|KITCHEN GADGETS|GM|-80.746334|80.746352221258178|68|1
35.41832|67c4b5d1dbeb1d189d8db51326afd7112e511d32|12.99|2014-11-16 13:05:00|80.749667378538092|2|7023666311|190|35.464876711042834|0|3|751|-80.662946|87|35.412407|NFS-BOUQUETS|0.0|9|$12.99 SUNNY DAY BOUQUET|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00070236663119|FLORAL|FLORAL|-80.746334|80.746352221258178|68|1
35.41832|15568c84f9eda5ad470907fb247db4bc7645e6d3|1.34|2014-12-02 17:48:00|80.749667378538092|2|7047045916|190|35.464876580478958|0|3|685|-80.8438|61|35.23102|GREEK|0.0|3|YOPLAIT GREEK BLEND STWBRY RAS|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00070470459158|YOGURT|DAIRY|-80.746334|80.746470557922436|205|1
35.41832|31feade000773bceb4d62a6b12814fb4c436336d|4.58|2014-09-27 15:33:00|80.749667378538092|2|7800023046|190|35.46487650500918|0|3|55|-80.85013|8|35.175855|REGULAR|0.79|23|7-UP 2 LTR NR|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00078000000344|CARBONATED BEVERAGES|BEVERAGE|-80.746334|80.74650498322184|218|2
35.41832|525411f1163f465a5c8664bdb327026e5b965b5e|2.49|2015-01-30 14:33:00|80.749667378538092|2|7203659022|190|35.464876711042834|0|3|312|-80.662946|51|35.412407|BUTTER|0.0|3|HT BUTTR QTR 1/2S|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00072036590220|BUTTER & MARGARINE|DAIRY|-80.746334|80.746352221258178|68|1
35.41832|8853a2baa11ce5ec94209b44a77fb50080ffc734|4.85|2014-10-25 17:30:00|80.749667378538092|2|20182000000|190|35.464876711042834|0|3|655|-80.662946|49|35.412407|STR MDE VALUE ADDED BEEF|0.54|2|STKHOUSE MARNTD BEEF ON STICK|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00201820000007|BEEF|MEAT|-80.746334|80.746352221258178|68|1
35.41832|742f2caf654e7d3d840b26dd7b3a4224290dcfc4|3.89|2014-11-25 20:19:00|80.749667378538092|2|8411410812|190|35.464876580478958|0|3|201|-80.8438|31|35.23102|POTATO CHIPS|0.0|1|KETTLE BACKYARD BBQ CHIPS|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00084114113917|SNACKS|G1 GROCERY|-80.746334|80.746470557922436|205|1
35.41832|ad56bbdc2e068662689646a48f110ed01d615767|9.99|2014-10-30 18:56:00|80.749667378538092|2|8858600416|190|35.464876711042834|0|3|9956|-80.662946|886|35.412407|NFS-PREM-REISLING|0.0|13|CHT ST MICH HARV SEL RIESLING|13cab2c167627b85538b24000837f2ba6851f62d|3.2169564661626153|35.465179900649026|00088586004162|PREMIUM ($8-$10.99)|WINE|-80.746334|80.746352221258178|68|1
35.323246|136f52695cccabe53f239c29a48c053ea5e83ceb|8.99|2015-02-13 14:28:00|1.4102725052409182|2|7203695528|166|0.6165069451919168|0|1|1659|-80.945176|381|35.323246|VARIETY SINGLE LAYER|0.0|14|SGL LYR DBL FUDGE CAKE.|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00072036955289|CAKES|BAKERY|-80.945176|1.4127598348062935|166|1
35.323246|c4264eb5fae8a368adfeb5f1c0a40e276cfcfe74|8.99|2015-01-27 14:55:00|1.4102725052409182|2|7203695528|166|0.6165069451919168|0|1|1659|-80.945176|381|35.323246|VARIETY SINGLE LAYER|0.0|14|SGL LYR DBL FUDGE CAKE.|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00072036955289|CAKES|BAKERY|-80.945176|1.4127598348062935|166|1
35.323246|8a4ce22e0315ae5dd3239bb36521e2cd810ff2c2|8.99|2014-11-05 15:47:00|1.4102725052409182|2|7203695528|166|0.6165069451919168|0|1|1659|-80.945176|381|35.323246|VARIETY SINGLE LAYER|2.0|14|SGL LYR DBL FUDGE CAKE.|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00072036955289|CAKES|BAKERY|-80.945176|1.4127598348062935|166|1
35.323246|1ada93f770da4385cba791528b721b85798b3a62|8.99|2014-09-13 16:41:00|1.4102725052409182|2|7203695528|166|0.6165069451919168|0|1|1659|-80.945176|381|35.323246|VARIETY SINGLE LAYER|0.0|14|SGL LYR DBL FUDGE CAKE.|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00072036955289|CAKES|BAKERY|-80.945176|1.4127598348062935|166|1
35.323246|6194fd23ab0e297472c0c4651f0f3a86947cae88|8.99|2014-11-10 15:30:00|1.4102725052409182|2|7203695528|166|0.6165069451919168|0|1|1659|-80.945176|381|35.323246|VARIETY SINGLE LAYER|2.0|14|SGL LYR DBL FUDGE CAKE.|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00072036955289|CAKES|BAKERY|-80.945176|1.4127598348062935|166|1
35.323246|09c78dacc57f259ca0b625dc476ef50b9d58f2cf|8.99|2014-10-11 14:03:00|1.4102725052409182|2|7203695528|166|0.6165069451919168|0|1|1659|-80.945176|381|35.323246|VARIETY SINGLE LAYER|0.0|14|SGL LYR DBL FUDGE CAKE.|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00072036955289|CAKES|BAKERY|-80.945176|1.4127598348062935|166|1
35.323246|841ff4906ea49667f0140f841da250d243b01566|1.25|2015-01-02 15:14:00|1.4102725052409182|2|7203698557|166|0.6165069451919168|0|1|424|-80.945176|72|35.323246|NFS-FACIAL TISSUE|0.25|1|HT FACIAL TISSUE LOTION|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00072036985583|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|1b3e0e49c430ed0e0cf7c9fbea61017f3c63737d|4.49|2014-09-23 12:02:00|1.4102725052409182|2|7410855526|166|0.6165069451919168|0|1|3677|-80.945176|1060|35.323246|HAIR HAIRNETS|0.0|17|CNR HAIR NETS 10PK MEDIUM|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00074108555267|HAIR CARE ACCESSORIES|HBC|-80.945176|1.4127598348062935|166|1
35.323246|8c750d566b10106bf8c1059edd82431d89a9e903|5.69|2014-09-20 14:42:00|1.4102725052409182|2|7756725423|166|0.6165069451919168|0|1|252|-80.945176|45|35.323246|PREMIUM ICE CREAM|2.85|5|BREYERS CHERRY/VANILLA  I/C|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00077567254276|ICE CREAM|FROZEN|-80.945176|1.4127598348062935|166|1
35.323246|c69f0393c7e6f16a809565fe27859b1262854f82|6.99|2014-10-30 18:04:00|1.4102725052409182|2|20219900000|166|0.6165069451919168|0|1|299|-80.945176|49|35.323246|ANGUS BEEF|0.71|2|ANGUS SIRLOIN FILET CUSTOM CUT|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00202242000002|BEEF|MEAT|-80.945176|1.4127598348062935|166|1
35.323246|6439ccca16808e435680657af868c6c939a4ace0|13.99|2014-11-22 11:55:00|1.4102725052409182|2|7675304456|166|0.6165069451919168|0|1|5813|-80.945176|1534|35.323246|METAL BAKEWARE (TINWARE)|7.0|18|CER BAKEWARE RECT 1.0 CT|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00076753044561|MEATAL/GLASS BAKEWARE|GM|-80.945176|1.4127598348062935|166|1
35.323246|019b495d1ffb4454bb66d24b89a29043a5d83ee6|1.3|2014-10-05 16:35:00|1.4102725052409182|2|5000000124|166|0.6165069451919168|0|1|154|-80.945176|24|35.323246|NFS-CAT FOOD WET|0.3|1|FANCY FEAST GRAVY LOVERS TURKY|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00050000580040|PET FOOD/SUPPLIES|G1 GROCERY|-80.945176|1.4127598348062935|166|2
35.323246|00286305f7d90fbbfa760b1a41ff4e853cc05c72|1.3|2014-10-03 16:48:00|1.4102725052409182|2|5000000124|166|0.6165069451919168|0|1|154|-80.945176|24|35.323246|NFS-CAT FOOD WET|0.3|1|FANCY FEAST GRAVY LOVERS TURKY|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00050000580040|PET FOOD/SUPPLIES|G1 GROCERY|-80.945176|1.4127598348062935|166|2
35.323246|a1d0a608c308d8fead17c21d710c97997b4ce87d|2.38|2015-02-14 11:19:00|1.4102725052409182|2|3940001747|166|0.6165069451919168|0|1|242|-80.945176|39|35.323246|CANNED BEANS|0.38|1|BUSH BEAN GARBANZOS|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00039400017004|VEGETABLES-CAN/JAR|G1 GROCERY|-80.945176|1.4127598348062935|166|2
35.323246|549edc45c1a34a3a7a1904783e4faad2f9d112f9|6.58|2014-12-12 15:31:00|1.4102725052409182|2|4144930140|166|0.6165069451919168|0|1|9|-80.945176|2|35.323246|DESSERT MIXES|1.65|1|KRUSTEAZ KEY LIME PIE|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00041449107929|BAKING MIXES|G1 GROCERY|-80.945176|1.4127598348062935|166|2
35.323246|3c2cdac8e8192353a8cf9d015bd2b9de2245089d|9.99|2015-02-28 15:53:00|1.4102725052409182|2|7987930192|166|0.6165069451919168|0|1|1687|-80.945176|385|35.323246|THAW & SELL (SWEET GOODS)|0.0|14|GLUTEN FREE CHOC CAKE|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00079879301921|SWEET GOODS|BAKERY|-80.945176|1.4127598348062935|166|1
35.323246|0a20dbf9d79f11c76d44ee5a3038b7321ce2d88f|9.99|2015-03-08 14:22:00|1.4102725052409182|2|7987930192|166|0.6165069451919168|0|1|1687|-80.945176|385|35.323246|THAW & SELL (SWEET GOODS)|0.0|14|GLUTEN FREE CHOC CAKE|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00079879301921|SWEET GOODS|BAKERY|-80.945176|1.4127598348062935|166|1
35.323246|4401f88b8fc23b3e594b1e7fadffe154db1cfe18|2.99|2014-11-24 15:36:00|1.4102725052409182|2|7231000145|166|0.6165069451919168|0|1|235|-80.945176|37|35.323246|GREEN TEA|1.5|1|BIGELOW TEA GREEN DECAF|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00072310042476|TEA|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|202cf5ae4d10298a4d606db8dec4b72913498c9b|6.11|2014-09-25 19:37:00|1.4102725052409182|2|27082900000|166|0.6165069451919168|0|1|973|-80.945176|201|35.323246|FRESH PERDUE CHICKEN|2.04|2|PERDUE BNLS CHICKEN BREAST|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00270829000004|POULTRY|MEAT|-80.945176|1.4127598348062935|166|1
35.323246|018e3fa40f984827b088a2f88fdc860465416095|1.0|2014-12-22 11:45:00|1.4102725052409182|2||166|0.6165069451919168|0|1|509|-80.945176|64|35.323246|FRESH CITRUS-REMAINING|0.0|4|COO LIMES, LRG|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00204048000002|FRESH PRODUCE|PRODUCE|-80.945176|1.4127598348062935|166|2
35.323246|37b87adfa3da959c2fba18f9048e230186bb7fdc|5.99|2014-12-20 11:22:00|1.4102725052409182|2|7756725423|166|0.6165069451919168|0|1|275|-80.945176|45|35.323246|SUPER PREMIUM ICE CREAM|3.0|5|BREYERS SALTED CARAMEL|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00077567254450|ICE CREAM|FROZEN|-80.945176|1.4127598348062935|166|1
35.323246|c51da777accbd1de4759d0de86a41e71932b35d9|5.99|2015-01-20 14:38:00|1.4102725052409182|2|7756725423|166|0.6165069451919168|0|1|275|-80.945176|45|35.323246|SUPER PREMIUM ICE CREAM|2.99|5|BREYERS SALTED CARAMEL|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00077567254450|ICE CREAM|FROZEN|-80.945176|1.4127598348062935|166|1
35.323246|d68a40080f24819c37e97cdede492d4d35bb2d12|3.89|2015-01-24 14:47:00|1.4102725052409182|2|1300000466|166|0.6165069451919168|0|1|70|-80.945176|11|35.323246|KETCHUP|1.39|1|HEINZ KETCHUP 38 OZ|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00013000004664|CONDIMENTS|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|2892e0ffbe903466b7fd8e8883a79c7cf6d16a13|8.99|2014-12-06 16:00:00|1.4102725052409182|2|89402970258|166|0.6165069451919168|0|1|7305|-80.945176|1600|35.323246|CHRISTMAS INDOOR DECOR IMP|3.0|18|"I/O 6"" BO CRYSTAL TREE"|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00894029702584|SEASONAL MERCHANDISE|GM|-80.945176|1.4127598348062935|166|1
35.323246|7a70b17556095b13767eb80181366ae6355586ac|3.19|2014-11-15 10:32:00|1.4102725052409182|2|1920081145|166|0.6165069451919168|0|1|399|-80.945176|69|35.323246|NFS-DISINFECTANTS|0.0|1|LYSOL WIPES POWER & FREE|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00019200880695|HOUSEHOLD CLEANERS/SUPPLIES|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|0b6a4d937651cfb0143a704366a58d25bd681416|0.88|2014-10-17 19:23:00|1.4102725052409182|2||166|0.6165069451919168|0|1|502|-80.945176|64|35.323246|FRESH BANANAS|0.0|4|BANANAS, YELLOW|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.945176|1.4127598348062935|166|1
35.323246|081894f790a4086afd6a823de7bf1ce3a4cdd6f3|5.99|2014-12-24 14:50:00|1.4102725052409182|2|1328632126|166|0.6165069451919168|0|1|7419|-80.945176|1600|35.323246|CHRISTMAS GIFT WRAP|2.0|18|"I/O 40"" JUVENLE CMAS WRAP 90SF"|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00013286321257|SEASONAL MERCHANDISE|GM|-80.945176|1.4127598348062935|166|1
35.323246|2fd277641f2123759a4e6388646cd7df84f34741|7.99|2014-10-21 13:42:00|1.4102725052409182|2|71981286251|166|0.6165069451919168|0|1|5939|-80.945176|1538|35.323246|UTENSILS-COOKING METAL|0.0|18|(JHK) OXO POTATO MASHER|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00719812862514|KITCHEN GADGETS|GM|-80.945176|1.4127598348062935|166|1
35.323246|748eac033d148ca7026d51f21e29688936c0ab6e|1.0|2015-01-13 11:46:00|1.4102725052409182|2||166|0.6165069451919168|0|1|522|-80.945176|64|35.323246|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00204664000004|FRESH PRODUCE|PRODUCE|-80.945176|1.4127598348062935|166|1
35.323246|a0e59663dd41fde660b64381226f521fdef5527a|5.99|2015-01-16 12:01:00|1.4102725052409182|2|7756725423|166|0.6165069451919168|0|1|275|-80.945176|45|35.323246|SUPER PREMIUM ICE CREAM|3.0|5|BREYERS BLK RASPBERRY CHOC|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00077567264794|ICE CREAM|FROZEN|-80.945176|1.4127598348062935|166|1
35.323246|338c81db30114d1ff968fcd2c2eec9e6257ec2c7|8.99|2014-12-31 15:42:00|1.4102725052409182|2|7675304010|166|0.6165069451919168|0|1|5813|-80.945176|1534|35.323246|METAL BAKEWARE (TINWARE)|0.9|18|GC NS BAKE & ROAST PAN 13X9|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00076753040105|MEATAL/GLASS BAKEWARE|GM|-80.945176|1.4127598348062935|166|1
35.323246|aff66eb4acc508291366b5db544df580bb8d08e5|5.16|2015-01-10 12:34:00|1.4102725052409182|2|3940001810|166|0.6165069451919168|0|1|242|-80.945176|39|35.323246|CANNED BEANS|1.16|1|BUSH PEAS BLACKEYE|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00039400013686|VEGETABLES-CAN/JAR|G1 GROCERY|-80.945176|1.4127598348062935|166|4
35.323246|bfd616df429d61b440bbb114735250166369ab9c|2.69|2014-11-28 14:53:00|1.4102725052409182|2|1600026460|166|0.6165069451919168|0|1|42|-80.945176|6|35.323246|GRANOLA/YOGURT BARS|0.0|1|NV BAR GF CRN ALMND RST NUT|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00016000146228|BREAKFAST FOODS|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|3468942ab25d26673b3b1267b4c143c1a74d154d|10.0|2015-01-29 10:49:00|1.4102725052409182|2|20229500000|166|0.6165069451919168|0|1|299|-80.945176|49|35.323246|ANGUS BEEF|0.0|2|ANGUS BEEF EYE OF ROUND ROAST|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00202295000004|BEEF|MEAT|-80.945176|1.4127598348062935|166|1
35.323246|299def4f3d568270f9eaf244e4ed5651a216d561|2.97|2014-11-26 14:23:00|80.945255278477163|2||166|35.350513409356338|0|13|523|-80.85013|64|35.175855|FRESH POTATOES|1.82|4|COO SWEET POTATOES, BULK|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|35.37387923947206|00204091000004|FRESH PRODUCE|PRODUCE|-80.945176|80.945212806973615|218|1
35.323246|083f98b209ca8a3b02c1c0a3eff45eee73579974|6.39|2014-12-30 15:10:00|1.4102725052409182|2|4480075010|166|0.6165069451919168|0|1|223|-80.945176|35|35.323246|SUGAR SUBSTITUTES|1.0|1|STEVIA EXTRACT IN THE RAW|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00044800750109|SUGAR/SUBSTITUTES|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|2ebff347276a2439f36b96064dfc39af790c24cf|3.69|2014-12-12 15:35:00|1.4102725052409182|2|4178000159|166|0.6165069451919168|0|1|201|-80.945176|31|35.323246|POTATO CHIPS|0.9|1|UTZ RF KETTLE CHIPS|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00041780001207|SNACKS|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|33735ea1558f5646c0529425e84d17bb4248244f|2.99|2015-02-26 12:22:00|1.4102725052409182|2|3120020007|166|0.6165069451919168|0|1|130|-80.945176|20|35.323246|CRANBERRY JUICE/DRINKS-SHELF|0.0|1|OSPRAY CRANBERRY JUICE|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00031200200075|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.323246|626d61a9c61b955fc97ec924e6a28ea0aaa64840|2.29|2015-01-04 14:04:00|1.4102725052409182|2|7203663996|166|0.6165069451919168|0|1|342|-80.945176|57|35.323246|FRESH MILK|0.82|3|HARRIS TEETER FF SKIM MILK|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00072036631299|MILK|DAIRY|-80.945176|1.4127598348062935|166|1
35.323246|e934499fc78a4d101e3b4dd120791d724509f507|2.29|2015-01-09 17:24:00|1.4102725052409182|2|4133533217|166|0.6165069451919168|0|1|184|-80.945176|28|35.323246|SALAD DRESSINGS-LIQUID|1.29|1|KENS DRS LO RANCH|206a4fd6bbee51152375fbba011e5d6a84a3179c|1.8841132803857976|0.61833652052202714|00041335000419|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.945176|1.4127598348062935|166|1
35.000049|a69d5e0a225e609732d2a902f226d0ac81059b44|3.75|2015-02-15 13:42:00|80.700248323638462|2|4139000107|249|35.103207963171322|0|7|79|-80.7007|273|35.06858|ASIAN SAUCES/SEASONINGS|0.0|1|KIKKOMAN SOY SAUCE LT 15|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00041390001079|ASIAN PREP. FOODS|G1 GROCERY|-80.699686|80.699775519439697|273|1
35.000049|1bfc65d0e070a2e041c9802f9b553f348681d013|2.49|2015-02-17 14:43:00|80.700248323638462|2|5040073942|249|35.103207963171322|0|7|1033|-80.7007|163|35.06858|HAMBURGER|0.0|7|BALL PARK WHITE HAMS 8PK PP|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00050400739420|BUNS/ROLLS|COMMERCIAL BAKERY|-80.699686|80.699775519439697|273|1
35.000049|84c2cb1196f9d192add77e5b6b632d3488174a33|3.49|2014-10-11 15:23:00|80.700248323638462|2|2733100023|249|35.103207963171322|0|7|495|-80.7007|108|35.06858|NON REFRIGERATED|0.0|19|LA BANDERITA L/CARB TORTILLAS|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00027331000233|TORTILLAS|CASE READY MEATS|-80.699686|80.699775519439697|273|1
35.000049|0f723e1d00a6c542733b4758cb262e7fd5128c29|3.35|2014-12-21 11:53:00|80.700248323638462|2|2840005597|249|35.10320798645877|0|7|199|-80.770346|31|35.052812|DIPS & SALSAS|0.35|1|TOSTITOS RESTRNT  STYLE SALSA|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00028400089364|SNACKS|G1 GROCERY|-80.699686|80.699715058480123|40|1
35.000049|679e1efb47360968a42e535e6a52cdbefbf4c897|3.65|2015-02-18 16:31:00|80.700248323638462|2|3010001610|249|35.103207962963474|0|7|1254|-80.732725|12|35.082768|FUDGE ENROBED|1.65|1|FUDGE SHOPPE GRASSHOPPER MINT|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00030100440574|COOKIES|G1 GROCERY|-80.699686|80.699775876128598|147|1
35.000049|31981cc297cd50bff5af50a34cb11a312e6bdc0a|3.29|2015-02-02 16:46:00|80.700248323638462|2|2840011895|249|35.103207963171322|0|7|204|-80.7007|31|35.06858|TORTILLA CHIPS|0.79|1|TOSTITOSTHIN & CRISPY|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00028400116886|SNACKS|G1 GROCERY|-80.699686|80.699775519439697|273|1
35.000049|b72dca64bed245168158f7c423b8be67a7ee2139|3.89|2014-09-17 17:07:00|80.700248323638462|2|3010001610|249|35.103207982226124|0|7|1254|-80.771677|12|35.066546|FUDGE ENROBED|1.39|1|FUDGE SHOPPE GRASSHOPPER MINT|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00030100440574|COOKIES|G1 GROCERY|-80.699686|80.69973234078671|45|1
35.000049|b2a167fe176e7f5163dbf66463121314859b1e35|2.19|2015-01-30 18:30:00|80.700248323638462|2|7203676220|249|35.103207963171322|0|7|886|-80.7007|150|35.06858|SAUCES|0.2|12|HT FISHERMANS COCKTAIL SAUCE.|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00072036762207|CONDIMENTS|SEAFOOD|-80.699686|80.699775519439697|273|1
35.000049|fba205d89129912ad09fa6437c3a957f76f0d53c|1.67|2014-09-13 12:46:00|1.4091206135396188|2|7203657031|249|0.6108660934093487|0|47|322|-80.699686|53|35.000049|SOUR CREAM|0.0|3|HT LIGHT SOUR CREAM|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|0.61242566243833529|00072036590343|CULTURES|DAIRY|-80.699686|1.4084752260255726|249|1
35.000049|734cb7afec4532fac560739dc3f5e094cd47adf5|1.99|2014-12-17 18:01:00|80.700248323638462|2|7203688096|249|35.103207963171322|0|7|526|-80.7007|64|35.06858|FRESH MUSHROOMS|0.1|4|HT SLICED WHITE MUSHROOMS|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00072036880963|FRESH PRODUCE|PRODUCE|-80.699686|80.699775519439697|273|1
35.000049|88b0fd062a7825ff60278ceef36c3d352c6841da|3.79|2014-11-17 18:06:00|80.700248323638462|2|7203688014|249|35.103207963171322|0|7|581|-80.7007|136|35.06858|FRESH SALSA|0.0|4|HT FRESH MILD SALSA|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00072036880215|OTHER MERCHANDISE|PRODUCE|-80.699686|80.699775519439697|273|1
35.000049|800657a9939e1278b9f67940f97d759d632235c9|3.79|2014-09-27 16:12:00|80.700248323638462|2|7203688014|249|35.103207962123129|0|7|581|-80.64817|136|35.04711|FRESH SALSA|0.0|4|HT FRESH MILD SALSA|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00072036880215|OTHER MERCHANDISE|PRODUCE|-80.699686|80.699777304047657|129|1
35.000049|18f2607ad79c64b949a8942aa68c2341ac3c3846|10.29|2015-01-05 16:52:00|80.700248323638462|2|20196400000|249|35.103207963171322|0|7|299|-80.7007|49|35.06858|ANGUS BEEF|0.0|2|HT RESERVE ANGUS SHAVED STK|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00201964000000|BEEF|MEAT|-80.699686|80.699775519439697|273|1
35.000049|2867deefa83b568f01b0c9886d4d7a6cda6efad7|2.0|2014-10-19 16:56:00|80.700248323638462|2|7464100079|249|35.103207963171322|0|7|562|-80.7007|64|35.06858|FRESH CUT FRUIT|0.0|4|APPLE CHEESE & CARMEL DIP|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00074641000798|FRESH PRODUCE|PRODUCE|-80.699686|80.699775519439697|273|1
35.000049|c749a4ca2a1502cc479ab7e0529319a619355212|2.5|2014-10-11 16:34:00|80.700248323638462|2|7774523089|249|35.103207963171322|0|7|563|-80.7007|64|35.06858|FRESH VEGETABLE/FRUIT TRAYS|0.0|4|R.P. APPLE/YOGURT/GRANOLA|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00077745230894|FRESH PRODUCE|PRODUCE|-80.699686|80.699775519439697|273|1
35.000049|0385709b71f16608f4f8b6f77a86b26ed231ec62|4.0|2015-03-02 17:24:00|80.700248323638462|2|7464100079|249|35.103207989172532|0|7|562|-80.760919|64|35.024332|FRESH CUT FRUIT|0.0|4|APPLE CHEESE & CARMEL DIP|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00074641000798|FRESH PRODUCE|PRODUCE|-80.699686|80.699688988614966|343|2
35.000049|2d74f25d1ed18912a0f9fb7cece47527f988e57d|0.81|2015-02-11 17:37:00|80.700248323638462|2||249|35.103207963171322|0|7|502|-80.7007|64|35.06858|FRESH BANANAS|0.0|4|BANANAS, YELLOW|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00204011000008|FRESH PRODUCE|PRODUCE|-80.699686|80.699775519439697|273|1
35.000049|3d1e3f8e8cd9c46993e4aa7dd4286586f5d09a34|4.49|2014-11-02 15:21:00|80.700248323638462|2|2531742000|249|35.103207963171322|0|7|659|-80.7007|103|35.06858|CHILDRENS LUNCH SNACKS|0.99|19|APPLEGATE HALF TIME TURK/CHSE|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00025317420006|LUNCH SNACKS|CASE READY MEATS|-80.699686|80.699775519439697|273|1
35.000049|49a1282f84b5bf42ae0f2f012826b3c7c1e04c3b|1.79|2015-03-09 19:32:00|80.700248323638462|2|2430004101|249|35.103207962123129|0|7|1044|-80.64817|173|35.04711|SW BAKD GOOD SNACK CAKES|0.0|7|LD HONEY BUNS|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00024300041020|SWEET BAKED GOODS|COMMERCIAL BAKERY|-80.699686|80.699777304047657|129|1
35.000049|f8184d623aa6a42c97950f7aa485a47183054333|4.29|2015-01-03 10:23:00|80.700248323638462|2|2840016014|249|35.103207963171322|0|7|201|-80.7007|31|35.06858|POTATO CHIPS|2.14|1|LAYS BBQ|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00028400160131|SNACKS|G1 GROCERY|-80.699686|80.699775519439697|273|1
35.000049|7e922d67c6e04eeee53f8c9fc75b4b134c4284b4|3.35|2015-02-22 14:19:00|80.700248323638462|2|1312000286|249|35.103207963171322|0|7|1469|-80.7007|278|35.06858|REGULAR CUT FRIES|0.0|5|ORE-IDA SHOESTRINGS|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00013120008283|FROZEN POTATO|FROZEN|-80.699686|80.699775519439697|273|1
35.000049|526fa73ea7ed0e3efe63d11991c4b57bf150e852|10.99|2014-10-23 17:18:00|80.700248323638462|2|83238600506|249|35.103207963171322|0|7|5734|-80.7007|1524|35.06858|TUMBLERS & DRINKWARE|0.0|18|VULCANO TRAVEL TUMBLER 16 OZ|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00832386005061|TUMBLERS|GM|-80.699686|80.699775519439697|273|1
35.000049|2f0366928cf4c5b3555a178d9f45ef8c00796a12|1.89|2014-12-31 16:21:00|80.700248323638462|2|73639310343|249|35.103207963171322|0|7|247|-80.7007|39|35.06858|VEGETABLES-FLANKER|0.64|1|GLORY TURKEY SND COLLARD GREEN|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00736393103232|VEGETABLES-CAN/JAR|G1 GROCERY|-80.699686|80.699775519439697|273|1
35.000049|76e47ef3f7e27f360984a0349f59380622ebc9c3|20.99|2014-12-06 17:51:00|80.700248323638462|2|20903500000|249|35.103207963171322|0|7|660|-80.7007|154|35.06858|FISH FILLETS WILD CGHT|7.35|12|WC FRESH YELLOWFIN TUNA ST (EC|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00209035000003|FISH FILLETS/STEAKS|SEAFOOD|-80.699686|80.699775519439697|273|1
35.000049|ea435c047491ff3ce0ead77fdf857dc3302dd99c|3.79|2014-11-04 17:16:00|80.700248323638462|2|1410007105|249|35.103207963171322|0|7|1025|-80.7007|162|35.06858|WHITE|0.0|7|PEP VERY THIN WHITE BRD PP|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00014100071051|SLICED BREAD|COMMERCIAL BAKERY|-80.699686|80.699775519439697|273|1
35.000049|b79d46ea58f2c4b62ffd5017bcf4f585f48a5fe6|6.79|2014-11-12 18:29:00|80.700248323638462|2|7800008216|249|35.103207963171322|0|7|54|-80.7007|8|35.06858|DIET|6.79|23|DT CHERRY DR PEPPER 12PK|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00078000099164|CARBONATED BEVERAGES|BEVERAGE|-80.699686|80.699775519439697|273|1
35.000049|683c7fd67283b26bdfb5dfa6faf8292a85807322|3.9|2015-02-09 13:36:00|80.700248323638462|2|20337400000|249|35.103207961024793|0|7|641|-80.758228|137|34.95459|PREMIUM PORK|0.0|2|PORK LOIN BNLS BUTTERFLY CHOPS|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00203382000006|PORK|MEAT|-80.699686|80.699779137358519|182|1
35.000049|3c709f04b5fe3bd2558cd495e7db264cec7a746c|1.2|2014-10-05 16:12:00|80.700248323638462|2||249|35.103207963171322|0|7|531|-80.7007|64|35.06858|FRESH CORN|0.0|4|COO YELLOW CORN|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00204078000003|FRESH PRODUCE|PRODUCE|-80.699686|80.699775519439697|273|2
35.000049|10a5c4147869caf84e5c0cfafa80e79608346523|13.58|2015-01-27 16:46:00|80.700248323638462|2|1200080994|249|35.103207963171322|0|7|54|-80.7007|8|35.06858|DIET|3.39|23|DT WILD CHERRY PEPSI FM|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00012000810176|CARBONATED BEVERAGES|BEVERAGE|-80.699686|80.699775519439697|273|2
35.000049|263253c319549ce73b4f8d5830608a2c24eb76bc|6.49|2014-10-09 08:12:00|80.700248323638462|2|1200080994|249|35.103207963171322|0|7|54|-80.7007|8|35.06858|DIET|1.5|23|DT WILD CHERRY PEPSI FM|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00012000810176|CARBONATED BEVERAGES|BEVERAGE|-80.699686|80.699775519439697|273|1
35.000049|f04380818688d956328020ee6504414ec1546067|2.29|2015-01-08 19:23:00|80.700248323638462|2|7800023046|249|35.103207873564727|0|7|55|-80.654118|8|35.123768|REGULAR|0.79|23|CHERRY 7 UP 2LTR NR|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00078000005318|CARBONATED BEVERAGES|BEVERAGE|-80.699686|80.699874680220944|473|1
35.000049|a02cb4697db897da7b829fbbe106327cd8a7794c|3.39|2014-12-23 19:15:00|80.700248323638462|2|5000012734|249|35.103207962963474|0|7|341|-80.732725|57|35.082768|CREAMERS|0.89|3|COFFEEMATE SF ITALIAN SWT CRM|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00050000145782|MILK|DAIRY|-80.699686|80.699775876128598|147|1
35.000049|d54c5834716f3852080fc619dcc06c19b1179e38|2.85|2014-11-14 17:33:00|80.700248323638462|2|8390000536|249|35.103207963171322|0|7|365|-80.7007|56|35.06858|REFRIGERATED TEAS|0.85|3|GOLD PEAK DIET TEA|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00083900005382|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.699686|80.699775519439697|273|1
35.000049|cce26b2cc6a90984dbe8f9b112e04df4ba40f1bb|2.85|2014-11-01 11:53:00|80.700248323638462|2|8390000536|249|35.103207963171322|0|7|365|-80.7007|56|35.06858|REFRIGERATED TEAS|0.85|3|GOLD PEAK DIET TEA|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00083900005382|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.699686|80.699775519439697|273|1
35.000049|c07ce49bd01601ad25f8e8fbe5960120e5e8b4d9|2.99|2014-09-18 08:10:00|80.700248323638462|2|61126962373|249|35.103207963171322|0|7|97|-80.7007|8|35.06858|ENERGY DRINKS|0.0|23|RED BULL TOTAL ZERO 12 OZ|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00611269623734|CARBONATED BEVERAGES|BEVERAGE|-80.699686|80.699775519439697|273|1
35.000049|8b7e0abebf891bdf0a31287ae033aa4b0f91473d|3.99|2014-09-24 16:56:00|80.700248323638462|2|5783602064|249|35.10320798645877|0|7|522|-80.770346|64|35.052812|FRESH TOMATOES|0.0|4|CAMPARI TOMATO 16 OZ|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00057836020641|FRESH PRODUCE|PRODUCE|-80.699686|80.699715058480123|40|1
35.000049|eaac9f292b66982737d8b29c4db9945fb6d584f0|2.29|2014-11-11 13:16:00|80.700248323638462|2|7357013000|249|35.103207963171322|0|7|1267|-80.7007|53|35.06858|DIPS AND SPREADS|0.0|3|HELUVA GOOD FRENCH ONION DIP|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00073570130002|CULTURES|DAIRY|-80.699686|80.699775519439697|273|1
35.000049|ab9a4c2db9b9b43db541f3309a4a26128adde004|6.87|2014-11-20 08:23:00|80.700248323638462|2|61126999100|249|35.103207963171322|0|7|97|-80.7007|8|35.06858|ENERGY DRINKS|1.87|23|RED BULL TOTAL ZERO 8.4 OZ|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00611269623727|CARBONATED BEVERAGES|BEVERAGE|-80.699686|80.699775519439697|273|3
35.000049|2cba3a113f8f2475a229cd91dd6eedc54abcfbeb|3.99|2015-01-22 16:54:00|1.4091206135396188|2|4525511880|249|0.6108660934093487|0|47|523|-80.699686|64|35.000049|FRESH POTATOES|0.0|4|DUTCH YELLOW POTATO 24 OZ|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|0.61242566243833529|00045255118803|FRESH PRODUCE|PRODUCE|-80.699686|1.4084752260255726|249|1
35.000049|3d8d71a589f47a2f7d3ab49fa19aea44ebf0c08e|4.49|2015-01-14 16:45:00|80.700248323638462|2|3663202782|249|35.103207963171322|0|7|685|-80.7007|61|35.06858|GREEK|0.99|3|DANNON OIKOS VANILLA 4 PK|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00036632027825|YOGURT|DAIRY|-80.699686|80.699775519439697|273|1
35.000049|e746409558bc96e50b9f8fa0c6e237d8d7de6fc5|5.69|2014-10-01 18:11:00|80.700248323638462|2|3680036723|249|35.103207873564727|0|7|4236|-80.654118|1200|35.123768|DEX ADULT/CHILDREN|0.0|17|TC DAYTIME PE ORIGINAL LIQ|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00036800367326|COUGH/COLD/SINUS|HBC|-80.699686|80.699874680220944|473|1
35.000049|560b305a85c54c089656d8a12411dfd7102373e0|1.69|2014-12-12 18:35:00|80.700248323638462|2|4178900621|249|35.103207963171322|0|7|1203|-80.7007|33|35.06858|RAMEN|0.69|1|MARUCHAN RAMEN CHICKEN 6PK|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00041789006210|SOUP|G1 GROCERY|-80.699686|80.699775519439697|273|1
35.000049|927e1268c0a26eb7508c5b54714618f5db0520ac|19.98|2014-10-22 17:44:00|80.700248323638462|2|64365400136|249|35.103207989166933|0|7|9945|-80.699909|885|35.002628|NFS POP OTHER WHITE|0.0|13|HINNANT CAROLINA WILDFLOWER|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00643654001360|POPULAR (4-$7.99)|WINE|-80.699686|80.699689264455898|477|2
35.000049|5085791c7fefc7c21148b040e73a112cf04a002e|1.99|2014-12-24 12:36:00|80.700248323638462|2|7203663220|249|35.103207963171322|0|7|330|-80.7007|55|35.06858|EGGS|0.0|3|HT GRADE A    LARGE EGGS|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00072036632203|EGGS FRESH|DAIRY|-80.699686|80.699775519439697|273|1
35.000049|5a1f0ee46b638fd9dceedceb5a35b485a0a0e220|2.19|2015-01-31 14:14:00|80.700248323638462|2|1200000230|249|35.103207819339772|0|7|55|-80.62331|8|35.140781|REGULAR|0.52|23|MTN DEW 2LTR NR|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00012000002335|CARBONATED BEVERAGES|BEVERAGE|-80.699686|80.699914678895297|39|1
35.000049|d51a4c8a3531d838983645055d0cc7dfd145723d|3.99|2015-01-31 14:13:00|80.700248323638462|2|2840000359|249|35.103207819339772|0|7|197|-80.62331|31|35.140781|POPPED POPCORN|0.0|1|SMARTFOOD POPCORN|224f5552bdcbbc3b7a0242ecbb09bcf9949b4b8e|7.128037033786112|35.096297298232479|00028400083591|SNACKS|G1 GROCERY|-80.699686|80.699914678895297|39|1
35.219587|72a6437a0d282066882d7dbb6215a1304fd370f4|16.98|2015-01-02 15:27:00|80.810069425230125|2|3570001820|401|35.246482287430709|0|23|36|-80.844274|10|35.204336|PREMIUM GROUND|4.25|1|COMM COFFEE GROUND CAFE SPEC|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00035700018550|COFFEE|G1 GROCERY|-80.810056|80.810066327628277|61|2
35.219587|c836356a0497778fe02f9ffea98e68660190f5c4|4.99|2015-02-01 13:54:00|80.810069425230125|2|3338390203|401|35.246482287430709|0|23|561|-80.844274|64|35.204336|FR PROD ORGANIC PRODUCE|0.0|4|ORG CARROTS 5LB BAG|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00033383902036|FRESH PRODUCE|PRODUCE|-80.810056|80.810066327628277|61|1
35.219587|170745df57af9bcd3b2697769ffde5c5c821e1f7|4.99|2014-11-30 13:10:00|80.810069425230125|2|3338390203|401|35.246482287341081|0|23|561|-80.826724|64|35.195689|FR PROD ORGANIC PRODUCE|0.0|4|ORG CARROTS 5LB BAG|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00033383902036|FRESH PRODUCE|PRODUCE|-80.810056|80.810066671740415|412|1
35.219587|167d1113f8015d14b52a34e18a961b42b672e3dc|4.99|2015-02-20 16:35:00|80.810069425230125|2|3338390203|401|35.246482287430709|0|23|561|-80.844274|64|35.204336|FR PROD ORGANIC PRODUCE|0.0|4|ORG CARROTS 5LB BAG|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00033383902036|FRESH PRODUCE|PRODUCE|-80.810056|80.810066327628277|61|1
35.219587|64afc889a4f9ff49f330937b327d46eeeb47ad99|4.99|2014-12-28 10:08:00|80.810069425230125|2|3338390203|401|35.246482286601598|0|23|561|-80.80146|64|35.17739|FR PROD ORGANIC PRODUCE|0.0|4|ORG CARROTS 5LB BAG|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00033383902036|FRESH PRODUCE|PRODUCE|-80.810056|80.810069172156702|208|1
35.219587|16b464c752fcfb314328e2951ae3103790a6b785|4.49|2014-11-21 19:16:00|80.810069425230125|2|2840009217|401|35.246482287430709|0|23|1981|-80.844274|480|35.204336|CHIPS|2.24|6|STACY'S MULTIGRAIN PITA CHIP|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00028400092326|DRY GOODS|DELI|-80.810056|80.810066327628277|61|1
35.219587|b103576255272c85347c494d3abb62db8f5e26db|4.49|2014-12-12 13:46:00|80.810069425230125|2|2840009217|401|35.246482287430709|0|23|1981|-80.844274|480|35.204336|CHIPS|2.25|6|STACY'S MULTIGRAIN PITA CHIP|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00028400092326|DRY GOODS|DELI|-80.810056|80.810066327628277|61|1
35.219587|ab016892b030e81338fcff37796c7b8aa5a7837c|14.99|2014-11-14 16:28:00|80.810069425230125|2|3125904695|401|35.246482287341081|0|23|9976|-80.826724|888|35.195689|NFS-U/PREM-PINOT NOIR|0.0|13|JOSH CELLARS PINOT NOIR|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00031259046952|ULTRA PREMIUM ($15-$19.99)|WINE|-80.810056|80.810066671740415|412|1
35.219587|e4771e82c7b7cafe78e0b6c28ef2ec496617a717|0.91|2014-09-28 16:17:00|80.810069425230125|2||401|35.246482287430709|0|23|524|-80.844274|64|35.204336|FRESH PROD FRESH ONIONS|0.0|4|COO YELLOW ONIONS, LRG|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00204665000003|FRESH PRODUCE|PRODUCE|-80.810056|80.810066327628277|61|1
35.219587|aa51d4e36b64b9eaa69df644ee72107671270a89|4.99|2014-09-10 17:13:00|80.810069425230125|2|4082201114|401|35.246482287430709|0|23|1878|-80.844274|435|35.204336|HUMMUS|0.0|6|SPINACH ARTICHOKE HUMMUS|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00040822027540|SALADS|DELI|-80.810056|80.810066327628277|61|1
35.219587|92a9ee5b1663cfc5503e36043ab041133d9fe170|4.99|2014-12-09 16:29:00|80.810069425230125|2|8817722767|401|35.246482287430709|0|23|79|-80.844274|273|35.204336|ASIAN SAUCES/SEASONINGS|0.0|1|SOY VAY HOISIN GARLIC|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00088177227697|ASIAN PREP. FOODS|G1 GROCERY|-80.810056|80.810066327628277|61|1
35.219587|e3a9467e0fb5838b9dee823e66e5e0df0b84d1c3|13.99|2015-01-17 14:17:00|80.810069425230125|2|8378322812|401|35.246482287430709|0|23|458|-80.844274|82|35.204336|CRAFT BEER|0.0|16|SIERRA NEVADA SEASONAL 12PK|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00083783228120|DOMESTIC BEER|BEER|-80.810056|80.810066327628277|61|1
35.219587|619c2e2219d4feb9fb77782cdb6ddac4ffc198c1|1.79|2014-10-15 12:10:00|80.810069425230125|2|2392333002|401|35.246482287430709|0|23|1257|-80.844274|1|35.204336|POUCH BABY FOOD|0.79|1|EB ORG PUMK CRANBRRY APPLE 3RD|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00023923320048|BABY FOOD|G1 GROCERY|-80.810056|80.810066327628277|61|1
35.219587|5ac94f99397961a95596bbc7e229954b2a713f71|7.38|2014-11-14 16:59:00|80.810069425230125|2|3361700703|401|35.246482287430709|0|23|92|-80.844274|13|35.204336|REMAINING CRACKERS|1.38|1|WASA FF MULTIGRAIN CRISPY|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00033617007032|CRACKERS|G1 GROCERY|-80.810056|80.810066327628277|61|2
35.219587|da8202ab9cea5e2a3d9aa2ad67e2117e1e2e59ea|6.79|2014-10-08 17:28:00|80.810069425230125|2|38151901931|401|35.246482287430709|0|23|3503|-80.844274|1045|35.204336|CONDITIONER-PREMIUM|0.8|17|HERBAL ESS H/HYDRA MOIS COND|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00381519019289|HAIR & SCALP CARE|HBC|-80.810056|80.810066327628277|61|1
35.219587|4c9e5b574d8d16973078058736c40ef12009ac6c|3.36|2014-12-13 10:18:00|80.810069425230125|2||401|35.246482286601598|0|23|502|-80.80146|64|35.17739|FRESH BANANAS|0.0|4|BANANAS, YELLOW|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00204011000008|FRESH PRODUCE|PRODUCE|-80.810056|80.810069172156702|208|2
35.219587|237cdf598638d8fa7d4e20625d04630f6d3bb6b4|1.59|2015-01-26 18:48:00|80.810069425230125|2||401|35.246482287430709|0|23|502|-80.844274|64|35.204336|FRESH BANANAS|0.0|4|BANANAS, YELLOW|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00204011000008|FRESH PRODUCE|PRODUCE|-80.810056|80.810066327628277|61|1
35.219587|ad6774ec5753c80090e1223a1bfb5c25c8ccfc45|1.99|2014-10-10 16:47:00|80.810069425230125|2|7225100154|401|35.246482287430709|0|23|240|-80.844274|38|35.204336|COUS/ALT GRAINS|0.0|1|NEAR EAST COUSCOUS CHKN HERB|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00072251001532|RICE GRAINS AND BEANS|G1 GROCERY|-80.810056|80.810066327628277|61|1
35.219587|015cef5264ecc7bbbd105ff247835845bc7dafd2|1.39|2014-10-22 12:48:00|80.810069425230125|2|2200000488|401|35.246482283307614|0|23|48|-80.85013|7|35.175855|REGISTER GUM|0.2|1|(FE)ORBIT PEPPERMINT GUM 14PC|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00022000004864|CANDY|G1 GROCERY|-80.810056|80.810076954188915|218|1
35.219587|e0f8678a7ad9e88dda66b4bd416d8d94d1eb6db9|3.99|2014-10-31 15:06:00|80.810069425230125|2|2800074797|401|35.246482287430709|0|23|727|-80.844274|7|35.204336|SEASONAL CANDY-SINGLE FAC|0.49|1|I/O(H15)BABY RUTH FUN SIZE|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00028000747978|CANDY|G1 GROCERY|-80.810056|80.810066327628277|61|1
35.219587|76fcae868a0a7145929773dd248b9eb56d1847e8|4.49|2014-10-30 18:31:00|80.810069425230125|2|2840009217|401|35.246482287430709|0|23|1981|-80.844274|480|35.204336|CHIPS|0.0|6|STACY'S PITA CHIPS NAKED|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00028400092173|DRY GOODS|DELI|-80.810056|80.810066327628277|61|1
35.219587|3d20516d2e86f9f17c03ae5a17ae3a8c55b6da49|5.98|2014-12-08 16:53:00|80.810069425230125|2||401|35.246482287430709|0|23|561|-80.844274|64|35.204336|FR PROD ORGANIC PRODUCE|0.99|4|COO ORG KALE|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00294627000004|FRESH PRODUCE|PRODUCE|-80.810056|80.810066327628277|61|2
35.219587|2a0a95cfbb4dfdfe62dc2f2ffe1337df737bae7c|2.59|2014-11-30 12:21:00|80.810069425230125|2|85832876218|401|35.246482287430709|0|23|1201|-80.844274|33|35.204336|RTS CANNED|0.0|1|WOLF PUCK ORGANIC CORN CHOWDER|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00858328761901|SOUP|G1 GROCERY|-80.810056|80.810066327628277|61|1
35.219587|237f0c0f06082b170341a199420b22f1d239b016|6.79|2015-01-19 18:14:00|1.4094857484078087|2|38151901931|401|0.6146977543425921|0|26|3536|-80.810056|1045|35.219587|SHAMPOO-PREMIUM|0.8|17|HERBAL ESS H/HYDRATE MOIS SHAM|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|0.61471665291522548|00381519019258|HAIR & SCALP CARE|HBC|-80.810056|1.4104015459209989|401|1
35.219587|ebf1e96622586ef8169c01980f38fb3981b426e5|3.38|2014-12-30 14:59:00|80.810069425230125|2|73801577715|401|35.246482287430709|0|23|545|-80.844274|64|35.204336|FRESH SPROUTS|0.19|4|BLACK-EYED PEAS, PKG|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00738015777159|FRESH PRODUCE|PRODUCE|-80.810056|80.810066327628277|61|2
35.219587|8f883045642da935569eca8f5db29afd7da86304|2.67|2014-11-02 14:57:00|80.810069425230125|2|7203698754|401|35.246482287430709|0|23|1265|-80.844274|57|35.204336|ALMOND MILK|0.17|3|HT ALMOND DRINK UNSWT ORIGINAL|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00072036707352|MILK|DAIRY|-80.810056|80.810066327628277|61|1
35.219587|d59f0d208fbe4a55d2b2b3c91cb860372c22edcc|5.69|2014-10-04 20:28:00|80.810069425230125|2|20541900000|401|35.246482280901937|0|23|1832|-80.825175|415|35.152722|BH SLICING CHEESE|0.57|6|BOARS HEAD LACEY SWISS CHEESE|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00205419000003|SLICING CHEESE|DELI|-80.810056|80.8100811601185|160|1
35.219587|7630f8852114137e1232e4d6e2341f41e60c068d|1.0|2014-10-13 17:51:00|80.810069425230125|2||401|35.246482283307614|0|23|509|-80.85013|64|35.175855|FRESH CITRUS-REMAINING|0.0|4|COO LIMES, LRG|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00204048000002|FRESH PRODUCE|PRODUCE|-80.810056|80.810076954188915|218|2
35.219587|ce2ef4be42a2b7b41b5a624545a16ba577ccd052|6.99|2014-10-27 15:40:00|80.810069425230125|2|7203670333|401|35.246482287430709|0|23|443|-80.844274|76|35.204336|NFS-GARBAGE BAGS|1.22|1|YH TALL KTCHN ODOR CNTL|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00072036703460|WRAPPING MATERIALS & BAGS|G1 GROCERY|-80.810056|80.810066327628277|61|1
35.219587|3df49fdcd66452457a155f181205548fb39d0425|3.29|2014-10-04 11:54:00|80.810069425230125|2|2840004768|401|35.246482287430709|0|23|202|-80.844274|31|35.204336|PRETZELS|0.29|1|ROLD GOLD PRETZEL TINY TWIST|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00028400047685|SNACKS|G1 GROCERY|-80.810056|80.810066327628277|61|1
35.219587|6f7bef0aada608c75a2662f8f7231d2bab54acbb|3.69|2014-12-02 16:41:00|80.810069425230125|2|2100062503|401|35.246482283307614|0|23|318|-80.85013|52|35.175855|SHREDDED/GRATED CHEESE|0.69|3|KRAFT 2% MEXICAN FOUR CHEESE|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00021000024612|CHEESE|DAIRY|-80.810056|80.810076954188915|218|1
35.219587|223d7edd973578ae44321ce5045f97c7057a1138|3.49|2015-01-23 08:09:00|80.810069425230125|2|7203697601|401|35.246482261662102|0|23|4612|-80.771677|1215|35.066546|VITAMIN-MINERALS|0.0|17|HT NAT ZINC 50MG TABS 97601|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00072036976017|VITAMINS & SUPPLEMENTS|HBC|-80.810056|80.810102735571007|45|1
35.219587|a64511b794e98a89cac0666b925ec653067111bf|3.49|2014-11-13 13:30:00|80.810069425230125|2|7203697601|401|35.246482287430709|0|23|4612|-80.844274|1215|35.204336|VITAMIN-MINERALS|0.0|17|HT NAT ZINC 50MG TABS 97601|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00072036976017|VITAMINS & SUPPLEMENTS|HBC|-80.810056|80.810066327628277|61|1
35.219587|993c321428eb02a0148b2637b68ff9be0707d63d|4.99|2015-02-06 16:43:00|80.810069425230125|2|4082201114|401|35.246482287430709|0|23|1878|-80.844274|435|35.204336|HUMMUS|1.0|6|HUMMUS W/ ROASTED PINE NUTS|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00040822011747|SALADS|DELI|-80.810056|80.810066327628277|61|1
35.219587|9727769da55771e2a8aa2b7bf3f6bea97b17c025|4.99|2014-11-23 18:28:00|80.810069425230125|2|7203688187|401|35.246482287430709|0|23|561|-80.844274|64|35.204336|FR PROD ORGANIC PRODUCE|0.0|4|ORG HT BABY SPINACH 11 OZ|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00072036881878|FRESH PRODUCE|PRODUCE|-80.810056|80.810066327628277|61|1
35.219587|b39a084c063136b6584a7e05e90f6af6b0ea35a2|4.69|2015-01-06 18:46:00|80.810069425230125|2|7203676448|401|35.246482287430709|0|23|239|-80.844274|38|35.204336|RICE-PACKAGED & BULK|0.0|1|HTO RICE BROWN BASMATI|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00072036764508|RICE GRAINS AND BEANS|G1 GROCERY|-80.810056|80.810066327628277|61|1
35.219587|d2051b12093a200c9bf73675245b698c6e49dd44|4.99|2014-10-19 18:17:00|80.810069425230125|2|7203688187|401|35.246482287430709|0|23|561|-80.844274|64|35.204336|FR PROD ORGANIC PRODUCE|0.0|4|ORG HT BABY SPINACH 11 OZ|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00072036881878|FRESH PRODUCE|PRODUCE|-80.810056|80.810066327628277|61|1
35.219587|be30d0a189dcf7ede5f60ff1e565009da6f3fefa|4.99|2015-02-25 15:43:00|80.810069425230125|2|7203688187|401|35.246482287430709|0|23|561|-80.844274|64|35.204336|FR PROD ORGANIC PRODUCE|0.0|4|ORG HT BABY SPINACH 11 OZ|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00072036881878|FRESH PRODUCE|PRODUCE|-80.810056|80.810066327628277|61|1
35.219587|898ba14b6eb5f57da69347d664a74717ff3ff66f|0.99|2014-11-30 15:16:00|80.810069425230125|2||401|35.246482287430709|0|23|540|-80.844274|64|35.204336|FRESH CELERY|0.0|4|COO CELERY (RPC) 24'S|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00204070000001|FRESH PRODUCE|PRODUCE|-80.810056|80.810066327628277|61|1
35.219587|5996ee6a1b665d2fdf7b49e41658378cbb1e4fc4|3.89|2014-11-08 18:07:00|80.810069425230125|2|7684010015|401|35.246482287430709|0|23|275|-80.844274|45|35.204336|SUPER PREMIUM ICE CREAM|0.0|5|BEN & JERRY FRO YO FDGE BRW|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00076840100569|ICE CREAM|FROZEN|-80.810056|80.810066327628277|61|1
35.219587|9e88642f75369d40f3d83fe2d3e3a00f8da48b6d|4.99|2014-11-20 15:23:00|80.810069425230125|2|7336070341|401|35.246482287341081|0|23|30|-80.826724|4|35.195689|CARBONATED WATER|1.49|1|LACROIX WTR PLAIN 12PK|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00073360703416|BOTTLED WATER|G1 GROCERY|-80.810056|80.810066671740415|412|1
35.219587|c9811a8fd8a60009fc86ac24ea7c1fd887b9fcf5|5.99|2015-01-12 08:22:00|80.810069425230125|2|7214045231|401|35.246482261662102|0|23|3202|-80.771677|1015|35.066546|HAND & BODY THERAPEUTIC|0.0|17|AQUAPHOR HEALING OINTMENT|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00072140452315|HAND & BODY LOTION/SUN CARE|HBC|-80.810056|80.810102735571007|45|1
35.219587|0665d1070b2682d846efcf3f07da563b05d18989|3.25|2015-01-13 16:25:00|80.810069425230125|2|4157005617|401|35.246482287430709|0|23|1265|-80.844274|57|35.204336|ALMOND MILK|0.0|3|ALMOND BREEZE UNSWEET ORIGINAL|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00041570056707|MILK|DAIRY|-80.810056|80.810066327628277|61|1
35.219587|5f847afc34f31b6af651fa2791bd6729debef57d|0.79|2014-09-21 14:02:00|80.810069425230125|2|7203688001|401|35.246482280557707|0|23|527|-80.849471|64|35.161696|FRESH CARROTS|0.0|4|HT WHOLE CARROTS 1LB BAG|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00072036880017|FRESH PRODUCE|PRODUCE|-80.810056|80.81008170574728|35|1
35.219587|46141bea99ccbd5b0d07279b0d3fa01ec66aefda|3.99|2015-02-11 16:49:00|80.810069425230125|2|7203676145|401|35.246482287430709|0|23|1211|-80.844274|272|35.204336|HISP SALSA/DIPS|0.99|1|HT TRADER SALSA BEAN&CORN|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00072036761514|HISPANIC PREP. FOODS|G1 GROCERY|-80.810056|80.810066327628277|61|1
35.219587|27afbac46b3a0e76e6901f6e3b415064ef938d5b|13.98|2014-09-20 10:42:00|80.810069425230125|2|7203698736|401|35.246482240020782|0|23|4454|-80.848528|1210|35.053394|DIGESTIVE AID-SWALLOWABLE|2.19|17|HT DAIRY RELIEF-DIG CAP|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00072036987365|STOMACH REMEDIES|HBC|-80.810056|80.810118681811019|11|2
35.219587|bb4132dad222f83a28d348a1ef6627063aa3ad76|2.26|2014-09-23 17:06:00|80.810069425230125|2||401|35.246482283307614|0|23|502|-80.85013|64|35.175855|FRESH BANANAS|0.0|4|BANANAS, YELLOW|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00204011000008|FRESH PRODUCE|PRODUCE|-80.810056|80.810076954188915|218|1
35.219587|3edf8955bf165f9cd66f461900e13fb5eb18ed2a|3.15|2014-09-15 15:14:00|80.810069425230125|2|7203603083|401|35.246482287430709|0|23|30|-80.844274|4|35.204336|CARBONATED WATER|0.0|1|HT ORIGINAL SELTZER 12 PK|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00072036030832|BOTTLED WATER|G1 GROCERY|-80.810056|80.810066327628277|61|1
35.219587|893ebb9725203489186fe54127baebc1b1e832d1|12.99|2015-02-09 16:31:00|80.810069425230125|2|8378316000|401|35.246482287430709|0|23|458|-80.844274|82|35.204336|CRAFT BEER|0.0|16|SIERRA NEVADA SEASONAL|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00083783160000|DOMESTIC BEER|BEER|-80.810056|80.810066327628277|61|1
35.219587|594431bdc41d22e88aae582a4d1e47ed6fb1fa6b|12.99|2015-02-04 17:07:00|80.810069425230125|2|8378316000|401|35.246482287430709|0|23|458|-80.844274|82|35.204336|CRAFT BEER|0.0|16|SIERRA NEVADA SEASONAL|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00083783160000|DOMESTIC BEER|BEER|-80.810056|80.810066327628277|61|1
35.219587|df1bd3c9f9d84b07397a5e7a30f2c0ba6ace8c02|13.99|2015-02-16 14:41:00|80.810069425230125|2|8378316000|401|35.246482287430709|0|23|458|-80.844274|82|35.204336|CRAFT BEER|0.0|16|SIERRA NEVADA SEASONAL|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00083783160000|DOMESTIC BEER|BEER|-80.810056|80.810066327628277|61|1
35.219587|50d2e62946dceee96d9c2e029b4dee23782a9268|13.99|2015-03-04 16:24:00|80.810069425230125|2|75452700201|401|35.246482287430709|0|23|458|-80.844274|82|35.204336|CRAFT BEER|0.0|16|NEW BELGIUM FOLLY VARIETY 12PK|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00754527002015|DOMESTIC BEER|BEER|-80.810056|80.810066327628277|61|1
35.219587|9e43a5f96a2b04cb898671caedbaee051234ee8e|7.99|2014-12-05 18:32:00|80.810069425230125|2|75452700122|401|35.246482287430709|0|23|458|-80.844274|82|35.204336|CRAFT BEER|0.0|16|NEW BELGUIM 1554 BLACK ALE 6PK|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00754527001223|DOMESTIC BEER|BEER|-80.810056|80.810066327628277|61|1
35.219587|08dc4a3fe68a88e77010886ee449eca5b4764c78|3.99|2015-01-09 15:23:00|80.810069425230125|2|7203602701|401|35.246482261662102|0|23|1878|-80.771677|435|35.066546|HUMMUS|1.99|6|FFM ARTISAN CARM. ONION HUMMUS|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00072036027047|SALADS|DELI|-80.810056|80.810102735571007|45|1
35.219587|93524a4fabcaeddb0d256499aec9748d92ec7be7|3.99|2014-11-12 20:49:00|80.810069425230125|2|7203602701|401|35.246482287430709|0|23|1878|-80.844274|435|35.204336|HUMMUS|1.99|6|FFM ARTISAN CARM. ONION HUMMUS|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00072036027047|SALADS|DELI|-80.810056|80.810066327628277|61|1
35.219587|1474663952bae769dbb2569531732ecf50864eb5|2.91|2014-12-24 16:05:00|80.810069425230125|2|7203698757|401|35.246482287430709|0|23|31|-80.844274|4|35.204336|NON CARBONATED WATER|0.0|1|HT PURIFIED WATER|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00072036987570|BOTTLED WATER|G1 GROCERY|-80.810056|80.810066327628277|61|3
35.219587|1dbc87e748158e2d514add44f0a98d5530383d20|4.9|2015-03-06 16:17:00|80.810069425230125|2||401|35.246482287430709|0|23|500|-80.844274|64|35.204336|FRESH APPLES|2.46|4|FUJI APPLES|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00204131000001|FRESH PRODUCE|PRODUCE|-80.810056|80.810066327628277|61|1
35.219587|4296c1942b48a4b69f61e0d4186db207af9014ab|4.49|2015-01-01 15:28:00|80.810069425230125|2|4812127707|401|35.246482287430709|0|23|1036|-80.844274|164|35.204336|BREAKFAST BAGELS|2.25|7|THOMAS  RAISIN BAGELS 6CT PP|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00048121292089|BREAKFAST|COMMERCIAL BAKERY|-80.810056|80.810066327628277|61|1
35.219587|4a21a815f3eeeb5da353061a7151f13895d3d2d1|4.59|2014-11-07 16:07:00|80.810069425230125|2|78142100128|401|35.246482287341081|0|23|1601|-80.826724|371|35.195689|BRANDED BREAD|1.15|14|LA BREA SOURDOUGH LOAF|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00781421001288|BREAD|BAKERY|-80.810056|80.810066671740415|412|1
35.219587|c20f8af9071a0defba5b5fa3d1898ce9315fb1a9|7.99|2014-12-24 13:37:00|80.810069425230125|2|7203676196|401|35.246482283307614|0|23|36|-80.85013|10|35.175855|PREMIUM GROUND|2.42|1|HT TRADERS TOASTED ALMOND|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00072036978592|COFFEE|G1 GROCERY|-80.810056|80.810076954188915|218|1
35.219587|19ed3db1c6fb5db5e933826e6df1d81e0641a38c|2.93|2014-12-19 14:25:00|80.810069425230125|2|20165900000|401|35.246482287430709|0|23|297|-80.844274|49|35.204336|GROUND BEEF|0.0|2|GROUND BEEF 93% LEAN|233ca925d5f30b2ccd610426cefd38acd1d33223|1.8583995030798608|35.240679762029046|00201659000001|BEEF|MEAT|-80.810056|80.810066327628277|61|1
34.937113|4f36174fce29676e74b348560afb0b7ee8fc38e3|5.34|2014-09-23 19:22:00|80.849735164501183|4|7203698754|372|35.606142586351922|0|11|1265|-80.764523|57|35.341927|ALMOND MILK|0.0|3|HT ALMOND DRINK UNSWT ORIGINAL|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00072036707352|MILK|DAIRY|-80.837892|80.841632113361626|220|2
34.937113|6a71f4c61c923ff3511a7e7f8fdf30726fb40eb6|2.67|2014-11-22 21:56:00|80.849735164501183|4|7203698754|372|35.606142586351922|0|11|1265|-80.764523|57|35.341927|ALMOND MILK|0.17|3|HT ALMOND DRINK UNSWT ORIGINAL|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00072036707352|MILK|DAIRY|-80.837892|80.841632113361626|220|1
34.937113|f97a5c4626ff604aa57515be19c03fd6232c2ad8|3.19|2014-10-25 20:19:00|80.849735164501183|4|7231000041|372|35.606143602027274|0|11|230|-80.737839|37|35.297134|HERBAL TEA|0.0|1|BIGELOW TEA HERB PEPPERMINT|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00072310000391|TEA|G1 GROCERY|-80.837892|80.841348801086681|258|1
34.937113|efae26a9e752ad3cff76a12af99e20aff0b19215|5.34|2015-03-04 14:26:00|80.849735164501183|4|7203698754|372|35.606148297678345|0|11|1265|-80.824767|57|35.116751|ALMOND MILK|0.0|3|HT ALMOND DRINK UNSWT ORIGINAL|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00072036707352|MILK|DAIRY|-80.837892|80.839480359505345|294|2
34.937113|8d849abae7f3f144b3859c22ed29227c39cb5812|2.67|2014-09-18 19:40:00|80.849735164501183|4|7203698754|372|35.606142586351922|0|11|1265|-80.764523|57|35.341927|ALMOND MILK|0.0|3|HT ALMOND DRINK UNSWT ORIGINAL|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00072036707352|MILK|DAIRY|-80.837892|80.841632113361626|220|1
34.937113|3e1ef9fa126d645b0e606368c6da8253ae3e74e7|2.49|2014-10-07 15:42:00|80.849735164501183|4|71157510200|372|35.606142586351922|0|11|1244|-80.764523|21|35.341927|OTHER NUTS|0.0|1|SEAPOINT FARM WASABI EDAMAME|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00711575102104|NUTS|G1 GROCERY|-80.837892|80.841632113361626|220|1
34.937113|f5973349286df87f29ca83943324d32b04391573|2.67|2014-09-16 17:30:00|80.849735164501183|4|7203698754|372|35.606143602027274|0|11|1265|-80.737839|57|35.297134|ALMOND MILK|0.0|3|HT ALMOND DRINK UNSWT VANILLA|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00072036987563|MILK|DAIRY|-80.837892|80.841348801086681|258|1
34.937113|182b1cbf6bea34172c909c2ab081c464e9c92c47|4.39|2015-02-28 12:53:00|80.849735164501183|4|4400002796|372|35.606142586351922|0|11|90|-80.764523|13|35.341927|SNACK CRACKERS|2.2|1|TRISCUITS THIN CRISPS WASABSOY|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00044000037826|CRACKERS|G1 GROCERY|-80.837892|80.841632113361626|220|1
34.937113|4bff09ecd0e5b307ea3409b4174694b3fb874a8f|4.39|2014-12-23 16:46:00|80.849735164501183|4|4400002796|372|35.606143602027274|0|11|90|-80.737839|13|35.297134|SNACK CRACKERS|2.2|1|TRISCUITS THIN CRISPS WASABSOY|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00044000037826|CRACKERS|G1 GROCERY|-80.837892|80.841348801086681|258|1
34.937113|2e85401811940a91fa9e9c50758305b3004777b8|3.49|2014-12-03 20:20:00|80.849735164501183|4|4180050126|372|35.606143602027274|0|11|123|-80.737839|19|35.297134|JELLY/JAMS|0.0|1|WELCH'S NATURAL SPREADS GRAPE|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00041800501267|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.837892|80.841348801086681|258|1
34.937113|430c038948795d2213f2a562b4dc98f9ebd4c1be|3.49|2014-10-21 20:49:00|80.849735164501183|4|4180050126|372|35.606143602027274|0|11|123|-80.737839|19|35.297134|JELLY/JAMS|0.0|1|WELCH'S NATURAL SPREADS GRAPE|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00041800501267|JAMS/JELLIES/SPREADS|G1 GROCERY|-80.837892|80.841348801086681|258|1
34.937113|47e6c9995e2612955ea86f2d2828d253c9eceed4|1.89|2015-02-03 17:32:00|80.849735164501183|4|7920022288|372|35.606143602027274|0|11|50|-80.737839|7|35.297134|PEG CANDY|0.39|1|SWEETART MINI CHEWY PEG BAG|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00079200222888|CANDY|G1 GROCERY|-80.837892|80.841348801086681|258|1
34.937113|319b493baa6427fce26a84342cbdd189d4049802|0.99|2014-11-25 12:20:00|80.849735164501183|4|7203695306|372|35.606143602027274|0|11|1895|-80.737839|450|35.297134|TEA|0.0|6|FFM DIET TEA W/SPLENDA|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00072036018892|BEVERAGES|DELI|-80.837892|80.841348801086681|258|1
34.937113|efd26d0545e9c1515efd64b1f83f014a8c223d17|0.99|2015-01-22 17:12:00|80.849735164501183|4|7203695306|372|35.606143602027274|0|11|1895|-80.737839|450|35.297134|TEA|0.0|6|FFM DIET TEA W/SPLENDA|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00072036018892|BEVERAGES|DELI|-80.837892|80.841348801086681|258|1
34.937113|af113ce9c1c40e0bfe69963a49b8c93ade01d396|7.98|2014-11-18 12:14:00|80.849735164501183|4|7203602701|372|35.606143602027274|0|11|1878|-80.737839|435|35.297134|HUMMUS|1.99|6|FFM ARTISAN PINE NUT HUMMUS|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00072036027054|SALADS|DELI|-80.837892|80.841348801086681|258|2
34.937113|a31c3c73a4aac77cd9f38a4d045d14e6b353feab|3.99|2014-12-05 12:03:00|80.849735164501183|4|7203602701|372|35.606143602027274|0|11|1878|-80.737839|435|35.297134|HUMMUS|0.5|6|FFM ARTISAN PINE NUT HUMMUS|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00072036027054|SALADS|DELI|-80.837892|80.841348801086681|258|1
34.937113|bd079681f1716c09f84deda27d127b7d12e2e63f|3.99|2014-10-23 19:59:00|80.849735164501183|4|7203602701|372|35.606143602027274|0|11|1878|-80.737839|435|35.297134|HUMMUS|1.99|6|FFM ARTISAN PINE NUT HUMMUS|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00072036027054|SALADS|DELI|-80.837892|80.841348801086681|258|1
34.937113|f9e5c75b012e4e78e90b7717623c460b1b28f4f2|3.99|2014-11-10 17:04:00|80.849735164501183|4|7203602701|372|35.606143602027274|0|11|1878|-80.737839|435|35.297134|HUMMUS|0.5|6|FFM ARTISAN PINE NUT HUMMUS|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00072036027054|SALADS|DELI|-80.837892|80.841348801086681|258|1
34.937113|eb067184f1c816d2d50be3e2ddde90d20b7c9a5a|3.99|2014-12-01 14:24:00|80.849735164501183|4|7203602701|372|35.606143602027274|0|11|1878|-80.737839|435|35.297134|HUMMUS|0.5|6|FFM ARTISAN PINE NUT HUMMUS|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00072036027054|SALADS|DELI|-80.837892|80.841348801086681|258|1
34.937113|16e7ef2781e3e670c6c7f68c42bbe06f74a05f1f|2.39|2014-09-23 16:25:00|80.849735164501183|4|5440000080|372|35.606143602027274|0|11|82|-80.737839|11|35.297134|VINEGAR|0.72|1|REGINA RED WINE VINEGAR|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00054400000801|CONDIMENTS|G1 GROCERY|-80.837892|80.841348801086681|258|1
34.937113|8f325442a465481eb9af67f7c2f87498f51f41a6|5.39|2015-03-04 14:17:00|80.849735164501183|4|4900006381|372|35.606148297678345|0|11|31|-80.824767|4|35.116751|NON CARBONATED WATER|0.4|1|DASANI SPARKLING BLK CHERRY|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00049000065527|BOTTLED WATER|G1 GROCERY|-80.837892|80.839480359505345|294|1
34.937113|dabf00dd8d1fa6c82c1772b411e91e311d5f5ff6|3.29|2014-10-27 19:31:00|80.849735164501183|4|2840018382|372|35.606143602027274|0|11|201|-80.737839|31|35.297134|POTATO CHIPS|0.79|1|BAKED CHEETOS REGULAR|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00028400183901|SNACKS|G1 GROCERY|-80.837892|80.841348801086681|258|1
34.937113|1252157cb91662417d11f01b72a6798c760574b9|11.59|2014-10-01 20:17:00|80.849735164501183|4|3680024419|372|35.606143602027274|0|11|4186|-80.737839|1200|35.297134|ALLERGY REMEDY-ADULT|0.0|17|TC A/D ALLRGY-CETIRIZINE 10MG|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00036800244191|COUGH/COLD/SINUS|HBC|-80.837892|80.841348801086681|258|1
34.937113|5a7abfe6547c2b028d45ad2218e75ec8a78dcc2b|3.49|2014-11-20 12:43:00|80.849735164501183|4|7797509126|372|35.606143602027274|0|11|202|-80.737839|31|35.297134|PRETZELS|0.49|1|SPECIAL DRK CHOC PRETZEL DIPS|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00077975082478|SNACKS|G1 GROCERY|-80.837892|80.841348801086681|258|1
34.937113|c6b46c25a13ace5a49503305001e827d9297badb|3.49|2014-12-02 08:48:00|80.849735164501183|4|7797509126|372|35.606143602027274|0|11|202|-80.737839|31|35.297134|PRETZELS|0.49|1|SPECIAL DRK CHOC PRETZEL DIPS|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00077975082478|SNACKS|G1 GROCERY|-80.837892|80.841348801086681|258|1
34.937113|12e94fec87d4d6e845566e6163bd8a74c4df3756|0.95|2014-11-11 13:23:00|80.849735164501183|4||372|35.606143602027274|0|11|502|-80.737839|64|35.297134|FRESH BANANAS|0.0|4|BANANAS, YELLOW|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00204011000008|FRESH PRODUCE|PRODUCE|-80.837892|80.841348801086681|258|1
34.937113|677dcc95c5e8b3316d8db5143ab5704555f46a56|1.4|2014-10-07 13:03:00|80.849735164501183|4||372|35.606143602027274|0|11|502|-80.737839|64|35.297134|FRESH BANANAS|0.0|4|BANANAS, YELLOW|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00204011000008|FRESH PRODUCE|PRODUCE|-80.837892|80.841348801086681|258|1
34.937113|ee5de7a7aea0afae468a18c14204f8eba17f8645|4.99|2014-12-11 12:02:00|80.849735164501183|4|4082201114|372|35.606143602027274|0|11|1878|-80.737839|435|35.297134|HUMMUS|4.99|6|ROASTED GARLIC HUMMUS|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00040822011242|SALADS|DELI|-80.837892|80.841348801086681|258|1
34.937113|77916a7804710d4bcedbf8d214c4e3d383fb0f70|2.0|2014-11-26 16:40:00|80.849735164501183|4|4000000435|372|35.606143602027274|0|11|47|-80.737839|7|35.297134|REGISTER BARS|0.2|1|(FE)SNICKERS CANDY BAR|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00040000424314|CANDY|G1 GROCERY|-80.837892|80.841348801086681|258|2
34.937113|767ca642c8f6317a159107d19d2d6c27acbbab3e|3.55|2014-10-15 16:14:00|80.849735164501183|4|4157005617|372|35.606142586351922|0|11|1265|-80.764523|57|35.341927|ALMOND MILK|1.05|3|ALMOND BREEZE UNSWEET ORIGINAL|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00041570056707|MILK|DAIRY|-80.837892|80.841632113361626|220|1
34.937113|15a7a796934ee50ab4cdd13994420735d3dff552|2.27|2015-02-28 13:16:00|80.849735164501183|4|2200015586|372|35.606142586351922|0|11|45|-80.764523|7|35.341927|PEG GUM|0.0|1|ORBIT PEPPERMINT|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00022000155863|CANDY|G1 GROCERY|-80.837892|80.841632113361626|220|1
34.937113|6ee2192ab22e539e791cf13e727c3d15d848baf6|1.99|2015-02-10 20:56:00|80.849735164501183|4|60322422423|372|35.606138359231167|0|11|533|-80.860108|64|35.500972|FRESH PEPPERS|0.0|4|MINI SWEET PEPPERS 1LB|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00603224224230|FRESH PRODUCE|PRODUCE|-80.837892|80.842632715528794|268|1
34.937113|ba5126d45667d2aa325f59e536a050045971072f|4.99|2014-11-26 16:37:00|80.849735164501183|4|4082201114|372|35.606143602027274|0|11|1878|-80.737839|435|35.297134|HUMMUS|1.99|6|HUMMUS W/ ROASTED PINE NUTS|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00040822011747|SALADS|DELI|-80.837892|80.841348801086681|258|1
34.937113|a3d924b1d287705eff6c5d04f1dad6195f3dd780|2.25|2014-10-27 19:25:00|80.849735164501183|4||372|35.606143602027274|0|11|502|-80.737839|64|35.297134|FRESH BANANAS|0.0|4|BANANAS, YELLOW|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00204011000008|FRESH PRODUCE|PRODUCE|-80.837892|80.841348801086681|258|1
34.937113|a6a1fdb365bf488770c580736efe7412b37848a1|5.99|2014-10-16 21:09:00|80.849735164501183|4|8043234107|372|35.606143602027274|0|11|9935|-80.737839|885|35.297134|NFS POP CAB SAUV|0.0|13|JACOBS CREEK CABERNET SAUV|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00080432341070|POPULAR (4-$7.99)|WINE|-80.837892|80.841348801086681|258|1
34.937113|b332a6d66c626db6efd9a48a0237a16a1c9c2622|1.19|2014-12-12 09:40:00|80.849735164501183|4|7433686394|372|35.606143602027274|0|11|342|-80.737839|57|35.297134|FRESH MILK|0.2|3|HUNTER 2% MILK 14 OZ|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00074336863950|MILK|DAIRY|-80.837892|80.841348801086681|258|1
34.937113|7ffc91099e87bede3727f125eb78ffff3fe3d7d7|1.19|2014-12-10 12:55:00|80.849735164501183|4|7433686394|372|35.606143602027274|0|11|342|-80.737839|57|35.297134|FRESH MILK|0.2|3|HUNTER 2% MILK 14 OZ|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00074336863950|MILK|DAIRY|-80.837892|80.841348801086681|258|1
34.937113|e279175d829dc46711b8a425f5d9f5f32be7299f|3.29|2014-11-24 12:36:00|80.849735164501183|4|2840004768|372|35.606143602027274|0|11|202|-80.737839|31|35.297134|PRETZELS|0.29|1|ROLD GOLD PRETZEL STICKS|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00028400047708|SNACKS|G1 GROCERY|-80.837892|80.841348801086681|258|1
34.937113|483e7475a1dfbdc3f7a49227cbb15b5cd9df2f6a|3.29|2015-01-29 12:57:00|80.849735164501183|4|2840018382|372|35.606143602027274|0|11|201|-80.737839|31|35.297134|POTATO CHIPS|0.29|1|BAKED LAYS BBQ|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00028400183833|SNACKS|G1 GROCERY|-80.837892|80.841348801086681|258|1
34.937113|821087dcd2829ee3b5da5fc8f3d134988189e8e4|7.98|2014-11-11 20:08:00|80.849735164501183|4|74447391224|372|35.606143602027274|0|11|1265|-80.737839|57|35.297134|ALMOND MILK|1.49|3|SO DELICIOUS UNSWT ALMOND MILK|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00744473912254|MILK|DAIRY|-80.837892|80.841348801086681|258|2
34.937113|16b8c3cdf48c5a6382e878708450bdf080cbc2e0|4.29|2014-10-28 14:37:00|80.849735164501183|4|84357100478|372|35.606143602027274|0|11|197|-80.737839|31|35.297134|POPPED POPCORN|1.29|1|POP IND AGED WHITE CHED POPCRN|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00843571004745|SNACKS|G1 GROCERY|-80.837892|80.841348801086681|258|1
34.937113|dc710f1db870e3cc763fd7921e93d5afcdd7a50f|3.99|2014-12-16 20:06:00|80.849735164501183|4|3338300084|372|35.606148915358652|0|11|500|-80.816172|64|35.059823|FRESH APPLES|0.0|4|GOLD DEL APPLE 3LB BAG|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00072036880277|FRESH PRODUCE|PRODUCE|-80.837892|80.839024642357572|66|1
34.937113|8d952c2fe25dce5a2bd42557703c2a33b16e376f|6.49|2014-10-27 14:59:00|80.849735164501183|4|2301200051|372|35.606143602027274|0|11|1475|-80.737839|485|35.297134|SUSHI CLASSIC|0.0|6|VEGETABLE COMBO (BROWN RICE)|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00023012000516|SUSHI|DELI|-80.837892|80.841348801086681|258|1
34.937113|f9eb0f5e2586e6fdf4667c9e5a364283a0897b70|7.99|2014-12-02 13:19:00|80.849735164501183|4|2301200207|372|35.606143602027274|0|11|1475|-80.737839|485|35.297134|SUSHI CLASSIC|0.0|6|CRUNCHY SHRIMP ROLL|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00023012002077|SUSHI|DELI|-80.837892|80.841348801086681|258|1
34.937113|9484a502fe36945d22b5b55d9aeec78b5894898a|7.13|2015-02-18 18:27:00|80.849735164501183|4|27061900000|372|35.606143602027274|0|11|973|-80.737839|201|35.297134|FRESH PERDUE CHICKEN|0.0|2|PERDUE THIN CUT BNLS BREAST|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00270619000009|POULTRY|MEAT|-80.837892|80.841348801086681|258|1
34.937113|c93879ae3176006bf6acb5fe4eff2efb4a178f3d|3.89|2014-10-29 20:02:00|80.849735164501183|4|4400003219|372|35.606143602027274|0|11|1249|-80.737839|12|35.297134|CHOCOLATE CHIP COOKIES|0.9|1|CHIPS AHOY ORIG CHOCOLATE CHIP|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00044000032197|COOKIES|G1 GROCERY|-80.837892|80.841348801086681|258|1
34.937113|14863ad12ba1f7b9350caf48a5fc34c31bc74817|2.38|2014-12-04 12:36:00|80.849735164501183|4|7433686394|372|35.606143602027274|0|11|342|-80.737839|57|35.297134|FRESH MILK|0.2|3|HUNTER 1% CHOCOLATE MILK 14 OZ|263dfee06a448f84776d585b9451127b8e7fa9be|46.22881024317351|35.604954314503821|00074336863974|MILK|DAIRY|-80.837892|80.841348801086681|258|2
35.17739|d913077e0ce8e7dec5e0bc8102e222f50ddcc94a|6.39|2014-09-22 20:25:00|80.801203185414451|1|4154800385|208|35.195441956916255|0|24|252|-80.825175|45|35.152722|PREMIUM ICE CREAM|1.61|5|EDY'S SLOW CHURNED CHOC CHIP|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00041548766867|ICE CREAM|FROZEN|-80.80146|80.801468041191526|160|1
35.17739|e1dac7ad1ff0604419c175371285a07881afba6b|6.39|2014-12-28 10:49:00|80.801203185414451|1|4154800385|208|35.195441956916255|0|24|252|-80.825175|45|35.152722|PREMIUM ICE CREAM|1.51|5|EDY'S SLOW CHURNED CHOC CHIP|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00041548766867|ICE CREAM|FROZEN|-80.80146|80.801468041191526|160|1
35.17739|b062f0bed4c6645edd1f68bd919283da04edd5a6|6.39|2015-01-31 17:17:00|80.801203185414451|1|4154800385|208|35.195441956916255|0|24|252|-80.825175|45|35.152722|PREMIUM ICE CREAM|1.51|5|EDY'S SLOW CHURNED CHOC CHIP|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00041548766867|ICE CREAM|FROZEN|-80.80146|80.801468041191526|160|1
35.17739|01190aa0edffd9a15572cd7935c107d3e13b187a|13.29|2014-11-01 14:37:00|80.801203185414451|1|3700013882|208|35.195441958045173|0|24|389|-80.844274|66|35.204336|NFS-LAUNDRY DETERGENTS|1.3|1|TIDE HE ORIGINAL 64 LD|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00037000088868|DETERGENTS|G1 GROCERY|-80.80146|80.801461908030433|61|1
35.17739|7b34da95e301219ca193498d87cb7eb2d9c761e6|2.79|2015-01-04 14:55:00|80.801203185414451|1|3800035900|208|35.195441957608423|0|24|41|-80.85013|6|35.175855|BREAKFAST BARS|0.0|1|KLGS NUTRI GRN BAR BLUEBERRY|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00038000357008|BREAKFAST FOODS|G1 GROCERY|-80.80146|80.801465219970751|218|1
35.17739|6b06876437e96921ae3d8a1927eb16df0629b70e|3.89|2014-11-11 11:41:00|80.801203185414451|1|3800043426|208|35.195441957608423|0|24|42|-80.85013|6|35.175855|GRANOLA/YOGURT BARS|0.89|1|KLG FIBER+ BAR CHOC PB|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00038000490460|BREAKFAST FOODS|G1 GROCERY|-80.80146|80.801465219970751|218|1
35.17739|c5f9e65de75ba453d4323644c863ff40bb670a4e|2.19|2015-01-08 13:53:00|80.801203185414451|1|4900005010|208|35.195441956916255|0|24|55|-80.825175|8|35.152722|REGULAR|0.94|23|MM LEMONADE 2 LITER|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00025000053818|CARBONATED BEVERAGES|BEVERAGE|-80.80146|80.801468041191526|160|1
35.17739|a8632cb71e8bd82d6bb2072c9369c4b2f68ac2ae|10.99|2014-09-30 20:58:00|80.801203185414451|1|2200012357|208|35.195441957608423|0|24|727|-80.85013|7|35.175855|SEASONAL CANDY-SINGLE FAC|1.1|1|I/O(H14)SWEET VS SOUR 95CT|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00022000123572|CANDY|G1 GROCERY|-80.80146|80.801465219970751|218|1
35.17739|2b3a88a34f079e933ca9311a9611800337694eef|4.29|2014-11-03 13:52:00|80.801203185414451|1|2840006399|208|35.195441958060485|0|24|204|-80.826724|31|35.195689|TORTILLA CHIPS|1.79|1|TOSTITOS RESTURANT STYLE PP|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00028400063999|SNACKS|G1 GROCERY|-80.80146|80.801461677209588|412|1
35.17739|875a220b60b7a51f0fd83b0798f82f7941f38f04|6.99|2015-01-25 16:35:00|80.801203185414451|1|2066200530|208|35.195441958045173|0|24|254|-80.844274|892|35.204336|PREMIUM PIZZA|1.0|5|NEWMANS FOUR CHEESE PIZZA|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00020662005311|FROZEN PIZZA|FROZEN|-80.80146|80.801461908030433|61|1
35.17739|9da55390118fa88b3c0b26ed25eb98a0f9bc05f3|4.89|2014-12-03 21:24:00|80.801203185414451|1|1600027529|208|35.195441956916255|0|24|74|-80.825175|9|35.152722|RTE CEREAL ALL FAMILY|0.0|1|GM BASIC 4|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00016000275362|CEREAL|G1 GROCERY|-80.80146|80.801468041191526|160|1
35.17739|fdad54d78a45cdc85c52dd89b3a28fbbf3d45d49|6.99|2015-02-16 15:56:00|1.4094857484078087|1|2066200530|208|0.613961277758128|0|26|254|-80.80146|892|35.17739|PREMIUM PIZZA|0.0|5|NEWMANS FOUR CHEESE PIZZA|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|0.61471665291522548|00020662005311|FROZEN PIZZA|FROZEN|-80.80146|1.4102515174184975|208|1
35.17739|e3612016c5498cbd9c3b757b476d3f1a7e7a3b30|2.99|2014-12-28 15:38:00|80.801203185414451|1|2066200002|208|35.195441956916255|0|24|184|-80.825175|28|35.152722|SALAD DRESSINGS-LIQUID|0.0|1|NEWMANS DRS VIN BALSAMIC|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00020662000064|SALAD DRESSING/MAYONNAISE|G1 GROCERY|-80.80146|80.801468041191526|160|1
35.17739|911310151858786d1a7c550ff441503e2f6222c2|4.89|2014-12-08 10:48:00|80.801203185414451|1|1600027529|208|35.195441958045173|0|24|74|-80.844274|9|35.204336|RTE CEREAL ALL FAMILY|0.0|1|GM BASIC 4|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00016000275362|CEREAL|G1 GROCERY|-80.80146|80.801461908030433|61|1
35.17739|8f2630d41b42f865e9c4f4f67cf1d4aeeb372746|6.99|2014-12-15 16:28:00|80.801203185414451|1|2066200530|208|35.195441958045173|0|24|254|-80.844274|892|35.204336|PREMIUM PIZZA|1.99|5|NEWMANS FOUR CHEESE PIZZA|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00020662005311|FROZEN PIZZA|FROZEN|-80.80146|80.801461908030433|61|1
35.17739|4df7a41ba33d1a3d216b8980f38da8c22a342b09|4.89|2014-12-12 11:16:00|80.801203185414451|1|1600027529|208|35.195441958060485|0|24|74|-80.826724|9|35.195689|RTE CEREAL ALL FAMILY|0.0|1|GM BASIC 4|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00016000275362|CEREAL|G1 GROCERY|-80.80146|80.801461677209588|412|1
35.17739|7ae6aa1aa78d0047a497af0a32660349252fac12|4.89|2014-09-11 12:23:00|1.4094857484078087|1|1600027529|208|0.613961277758128|0|26|74|-80.80146|9|35.17739|RTE CEREAL ALL FAMILY|0.0|1|GM BASIC 4|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|0.61471665291522548|00016000275362|CEREAL|G1 GROCERY|-80.80146|1.4102515174184975|208|1
35.17739|1ed4e37d3623f9904dfc056c0c22973be8c195d4|4.89|2014-11-19 15:03:00|80.801203185414451|1|1600027529|208|35.195441958060485|0|24|74|-80.826724|9|35.195689|RTE CEREAL ALL FAMILY|0.0|1|GM BASIC 4|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00016000275362|CEREAL|G1 GROCERY|-80.80146|80.801461677209588|412|1
35.17739|c84790eb5295c1208341bf777c8f8f4496a5d61a|4.59|2015-03-01 15:41:00|80.801203185414451|1|2430009001|208|35.195441956916255|0|24|1433|-80.825175|9|35.152722|GRANOLA|0.0|1|HEARTLAND ORIGINAL GRANOLA|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00024300090011|CEREAL|G1 GROCERY|-80.80146|80.801468041191526|160|1
35.17739|8136cc182366b9644e2c2c24e0470fe3e8b6c82e|4.89|2014-09-25 19:35:00|80.801203185414451|1|1600027529|208|35.195441957608423|0|24|74|-80.85013|9|35.175855|RTE CEREAL ALL FAMILY|0.0|1|GM BASIC 4|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00016000275362|CEREAL|G1 GROCERY|-80.80146|80.801465219970751|218|1
35.17739|565b2e47e10ebea7e6a8c00f68450897952e4289|4.89|2015-03-03 15:34:00|80.801203185414451|1|1600027529|208|35.195441958060485|0|24|74|-80.826724|9|35.195689|RTE CEREAL ALL FAMILY|0.0|1|GM BASIC 4|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00016000275362|CEREAL|G1 GROCERY|-80.80146|80.801461677209588|412|1
35.17739|c29e67bc7aeb9e4ba3829e2dee3c5a00adaaf6ca|4.89|2014-12-30 19:06:00|80.801203185414451|1|1600027529|208|35.195441956916255|0|24|74|-80.825175|9|35.152722|RTE CEREAL ALL FAMILY|0.0|1|GM BASIC 4|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00016000275362|CEREAL|G1 GROCERY|-80.80146|80.801468041191526|160|1
35.17739|d45903c1a822c8fe39855fbaf702acc38ad2c755|6.99|2014-12-18 15:33:00|80.801203185414451|1|7981306060|208|35.19544195666824|0|24|2021|-80.810056|505|35.219587|FRESH CHEESE|3.5|6|BOURSIN SPINACH & ART. CUP|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00079813060631|SPECIALTY CHEESE|DELI|-80.80146|80.801468835515195|401|1
35.17739|b71b55f835f2405666db16c4f0eddd6fdaf690b8|8.49|2014-11-10 07:22:00|80.801203185414451|1||208|35.195441956916255|0|24|503|-80.825175|64|35.152722|FRESH GRAPES|2.07|4|RED GRAPES,SEEDLESS 12/16|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00204023000003|FRESH PRODUCE|PRODUCE|-80.80146|80.801468041191526|160|1
35.17739|f903f72b3c33d0daac71d65280f9599cf242df9c|5.15|2015-01-13 15:45:00|80.801203185414451|1|20128900000|208|35.195441958045173|0|24|297|-80.844274|49|35.204336|GROUND BEEF|0.0|2|VALUE PK HT PREMIUM GROUND BF|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00201289000006|BEEF|MEAT|-80.80146|80.801461908030433|61|1
35.17739|a878a92d378f21ca7a11b5a6528a4d2d9f02fcec|5.56|2014-10-24 08:45:00|80.801203185414451|1||208|35.195441958045173|0|24|503|-80.844274|64|35.204336|FRESH GRAPES|0.37|4|RED GRAPES,SEEDLESS 12/16|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00204023000003|FRESH PRODUCE|PRODUCE|-80.80146|80.801461908030433|61|1
35.17739|975f2b80c2bd3c3cf61f8a8c43a90bc370b875e9|2.04|2015-01-20 16:40:00|1.4094857484078087|1||208|0.613961277758128|0|26|500|-80.80146|64|35.17739|FRESH APPLES|0.0|4|GOLD DEL APPLE EASTERN|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|0.61471665291522548|00204137000005|FRESH PRODUCE|PRODUCE|-80.80146|1.4102515174184975|208|1
35.17739|e889e212b38903307ece0a7b1bc3b5e604df183d|2.79|2014-11-16 15:50:00|80.801203185414451|1|4144930022|208|35.195441956916255|0|24|8|-80.825175|2|35.152722|BROWNIE MIXES|0.0|1|GHIRADELLI TRIPL FUDGE BROWNIE|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00041449302706|BAKING MIXES|G1 GROCERY|-80.80146|80.801468041191526|160|1
35.17739|f48835481ec8057936317a7877647f3c8727aadc|8.58|2015-01-01 19:10:00|80.801203185414451|1|3700046967|208|35.195441956916255|0|24|3990|-80.825175|1080|35.152722|ORAL HYGIENE DENTAL FLOS|2.6|17|(JHK) GLIDE DENTAL FLOSS MNT|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00037000469568|ORAL HYGIENE|HBC|-80.80146|80.801468041191526|160|2
35.17739|9049279f275b77bfded9eabb43281e85a14067ac|3.49|2014-11-16 09:54:00|80.801203185414451|1|7760750649|208|35.195441958060485|0|24|1013|-80.826724|207|35.195689|SPECIALTY SEAS GROCERY 1|0.99|1|NOEL ADVENT CALENDARS|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00077607506495|SPECIALTY-SEASONAL|G1 GROCERY|-80.80146|80.801461677209588|412|1
35.17739|b2509da706bbb8b32776d0909873c5c4b204065f|7.98|2015-02-25 14:16:00|80.801203185414451|1|7341001375|208|35.195441956916255|0|24|1027|-80.825175|162|35.152722|GRAIN|1.99|7|ARNOLD OATNUT WP BRD PP|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00073410013557|SLICED BREAD|COMMERCIAL BAKERY|-80.80146|80.801468041191526|160|2
35.17739|cb0cedbe55b3c512e0673cd4adf73497f1abe9f8|8.58|2014-10-05 11:58:00|80.801203185414451|1|7341001375|208|35.195441956916255|0|24|1027|-80.825175|162|35.152722|GRAIN|2.14|7|ARN HEALTHNUT BRD WP PP|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00073410013656|SLICED BREAD|COMMERCIAL BAKERY|-80.80146|80.801468041191526|160|2
35.17739|11f6c83a3f636d29b4f65341c28a5e6b99778ed3|3.99|2015-02-13 15:23:00|80.801203185414451|1|7341001375|208|35.195441958045173|0|24|1027|-80.844274|162|35.204336|GRAIN|0.0|7|ARN HEALTHNUT BRD WP PP|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00073410013656|SLICED BREAD|COMMERCIAL BAKERY|-80.80146|80.801461908030433|61|1
35.17739|7245edc2511019b5f180f8c4257cf45692caeb25|3.29|2014-12-17 22:32:00|80.801203185414451|1|7373108300|208|35.195441958045173|0|24|204|-80.844274|31|35.204336|TORTILLA CHIPS|0.0|1|MISSION TORTILLA STRIPS|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00073731081037|SNACKS|G1 GROCERY|-80.80146|80.801461908030433|61|1
35.17739|11ac8a977115ca793b028f0b37b10b8368d8b802|2.99|2015-02-14 17:24:00|80.801203185414451|1|68725002611|208|35.195441956916255|0|24|1982|-80.825175|480|35.152722|DRY GOODS CRACKERS|0.0|6|DIVINA FRENCH MINI TOAST|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00687250026112|DRY GOODS|DELI|-80.80146|80.801468041191526|160|1
35.17739|ed92e36cea68881bc12b45e29c1f057f1243e205|7.68|2014-09-24 10:04:00|80.801203185414451|1||208|35.195441956916255|0|24|503|-80.825175|64|35.152722|FRESH GRAPES|1.54|4|GREEN GRAPES, SEEDLESS 12/16|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00204022000004|FRESH PRODUCE|PRODUCE|-80.80146|80.801468041191526|160|1
35.17739|7a311d4a4325b9528d0575878ec2a940f1d2b67f|1.31|2014-10-21 18:40:00|80.801203185414451|1||208|35.195441956916255|0|24|502|-80.825175|64|35.152722|FRESH BANANAS|0.0|4|BANANAS, YELLOW|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00204011000008|FRESH PRODUCE|PRODUCE|-80.80146|80.801468041191526|160|1
35.17739|d6b132bdd080e5fa9336597d7c15eb242282b07b|1.21|2014-09-30 16:16:00|80.801203185414451|1||208|35.195441958060485|0|24|502|-80.826724|64|35.195689|FRESH BANANAS|0.0|4|BANANAS, YELLOW|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00204011000008|FRESH PRODUCE|PRODUCE|-80.80146|80.801461677209588|412|1
35.17739|d751cef4951f936cec093b299980ba15c3cf2cb1|1.37|2014-09-30 07:45:00|80.801203185414451|1||208|35.195441956916255|0|24|502|-80.825175|64|35.152722|FRESH BANANAS|0.0|4|BANANAS, YELLOW|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00204011000008|FRESH PRODUCE|PRODUCE|-80.80146|80.801468041191526|160|1
35.17739|f4f8b53262f6c7121ef6fe1dea0f3a7faeec41c6|1.07|2015-02-19 10:37:00|80.801203185414451|1||208|35.195441958045173|0|24|502|-80.844274|64|35.204336|FRESH BANANAS|0.0|4|BANANAS, YELLOW|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00204011000008|FRESH PRODUCE|PRODUCE|-80.80146|80.801461908030433|61|1
35.17739|e3b14ded35b97e764ac5cc9b7fbe7e9b66fb59a0|8.67|2014-10-22 19:44:00|80.801203185414451|1|7203631051|208|35.195441958060485|0|24|192|-80.826724|30|35.195689|COOKING SPRAYS|2.67|1|HT COOKING SPRAY EXT OLIVE OIL|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00072036310521|SHORTENING/OIL|G1 GROCERY|-80.80146|80.801461677209588|412|3
35.17739|d7c777b55d132d782223fa57c306c1debd46be9b|3.97|2014-10-17 11:56:00|80.801203185414451|1|7203659020|208|35.195441958045173|0|24|312|-80.844274|51|35.204336|BUTTER|0.0|3|HARRIS TEETER UNSALTED BUTTER|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00072036590213|BUTTER & MARGARINE|DAIRY|-80.80146|80.801461908030433|61|1
35.17739|91cdefad7e118ded34b70240c77ef5c3f54a0468|3.39|2014-11-12 20:55:00|80.801203185414451|1|2529300098|208|35.195441956916255|0|24|1265|-80.825175|57|35.152722|ALMOND MILK|0.0|3|SILK PURE ALMOND UNSWEETEN VAN|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00025293001367|MILK|DAIRY|-80.80146|80.801468041191526|160|1
35.17739|7493bc2bd0dc55a4643f62c23cdf32fb02f3a340|3.34|2014-11-23 11:18:00|80.801203185414451|1|3600025824|208|35.195441956804878|0|24|424|-80.849471|72|35.161696|NFS-FACIAL TISSUE|0.84|1|KLEENEX FACIAL TIS UPRIGHT AST|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00036000374032|PAPER/PLASTIC PRODUCTS|G1 GROCERY|-80.80146|80.801468407184188|35|2
35.17739|e23d98d5528fdeb5465b060c0a1e30eba5a4cc8a|7.98|2015-02-27 07:37:00|80.801203185414451|1|69499008364|208|35.195441956916255|0|24|1250|-80.825175|12|35.152722|SPECIALTY COOKIES|0.98|1|LU LE PETITE ECOLIER XDK CHOC|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00694990013500|COOKIES|G1 GROCERY|-80.80146|80.801468041191526|160|2
35.17739|a8e2231cd114bb64f809f298ca6da4ae7a647457|1.5|2014-11-19 17:51:00|80.801203185414451|1|7203663107|208|35.195441956916255|0|24|1262|-80.825175|57|35.152722|HALF N HALF WHIPPING CREAM|0.0|3|HT HALF & HALF|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00072036632036|MILK|DAIRY|-80.80146|80.801468041191526|160|1
35.17739|6ae528fdef60a0dd517216e2ca223adf85fe3e12|4.79|2015-02-08 14:19:00|80.801203185414451|1|2100001860|208|35.195441957608423|0|24|331|-80.85013|52|35.175855|NATURAL SLICED|0.5|3|CRACKER BARRELL HAVARITI|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00021000018482|CHEESE|DAIRY|-80.80146|80.801465219970751|218|1
35.17739|a819864c803a9ebb08010e0d284e21cc577913ea|1.29|2014-11-11 12:41:00|80.801203185414451|1|8379152001|208|35.195441956916255|0|24|1981|-80.825175|480|35.152722|CHIPS|0.0|6|DIRTY POT CHIP LIGHTLY SALTED|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00083791520018|DRY GOODS|DELI|-80.80146|80.801468041191526|160|1
35.17739|257d3f34457c1f8bf6cff382802267c88b9c007d|5.99|2015-02-09 14:20:00|80.801203185414451|1|74759931462|208|35.195441957608423|0|24|727|-80.85013|7|35.175855|SEASONAL CANDY-SINGLE FAC|1.0|1|I/O(V15)CARAMEL TRIC|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00747599314629|CANDY|G1 GROCERY|-80.80146|80.801465219970751|218|1
35.17739|f3dbcaeb2f52fa79d7d5f1546f37bc28ecc018d6|3.39|2014-12-04 20:42:00|80.801203185414451|1|2529300098|208|35.195441957608423|0|24|1265|-80.85013|57|35.175855|ALMOND MILK|0.4|3|SILK PURE ALMOND DARKCHOCOLATE|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00025293001190|MILK|DAIRY|-80.80146|80.801465219970751|218|1
35.17739|b91c3b4fc3bc357baa263e2aed5efc31292066a7|13.99|2014-09-12 20:47:00|80.801203185414451|1|1626400786|208|35.195441956916255|0|24|1661|-80.825175|381|35.152722|ICE CREAM BRANDED|6.0|14|CARVEL LIL LOVE IC CAKE|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00016264007860|CAKES|BAKERY|-80.80146|80.801468041191526|160|1
35.17739|62572347e99fea7ecfca4d3780468fdf3195ad2e|12.49|2014-12-18 17:32:00|80.801203185414451|1|6206704955|208|35.195441956916255|0|24|459|-80.825175|83|35.152722|IMPORT BEER|0.0|16|LABATT'S BLUE LT 12PK BOTTLES|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00062067049552|IMPORT BEER|BEER|-80.80146|80.801468041191526|160|1
35.17739|eec066b352b39ac3cad7eeec0b54b90362af40b3|12.49|2014-10-09 17:27:00|80.801203185414451|1|6206704955|208|35.195441956916255|0|24|459|-80.825175|83|35.152722|IMPORT BEER|0.0|16|LABATT'S BLUE LT 12PK BOTTLES|2ddc277529c779354425e14adc6ea7effd4c5242|1.247346711657224|35.194272495053255|00062067049552|IMPORT BEER|BEER|-80.80146|80.801468041191526|160|1
34.977331|885d4d335498409fa6b791e840d7c999be4c4d73|1.94|2014-12-16 21:06:00|1.41290891556208|4|7203698254|149|0.6104695895098807|0|33|115|-81.027334|16|34.977331|REMAINING FRUIT|0.0|1|HT PINEAPPLE CRUSHED JC 20|30b1278253476adbcf4d5571180503d56a7f8aba|2.288476636401017|0.61055446569467375|00072036982520|FRUIT-CAN/JAR|G1 GROCERY|-81.027334|1.4141937624131469|149|2
35.103409|3bb1dc6867fdb378d0b6d992f4886e736c1f1baa|1.49|2015-01-23 11:40:00|80.992192682720116|3|2840002819|88|35.113861127407084|0|56|206|-80.85753|31|35.116638|FRONT END SNACKS|0.0|1|BAKED LAYS|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|35.113093007298254|00028400032087|SNACKS|G1 GROCERY|-80.992182|80.992191520780622|204|1
35.103409|470fa20a33912976a4745a3002493fc2cff1a4f8|1.49|2015-01-02 11:34:00|80.992192682720116|3|2840002819|88|35.113861127407084|0|56|206|-80.85753|31|35.116638|FRONT END SNACKS|0.0|1|BAKED LAYS|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|35.113093007298254|00028400032087|SNACKS|G1 GROCERY|-80.992182|80.992191520780622|204|1
35.103409|868cd0988bd52ce055bdb6dcf79e8483b2cce71d|1.49|2015-01-29 11:34:00|80.992192682720116|3|2840002819|88|35.113861127407084|0|56|206|-80.85753|31|35.116638|FRONT END SNACKS|0.0|1|BAKED LAYS|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|35.113093007298254|00028400032087|SNACKS|G1 GROCERY|-80.992182|80.992191520780622|204|1
35.103409|e81f311c67eb55cd540700000ed99e1e2cd692ac|7.99|2015-01-06 18:32:00|1.4132775322775095|3|3114252685|88|0.6126700657242101|0|58|2019|-80.992182|505|35.103409|PRESSED COOKED CHEESE|3.0|6|BELGIOISO ROMANO WEDGE|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00031142526851|SPECIALTY CHEESE|DELI|-80.992182|1.413580244274486|88|1
35.103409|c0a7a2e41ca4213af923a78599665439ccbe6a6d|4.99|2014-10-10 10:22:00|1.4132775322775095|3|2840008313|88|0.6126700657242101|0|58|204|-80.992182|31|35.103409|TORTILLA CHIPS|1.0|1|TOSTITOS RSTC FAMILY SIZE|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00028400083133|SNACKS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|876a8033a49beda06acf4ee314f31f1d4e198880|1.42|2015-01-20 18:03:00|1.4132775322775095|3||88|0.6126700657242101|0|58|502|-80.992182|64|35.103409|FRESH BANANAS|0.0|4|BANANAS, YELLOW|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00204011000008|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|1
35.103409|3a1fe11f6e6ccb54c3ca5fa7b3cb3e9b7a426a79|4.29|2014-12-30 16:06:00|1.4132775322775095|3|2840016014|88|0.6126700657242101|0|58|201|-80.992182|31|35.103409|POTATO CHIPS|0.29|1|LAYS HONEY BBQ|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00028400160537|SNACKS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|d5322a90ea29d72b0d908a1c619cc97e16495cdf|3.49|2014-12-26 11:17:00|80.992192682720116|3|2840008294|88|35.113861097757884|0|56|201|-80.945176|31|35.323246|POTATO CHIPS|0.99|1|LAYS KETTLE SALT & VINEGAR|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|35.113093007298254|00028400082921|SNACKS|G1 GROCERY|-80.992182|80.992213886969296|166|1
35.103409|e1dff2ecabce7fff30c05fcb03ef243ad0adab5a|4.35|2015-03-07 18:10:00|1.4132775322775095|3|2840003282|88|0.6126700657242101|0|58|199|-80.992182|31|35.103409|DIPS & SALSAS|0.0|1|TOSTITOS MED SALSA|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00028400032827|SNACKS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|cbf56a792bf27d573caf209467411d59a6fe4b0b|2.59|2015-01-24 18:03:00|1.4132775322775095|3|1480000034|88|0.6126700657242101|0|58|128|-80.992182|20|35.103409|APPLE JUICE-SHELF|0.0|1|MOTTS FOR TOTS APPLE JUICE|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00014800318203|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|8b68ec86291a1c154b2c42a05990d8d9e3c35413|1.89|2014-12-27 14:10:00|80.992192682720116|3|4850001775|88|35.113861097757884|0|56|335|-80.945176|56|35.323246|ORANGE JUICE-REGRIGERATED|0.0|3|TROPICANA PP CALCIUM 12 OZ|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|35.113093007298254|00048500017760|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.992182|80.992213886969296|166|1
35.103409|662a2fd6474b76bee2ba1c74d63c21f448ff1e31|6.49|2015-02-25 13:32:00|1.4132775322775095|3|7841112105|88|0.6126700657242101|0|58|350|-80.992182|196|35.103409|FROZEN PASTA|0.0|5|CAESARS PASTA GF STUFFED SHELL|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00078411121058|PASTA-FROZEN|FROZEN|-80.992182|1.413580244274486|88|1
35.103409|3abda53692bcac9d008f11bacca4b638677d45fd|4.49|2014-10-28 19:35:00|1.4132775322775095|3|81651201038|88|0.6126700657242101|0|58|141|-80.992182|21|35.103409|TRAIL MIXES AND BLENDS|0.0|1|CR SN MILK CHOC PRETZELS|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00816512010389|NUTS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|d5305c49e6aa24324aefc04e65069f9207bef50b|8.38|2014-11-02 20:58:00|1.4132775322775095|3|3800031846|88|0.6126700657242101|0|58|81|-80.992182|9|35.103409|RTE CEREAL KIDS|0.0|1|KELL COCOA KRISPIES|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00038000768620|CEREAL|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|9a7730f1590162f927156ebeb2adc08a0e870e9d|2.0|2014-09-27 20:08:00|1.4132775322775095|3||88|0.6126700657242101|0|58|511|-80.992182|64|35.103409|FRESH AVOCADOS|0.0|4|AVOCADOS, HASS XL 36CT|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00204770000004|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|1
35.103409|451daea3b50b1b921a987d0f522ef46c72a1a6a6|1.0|2014-12-28 13:28:00|80.992192682720116|3|4000000435|88|35.113861076899745|0|56|47|-80.780702|7|35.318911|REGISTER BARS|0.0|1|(FE)SNICKERS CANDY BAR|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|35.113093007298254|00040000424314|CANDY|G1 GROCERY|-80.992182|80.992222844945303|167|1
35.103409|ea9d2947c9f3361d88bb55eca4d35fa96ce85938|2.09|2015-01-14 18:36:00|1.4132775322775095|3||88|0.6126700657242101|0|58|542|-80.992182|64|35.103409|FRESH VEGETABLES REMAIN|0.0|4|COO BOK CHOY|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00204545000000|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|1
35.103409|04e77751579888f7cc8d8be0919efe5f78a7a0ed|3.34|2015-02-10 17:10:00|1.4132775322775095|3|7203643010|88|0.6126700657242101|0|58|252|-80.992182|45|35.103409|PREMIUM ICE CREAM|0.0|5|HT PREM CHOCOLATE IC|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00072036430113|ICE CREAM|FROZEN|-80.992182|1.413580244274486|88|1
35.103409|84f14eacc4ddf3d429fc9ca3e2cf8e7e958e68dd|3.29|2014-11-05 12:03:00|80.992192682720116|3|2840018382|88|35.113861127407084|0|56|201|-80.85753|31|35.116638|POTATO CHIPS|0.0|1|BAKED LAYS BBQ|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|35.113093007298254|00028400183833|SNACKS|G1 GROCERY|-80.992182|80.992191520780622|204|1
35.103409|da676c686901fed7989f5fd0d65f242be0f8f239|1.69|2014-12-06 13:54:00|1.4132775322775095|3|7203617992|88|0.6126700657242101|0|58|5618|-80.992182|1512|35.103409|RUBBER/HOUSEHOLD GLOVES|0.0|18|(PPL) (JHK) HT LATEX GLVES MED|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00072036179920|BROOMS/MOPS & BRUSHES|GM|-80.992182|1.413580244274486|88|1
35.103409|7809559da0d35ae763b18df6a6c2bca598f73b12|1.49|2015-01-04 13:26:00|80.992192682720116|3|2840002819|88|35.113861076899745|0|56|206|-80.780702|31|35.318911|FRONT END SNACKS|0.0|1|LAYS SALT & VINEGAR|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|35.113093007298254|00028400032575|SNACKS|G1 GROCERY|-80.992182|80.992222844945303|167|1
35.103409|1003fa2169f7d2da3311bb3cd3bd82d285a73816|5.1|2014-12-21 21:08:00|1.4132775322775095|3|4156514116|88|0.6126700657242101|0|58|1211|-80.992182|272|35.103409|HISP SALSA/DIPS|1.1|1|PACE T&C SALSA HOT|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00041565142163|HISPANIC PREP. FOODS|G1 GROCERY|-80.992182|1.413580244274486|88|2
35.103409|3158e0fb5514371c330b3c290e979d87a4a7d214|6.79|2014-11-17 19:46:00|1.4132775322775095|3|4850001833|88|0.6126700657242101|0|58|335|-80.992182|56|35.103409|ORANGE JUICE-REGRIGERATED|0.8|3|TROPICANA CALCIUM ORANGE JUICE|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00048500018309|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|49563a1034dcf36a9c13bb33752ad6a043463e7f|6.38|2014-11-16 00:44:00|1.4132775322775095|3||88|0.6126700657242101|0|58|562|-80.992182|64|35.103409|FRESH CUT FRUIT|0.0|4|MIXED FRUIT (IN-STORE)|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00204472000005|FRESH PRODUCE|PRODUCE|-80.992182|1.413580244274486|88|1
35.103409|fe32a440610268b092758dbdaefb6b3ec21ccf99|5.99|2015-03-01 15:55:00|80.992192682720116|3|2301200343|88|35.113861076899745|0|56|1477|-80.780702|485|35.318911|SUSHI HYBRID|0.0|6|Sushi Volcano|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|35.113093007298254|00023012003432|SUSHI|DELI|-80.992182|80.992222844945303|167|1
35.103409|c84784ef4c0e73b73936b2599ce809654d05e6c8|4.39|2014-09-10 19:45:00|1.4132775322775095|3|2446306109|88|0.6126700657242101|0|58|79|-80.992182|273|35.103409|ASIAN SAUCES/SEASONINGS|0.0|1|HUY FONG SC CHILI GARL DISPENS|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00024463061095|ASIAN PREP. FOODS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|bd6999e3658f9568092f70e8721928ab0ed4cfc6|2.69|2014-09-23 22:21:00|1.4132775322775095|3|7203663996|88|0.6126700657242101|0|58|342|-80.992182|57|35.103409|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00072036631299|MILK|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|7feeb4d522dcd0afba7f7bfc57ac805caa26c1f0|2.69|2014-09-29 21:18:00|1.4132775322775095|3|7203663996|88|0.6126700657242101|0|58|342|-80.992182|57|35.103409|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00072036631299|MILK|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|e1889725d3e01e2e65f5e9c996504d7cd143dc56|3.99|2014-11-11 16:05:00|1.4132775322775095|3|7203663995|88|0.6126700657242101|0|58|342|-80.992182|57|35.103409|FRESH MILK|0.0|3|HARRIS TEETER WHOLE MILK|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00072036639950|MILK|DAIRY|-80.992182|1.413580244274486|88|1
35.103409|83f31dcf267f4a678bb929366df6695cd1b697fc|5.49|2014-11-14 11:45:00|80.992192682720116|3|2301290132|88|35.113861127407084|0|56|1477|-80.85753|485|35.116638|SUSHI HYBRID|0.0|6|SPICY CALIFORNIA ROLL SP|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|35.113093007298254|00023012901325|SUSHI|DELI|-80.992182|80.992191520780622|204|1
35.103409|f4da8819edfd1cd1bc504dcc0b3ab1e3e2d24cfb|6.49|2014-12-07 13:10:00|80.992192682720116|3|2301200002|88|35.113861076899745|0|56|1475|-80.780702|485|35.318911|SUSHI CLASSIC|0.0|6|CALIFORNIA ROLL|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|35.113093007298254|00023012000028|SUSHI|DELI|-80.992182|80.992222844945303|167|1
35.103409|193572187811e2099293176c9414acb7412279db|4.19|2015-02-17 16:24:00|1.4132775322775095|3|2900007212|88|0.6126700657242101|0|58|1149|-80.992182|21|35.103409|PEANUTS|0.0|1|PLNTRS COCKTAIL PEANUTS|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00029000072121|NUTS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|1a70237c09fcaf4cec8e261eaede287e8af39245|3.29|2014-10-13 11:34:00|80.992192682720116|3|2840018382|88|35.113861127407084|0|56|201|-80.85753|31|35.116638|POTATO CHIPS|0.79|1|BAKED LAYS|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|35.113093007298254|00028400183826|SNACKS|G1 GROCERY|-80.992182|80.992191520780622|204|1
35.103409|ad062c75fb971717e1606612bf62db1b12cc4342|3.29|2014-09-14 12:18:00|1.4132775322775095|3|2840018382|88|0.6126700657242101|0|58|201|-80.992182|31|35.103409|POTATO CHIPS|0.0|1|BAKED LAYS|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00028400183826|SNACKS|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|b7400b6bc31913920fb6c9451cbb1c5d1422a028|3.29|2014-09-11 11:49:00|80.992192682720116|3|2840018382|88|35.113861127407084|0|56|201|-80.85753|31|35.116638|POTATO CHIPS|0.0|1|BAKED LAYS|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|35.113093007298254|00028400183826|SNACKS|G1 GROCERY|-80.992182|80.992191520780622|204|1
35.103409|811b3d037ed48fef4134ee93c74141d544652875|1.29|2015-01-15 18:22:00|1.4132775322775095|3|6414428243|88|0.6126700657242101|0|58|257|-80.992182|39|35.103409|TOMATOES|0.29|1|ROTEL TOMATOES HOT|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00064144282661|VEGETABLES-CAN/JAR|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|a7439d97afb5365fa8490753310d6c793012491b|7.99|2014-09-17 09:58:00|1.4132775322775095|3|5200020805|88|0.6126700657242101|0|58|171|-80.992182|20|35.103409|ISOTONIC DRINKS|2.99|1|GATORADE ORANGE 8PK|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00052000208078|JUICES/DRINKS-SHELF STABLE|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|7d0ed91c8c1d3f605fcb7de0be1f390dd639202e|6.57|2015-02-12 10:50:00|1.4132775322775095|3|4900005010|88|0.6126700657242101|0|58|55|-80.992182|8|35.103409|REGULAR|0.8500000000000001|23|CLASSIC COKE 2 LT CONTOUR|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00049000050103|CARBONATED BEVERAGES|BEVERAGE|-80.992182|1.413580244274486|88|3
35.103409|4b1ca538b48126b397dc7fe565f7ac3f6960734c|1.59|2014-11-19 20:40:00|1.4132775322775095|3|38137009217|88|0.6126700657242101|0|58|3990|-80.992182|1080|35.103409|ORAL HYGIENE DENTAL FLOS|0.0|17|J&J DENT FLOSS MINT WAX -09217|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00381370092179|ORAL HYGIENE|HBC|-80.992182|1.413580244274486|88|1
35.103409|cebeb32f0831dcadeb15cdbd08edb9d0be24730a|1.69|2015-01-25 11:27:00|80.992192682720116|3|4900000044|88|35.113861076899745|0|56|55|-80.780702|8|35.318911|REGULAR|0.0|23|CB COKE SINGLE 20 OZ.|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|35.113093007298254|00049000000443|CARBONATED BEVERAGES|BEVERAGE|-80.992182|80.992222844945303|167|1
35.103409|9540fb51af31bc984c57de8f196d21b1d5ebffd6|6.57|2015-02-14 15:12:00|80.992192682720116|3|4900005010|88|35.113861065530969|0|56|54|-80.995484|8|35.444064|DIET|0.8500000000000001|23|COKE ZERO 2 LITER|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|35.113093007298254|00049000050141|CARBONATED BEVERAGES|BEVERAGE|-80.992182|80.992226982524201|121|3
35.103409|eb4a0381f028a88855762eb19cbabbeabc8190ea|1.69|2014-12-17 10:56:00|1.4132775322775095|3|4900000044|88|0.6126700657242101|0|58|55|-80.992182|8|35.103409|REGULAR|0.0|23|CB COKE SINGLE 20 OZ.|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00049000000443|CARBONATED BEVERAGES|BEVERAGE|-80.992182|1.413580244274486|88|1
35.103409|9e667430f4fab31847840dbcadc132835153c587|7.49|2014-12-17 10:55:00|1.4132775322775095|3|7203695788|88|0.6126700657242101|0|58|1403|-80.992182|389|35.103409|THAW AND SELL PIES|1.5|14|"8"" PECAN PIE"|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00072036957887|PIES|BAKERY|-80.992182|1.413580244274486|88|1
35.103409|2e8617b21772518d6bfc0dce5493b33c586fc5bb|1.79|2014-09-23 18:51:00|1.4132775322775095|3|3940001614|88|0.6126700657242101|0|58|243|-80.992182|39|35.103409|BAKED BEANS|0.0|1|BUSH BKD BEAN ORIGINAL 28|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00039400016144|VEGETABLES-CAN/JAR|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.103409|48acaaff97c2c1840a84931382441117349b07af|2.99|2015-02-27 19:58:00|1.4132775322775095|3|61300873513|88|0.6126700657242101|0|58|99|-80.992182|32|35.103409|LIQUID TEA|0.3|1|ARNOLD PALMER LITE TEA|320e6f0351e8adf9b93bcdc7fb38c77f6567d53c|0.7222169633607147|0.61177642288969325|00613008720858|SOFT DRINKS-NON-CARBONATED|G1 GROCERY|-80.992182|1.413580244274486|88|1
35.43259|fc74a2985572a4279b71e49df4aec6904ca92914|1.58|2015-01-05 17:58:00|1.4057311447477159|4|2700039005|202|0.6184153580092175|0|52|257|-80.605588|39|35.43259|TOMATOES|0.08|1|HUNTS TOMATO SAUCE BSL GAR OGN|327d6b10b7629dc663755f42fdfdd0c8e080a6e4|4.957954468528736|0.6209993146566879|00027000391037|VEGETABLES-CAN/JAR|G1 GROCERY|-80.605588|1.406832906106031|202|2
35.43259|3df497d2a205eb8b33e3aa254a8c2149d47cfe1f|3.79|2014-10-29 20:00:00|1.4057311447477159|4|1410007105|202|0.6184153580092175|0|52|1025|-80.605588|162|35.43259|WHITE|0.0|7|PEP VERY THIN WHITE BRD PP|327d6b10b7629dc663755f42fdfdd0c8e080a6e4|4.957954468528736|0.6209993146566879|00014100071051|SLICED BREAD|COMMERCIAL BAKERY|-80.605588|1.406832906106031|202|1
35.061685|f937d07085e08254e5aecda21b4852afc5dc916a|0.5|2014-12-31 01:34:00|80.994598860450068|4||475|35.076384348219754|0|53|524|-80.992182|64|35.103409|FRESH PROD FRESH ONIONS|0.0|4|COO YELLOW ONIONS, LRG|36a0a3db463d910e95e0f7e25cd96ef14ebc4f59|1.015689564750435|35.072594466811061|00204665000003|FRESH PRODUCE|PRODUCE|-80.994596|80.99460398633228|88|1
35.061685|4b3e751a528b849341af50e788792dbafb9d01bc|2.85|2014-10-21 01:47:00|80.994598860450068|4|4600028869|475|35.076384348219754|0|53|77|-80.992182|272|35.103409|HISP SAUCES/SEASONINGS|0.0|1|E  OEP SEASONING TACO|36a0a3db463d910e95e0f7e25cd96ef14ebc4f59|1.015689564750435|35.072594466811061|00046000288697|HISPANIC PREP. FOODS|G1 GROCERY|-80.994596|80.99460398633228|88|3
35.061685|338285e7d75f1cf1ff40c65c77d505714318f9ab|5.99|2014-10-21 01:45:00|80.994598860450068|4|4470007502|475|35.076384348219754|0|53|484|-80.992182|101|35.103409|BEEF WIENERS|3.0|19|OSCAR MAYER BUNLENGTH BF FRANK|36a0a3db463d910e95e0f7e25cd96ef14ebc4f59|1.015689564750435|35.072594466811061|00044700000779|WIENERS|CASE READY MEATS|-80.994596|80.99460398633228|88|1
35.061685|33bd600cb7b9fbb7c61be0e5246226b3bb18b0c0|5.29|2014-12-31 00:22:00|80.994598860450068|4|7203670779|475|35.076384348219754|0|53|4296|-80.992182|1205|35.103409|ACETAMINOPHEN|1.3|17|HT ES COOL CAPLETS|36a0a3db463d910e95e0f7e25cd96ef14ebc4f59|1.015689564750435|35.072594466811061|00072036707796|PAIN RELIEF|HBC|-80.994596|80.99460398633228|88|1
35.000049|2652fc8d795a1284ee524019ec26d654aecee6be|7.98|2014-09-18 19:37:00|1.4091206135396188|1|4850002013|249|0.6108660934093487|0|47|335|-80.699686|56|35.000049|ORANGE JUICE-REGRIGERATED|0.99|3|TROPICANA PP LOW ACID|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00048500309223|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.699686|1.4084752260255726|249|2
35.000049|882813ffbaa1b04b66b5270beeefca73edaeaaf8|4.29|2014-11-13 15:22:00|1.4091206135396188|1|4400002747|249|0.6108660934093487|0|47|91|-80.699686|13|35.000049|SPRAYED BUTTER CRACKERS|1.29|1|S RITZ SNOWFLAKE|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00044000031237|CRACKERS|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|d058b563709b729348eab39141133f7a267c1dd7|1.18|2014-12-06 16:46:00|1.4091206135396188|1|7066203001|249|0.6108660934093487|0|47|1203|-80.699686|33|35.000049|RAMEN|0.15|1|CUP O' NOODLES BEEF FLAVOR|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00070662030011|SOUP|G1 GROCERY|-80.699686|1.4084752260255726|249|2
35.000049|c21b8d450717109a0dde4e981da770db238d795a|4.99|2015-02-11 18:33:00|1.4091206135396188|1|5844977180|249|0.6108660934093487|0|47|1433|-80.699686|9|35.000049|GRANOLA|1.0|1|NAT PATH ORG GRANOLA HONEY ALM|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00058449890379|CEREAL|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|ea68fc294bdd153c41015df6c63cf691b30e7779|1.87|2014-09-26 19:07:00|1.4091206135396188|1|7203670901|249|0.6108660934093487|0|47|214|-80.699686|33|35.000049|BROTH|0.0|1|HT FF BEEF BROTH 32 OZ|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00072036709004|SOUP|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|f2dbb2f144c6bfb1a1ba913db5fda8dd3dd82a43|2.49|2015-02-16 15:47:00|1.4091206135396188|1|7203670908|249|0.6108660934093487|0|47|214|-80.699686|33|35.000049|BROTH|0.0|1|HARRIS TEETER BEEF STOCK|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00072036709103|SOUP|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|14436843c26b3497dc73371d6d614375860f813b|12.99|2014-12-20 16:49:00|1.4091206135396188|1|36382400820|249|0.6108660934093487|0|47|4216|-80.699686|1200|35.000049|DECONGEST REMEDY-ADULT|0.0|17|MUCINEX EXPCTORANT 600MG 00820|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00363824008202|COUGH/COLD/SINUS|HBC|-80.699686|1.4084752260255726|249|1
35.000049|c72ff12dca3a3db604671c355c59d1fd4de047c2|7.77|2014-10-16 16:38:00|1.4091206135396188|1||249|0.6108660934093487|0|47|1347|-80.699686|64|35.000049|PUMPKINS|0.0|4|LONG ISLAND CHEESE PUMPKIN|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00204500000007|FRESH PRODUCE|PRODUCE|-80.699686|1.4084752260255726|249|1
35.000049|e65656195bcc43b54fa5934191de933fd3cf1409|7.1|2014-11-30 17:46:00|1.4091206135396188|1|7433610102|249|0.6108660934093487|0|47|342|-80.699686|57|35.000049|FRESH MILK|2.16|3|HIGHLAND CREST WHOLE MILK|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00074336879203|MILK|DAIRY|-80.699686|1.4084752260255726|249|2
35.000049|f8a4b44a993457f60ddf9215811222d83f3b86ee|3.99|2015-01-12 19:04:00|1.4091206135396188|1|7433610006|249|0.6108660934093487|0|47|342|-80.699686|57|35.000049|FRESH MILK|0.0|3|HUNTER WHOLE MILK GALLON|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00074336100062|MILK|DAIRY|-80.699686|1.4084752260255726|249|1
35.000049|8c326363fc24131ba1bac68c75939241ae6d7512|3.55|2014-11-15 20:09:00|1.4091206135396188|1|7433610102|249|0.6108660934093487|0|47|342|-80.699686|57|35.000049|FRESH MILK|0.0|3|HIGHLAND CREST WHOLE MILK|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00074336879203|MILK|DAIRY|-80.699686|1.4084752260255726|249|1
35.000049|3b14514b36ac1899056ebe0322051e3eba70fdf7|2.99|2015-01-03 20:31:00|1.4091206135396188|1|7433610102|249|0.6108660934093487|0|47|342|-80.699686|57|35.000049|FRESH MILK|0.0|3|HIGHLAND CREST WHOLE MILK|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00074336879203|MILK|DAIRY|-80.699686|1.4084752260255726|249|1
35.000049|35b74075f1412b1232145b39a48c3d84c1e315fb|3.59|2014-10-07 16:45:00|1.4091206135396188|1|7433610102|249|0.6108660934093487|0|47|342|-80.699686|57|35.000049|FRESH MILK|0.0|3|HIGHLAND CREST WHOLE MILK|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00074336879203|MILK|DAIRY|-80.699686|1.4084752260255726|249|1
35.000049|3d5db0a1f907181d3528fd7f81d5f7120ae463ee|7.18|2014-11-26 17:37:00|1.4091206135396188|1|7342000024|249|0.6108660934093487|0|47|322|-80.699686|53|35.000049|SOUR CREAM|0.0|3|DAISY SOUR CREAM|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00073420000240|CULTURES|DAIRY|-80.699686|1.4084752260255726|249|2
35.000049|f37e4c598bd9465ac7e07bffbbdf753acf47f1de|2.99|2015-01-27 18:43:00|1.4091206135396188|1|7433610102|249|0.6108660934093487|0|47|342|-80.699686|57|35.000049|FRESH MILK|0.0|3|HIGHLAND CREST WHOLE MILK|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00074336879203|MILK|DAIRY|-80.699686|1.4084752260255726|249|1
35.000049|987d8b6328776c296340841b489673688b660cd9|6.9|2014-12-13 08:14:00|1.4091206135396188|1|7433610102|249|0.6108660934093487|0|47|342|-80.699686|57|35.000049|FRESH MILK|0.0|3|HIGHLAND CREST WHOLE MILK|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00074336879203|MILK|DAIRY|-80.699686|1.4084752260255726|249|2
35.000049|f039e3f44bc8b506039023051f2f5038b16263af|2.25|2014-10-31 08:12:00|1.4091206135396188|1|3890000407|249|0.6108660934093487|0|47|105|-80.699686|16|35.000049|FRUIT CUPS AND GELS|0.25|1|DOLE 4PK MANDRN ORANGE|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00038900042073|FRUIT-CAN/JAR|G1 GROCERY|-80.699686|1.4084752260255726|249|1
35.000049|6df6bbd875c0e52e1104e996e62bb510f13b0850|1.34|2014-10-21 17:53:00|1.4091206135396188|1|7203641111|249|0.6108660934093487|0|47|242|-80.699686|39|35.000049|CANNED BEANS|0.0|1|HT BEANS GREAT NORTHERN|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00072036411129|VEGETABLES-CAN/JAR|G1 GROCERY|-80.699686|1.4084752260255726|249|2
35.000049|d576927bce9d680b518035877ef7a02de89f1f38|2.0|2014-11-13 16:37:00|80.699698036522989|1|7464100079|249|35.025198149312338|0|18|562|-80.810056|64|35.219587|FRESH CUT FRUIT|0.0|4|APPLE CHEESE & CARMEL DIP|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|35.030887098939942|00074641000798|FRESH PRODUCE|PRODUCE|-80.699686|80.699740869428311|401|1
35.000049|2b5d9be76d95bbd36381077ac158a09183c3a6c0|0.75|2014-12-04 11:30:00|80.699698036522989|1|7653906610|249|35.025198162170462|0|18|1984|-80.844274|480|35.204336|PC CONDIMENTS|0.0|6|NATURALLY FRESH RANCH DRESSING|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|35.030887098939942|00076539066107|DRY GOODS|DELI|-80.699686|80.699731238516421|61|1
35.000049|c71258992e1c2bad35b19702c7516240bdc15ab7|3.19|2014-12-15 11:49:00|1.4091206135396188|1|3700084602|249|0.6108660934093487|0|47|3530|-80.699686|1045|35.000049|SHAMPOO-MID PRICE|0.69|17|VIDAL SASSOON SHAM SMOOTH|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00037000846659|HAIR & SCALP CARE|HBC|-80.699686|1.4084752260255726|249|1
35.000049|2efbcc174eb27f14ffbeec21b954ea32736abba6|3.5|2014-10-24 16:48:00|1.4091206135396188|1|20496000000|249|0.6108660934093487|0|47|755|-80.699686|87|35.000049|NFS-BALLOONS|0.0|9|*BALLOONS|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00204960000005|FLORAL|FLORAL|-80.699686|1.4084752260255726|249|1
35.000049|6d599b652c67c1925d8a4223f98ee2260e1c9fcf|1.49|2015-02-28 15:56:00|1.4091206135396188|1||249|0.6108660934093487|0|47|522|-80.699686|64|35.000049|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00204664000004|FRESH PRODUCE|PRODUCE|-80.699686|1.4084752260255726|249|1
35.000049|8029144917349f1a662730bc88dad0571e0ea051|15.0|2015-01-30 19:18:00|80.699698036522989|1|8130831763|249|35.025198189455452|0|18|9934|-80.699909|885|35.002628|NFS POP CHARDONNAY|0.0|13|CB-OAK CREEK CHARDONNAY|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|35.030887098939942|00081308317632|POPULAR (4-$7.99)|WINE|-80.699686|80.699686795083821|477|6
35.000049|fc40921942922d314a505fff848ffba6f9963dec|30.0|2014-10-21 17:33:00|80.699698036522989|1|8130831763|249|35.025198189455452|0|18|9934|-80.699909|885|35.002628|NFS POP CHARDONNAY|0.0|13|CB-OAK CREEK CHARDONNAY|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|35.030887098939942|00081308317632|POPULAR (4-$7.99)|WINE|-80.699686|80.699686795083821|477|12
35.000049|43505f4c5dcdc2c2519260932a043dc775cd589f|10.0|2015-02-25 13:22:00|80.699698036522989|1|8130831763|249|35.025198189455452|0|18|9934|-80.699909|885|35.002628|NFS POP CHARDONNAY|0.0|13|CB-OAK CREEK CHARDONNAY|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|35.030887098939942|00081308317632|POPULAR (4-$7.99)|WINE|-80.699686|80.699686795083821|477|4
35.000049|93d42c4f47f45ff9385bf6e7cc3687d45e14f597|6.49|2014-12-17 16:25:00|1.4091206135396188|1|73150953236|249|0.6108660934093487|0|47|3087|-80.699686|1000|35.000049|FALSE NAIL KIT-OTHER MANUF|0.0|17|KISS EVRLASTNG FRENCH-INFINITE|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00731509532401|COSMETICS|HBC|-80.699686|1.4084752260255726|249|1
35.000049|85356ca239f88e5a74459c7921792f01e3cd91ad|4.5|2014-12-24 11:55:00|1.4091206135396188|1||249|0.6108660934093487|0|47|528|-80.699686|64|35.000049|FRESH BROCCOLI|0.45|4|COO BROCCOLI CROWNS (RPC)|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00204549000006|FRESH PRODUCE|PRODUCE|-80.699686|1.4084752260255726|249|1
35.000049|ab8ceb301cb5066d6d318c2f3174198a568ba32c|4.01|2015-01-04 02:45:00|80.699698036522989|1||249|35.02519818934708|0|18|562|-80.816172|64|35.059823|FRESH CUT FRUIT|0.0|4|(SEEDLESS) WATERMELON CHUNKS|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|35.030887098939942|00204485000009|FRESH PRODUCE|PRODUCE|-80.699686|80.699688959465433|66|1
35.000049|f12493f2f7f46499280389dade4b7157d6391dc0|8.97|2014-10-23 20:26:00|80.699698036522989|1|3993805735|249|35.02519818934708|0|18|7278|-80.816172|1600|35.059823|HALLOWEEN PARTY GOODS/DECOR|2.0999999999999996|18|PUMPKIN ZIPPER BAG|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|35.030887098939942|00039938057350|SEASONAL MERCHANDISE|GM|-80.699686|80.699688959465433|66|3
35.000049|6e07fef32d4922db374c85bf3415f7aba221c9b3|4.49|2014-09-26 07:51:00|1.4091206135396188|1|4812127707|249|0.6108660934093487|0|47|1036|-80.699686|164|35.000049|BREAKFAST BAGELS|2.24|7|THOMAS' EVERYTHING  BGL 6CT PP|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|0.61242566243833529|00048121253196|BREAKFAST|COMMERCIAL BAKERY|-80.699686|1.4084752260255726|249|1
35.000049|4e309e0a940b5ee04ac7345b196439556d81645f|3.38|2014-11-11 17:51:00|80.699698036522989|1|4900000044|249|35.025197883485873|0|18|54|-80.605588|8|35.43259|DIET|0.0|23|CB COKE ZERO 20 OZ|38b65cc7a344f9ce73ab05d81f9ae501cef05043|1.7377482588364541|35.030887098939942|00049000040869|CARBONATED BEVERAGES|BEVERAGE|-80.699686|80.699837468834744|202|2
35.116638|9bd5e35d25ff054ef56013f14c27b7bf53d518dd|1.37|2014-09-20 12:52:00|80.856688219393845|4||204|35.142337291460073|0|15|561|-80.992182|64|35.103409|FR PROD ORGANIC PRODUCE|0.0|4|COO ORG RED ONIONS|3a8a98a8b95a3e7cc3a1b20ab44e2df562fe3cb0|1.7757594714353826|35.134355925261694|00294082000007|FRESH PRODUCE|PRODUCE|-80.85753|80.857553417517764|88|1
35.116638|bc7a9fc3583560be359e1458decdacb23b93916d|1.19|2014-10-25 15:55:00|80.856688219393845|4|1090063384|204|35.142337291460073|0|15|428|-80.992182|3|35.103409|NFS-BAKING CUPS|0.0|1|REYNOLDS PASTEL BAKNG CUP 50CT|3a8a98a8b95a3e7cc3a1b20ab44e2df562fe3cb0|1.7757594714353826|35.134355925261694|00010900633840|BAKING SUPPLIES|G1 GROCERY|-80.85753|80.857553417517764|88|1
35.116638|c678beb60d6684b3d4407503bf9b9046246e2a08|4.99|2015-01-02 15:53:00|80.856688219393845|4|4900002468|204|35.142337291460073|0|15|54|-80.992182|8|35.103409|DIET|1.0|23|C/F DIET COKE .5 LITER/6 PK.|3a8a98a8b95a3e7cc3a1b20ab44e2df562fe3cb0|1.7757594714353826|35.134355925261694|00049000025422|CARBONATED BEVERAGES|BEVERAGE|-80.85753|80.857553417517764|88|1
35.116638|8069c369ecfe0b7e8d5870246f96c79722e0383a|4.99|2015-01-02 16:06:00|80.856688219393845|4|4082201114|204|35.142337291460073|0|15|1878|-80.992182|435|35.103409|HUMMUS|2.49|6|GREEK OLIVE HUMMUS|3a8a98a8b95a3e7cc3a1b20ab44e2df562fe3cb0|1.7757594714353826|35.134355925261694|00040822011341|SALADS|DELI|-80.85753|80.857553417517764|88|1
35.116638|0ae92cda7002bd577a18015761a4ce65805e33e9|2.16|2014-11-15 17:38:00|80.856688219393845|4|20540500000|204|35.142337291460073|0|15|1832|-80.992182|415|35.103409|BH SLICING CHEESE|0.0|6|BR HD VERMONT CHEDDAR WHITE|3a8a98a8b95a3e7cc3a1b20ab44e2df562fe3cb0|1.7757594714353826|35.134355925261694|00205405000000|SLICING CHEESE|DELI|-80.85753|80.857553417517764|88|1
35.116638|d0122e2c40e34a8ccab2221a2b52909fb9ab9ae9|3.99|2015-01-26 12:32:00|80.856688219393845|4|2951923211|204|35.14233729509747|0|15|1687|-80.825175|385|35.152722|THAW & SELL (SWEET GOODS)|1.0|14|WW LEMON CREME SNACK|3a8a98a8b95a3e7cc3a1b20ab44e2df562fe3cb0|1.7757594714353826|35.134355925261694|00029519232177|SWEET GOODS|BAKERY|-80.85753|80.857546397398522|160|1
35.116638|da5b052639eb1640e533974f2c0932ff1777e3a3|0.69|2015-01-25 13:57:00|80.856688219393845|4|71070840284|204|35.142337291460073|0|15|580|-80.992182|136|35.103409|OTHER MERCH DRESSINGS|0.0|4|ORGANIC CAESAR DRESSING|3a8a98a8b95a3e7cc3a1b20ab44e2df562fe3cb0|1.7757594714353826|35.134355925261694|00710708402845|OTHER MERCHANDISE|PRODUCE|-80.85753|80.857553417517764|88|1
35.116638|a7571f4f507f517946d2e605ae4b034ea841bcef|0.69|2015-01-11 15:00:00|80.856688219393845|4|71070840284|204|35.142337291460073|0|15|580|-80.992182|136|35.103409|OTHER MERCH DRESSINGS|0.0|4|ORGANIC CAESAR DRESSING|3a8a98a8b95a3e7cc3a1b20ab44e2df562fe3cb0|1.7757594714353826|35.134355925261694|00710708402845|OTHER MERCHANDISE|PRODUCE|-80.85753|80.857553417517764|88|1
35.03469|9625cb47cf7d2194e2f96087a3929c765e232f46|0.66|2014-10-04 19:49:00|80.970590786568081|4||82|35.079009736394411|0|55|502|-80.994596|64|35.061685|FRESH BANANAS|0.0|4|BANANAS, YELLOW|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00204011000008|FRESH PRODUCE|PRODUCE|-80.97058|80.97058935057278|475|1
35.03469|4d10a701edc4fe60a6ec92abf86e2bdd6be3c8cf|1.0|2014-12-17 15:45:00|80.970590786568081|4|812|82|35.07900972860665|0|55|1639|-80.992182|377|35.103409|BULK (DONUTS)|0.0|14|NEW BULK DONUT CODE|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00000000008120|DONUTS|BAKERY|-80.97058|80.970613430786784|88|1
35.03469|de78e1fe560a62ff19e0457925970248401255b2|8.99|2014-12-21 17:49:00|80.970590786568081|4|78778077016|82|35.079009736394411|0|55|36|-80.994596|10|35.061685|PREMIUM GROUND|2.0|1|NEC HAZLENUT|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00787780770148|COFFEE|G1 GROCERY|-80.97058|80.97058935057278|475|1
35.03469|a48f30d4256b41d49435555a15d398908c46670f|1.0|2014-11-09 14:48:00|80.970590786568081|4|812|82|35.079009736394411|0|55|1639|-80.994596|377|35.061685|BULK (DONUTS)|0.0|14|NEW BULK DONUT CODE|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00000000008120|DONUTS|BAKERY|-80.97058|80.97058935057278|475|1
35.03469|d6ea10586fb74ec9cc23a839d14301697cc377e9|2.79|2015-01-29 13:00:00|80.970590786568081|4|5210000676|82|35.079009736394411|0|55|220|-80.994596|34|35.061685|PEPPER|0.0|1|E  MC CRUSHED RED PEPPER|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00052100006765|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.97058|80.97058935057278|475|1
35.03469|1419c4e67d3ba73b6fb839907103ab41032d174e|2.49|2014-11-02 15:12:00|80.970590786568081|4|7203688048|82|35.079009736394411|0|55|526|-80.994596|64|35.061685|FRESH MUSHROOMS|0.0|4|HT SLICED BABY BELLAS|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00072036880482|FRESH PRODUCE|PRODUCE|-80.97058|80.97058935057278|475|1
35.03469|905fddabaa016d8ad3fe9db36e842418d682576d|8.99|2014-11-22 18:11:00|80.970590786568081|4|7203695149|82|35.079009736394411|0|55|1937|-80.994596|465|35.061685|COLD PREP FOODS ENTREES|0.0|6|SPINACH & CHEESE QUICHE|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00072036951465|COLD PREPARED FOODS|DELI|-80.97058|80.97058935057278|475|1
35.03469|e377d0d5453ac35aec1b05481529627072cb0b2f|8.99|2014-09-26 14:32:00|80.970590786568081|4|7203695149|82|35.079009736394411|0|55|1937|-80.994596|465|35.061685|COLD PREP FOODS ENTREES|0.0|6|SPINACH & CHEESE QUICHE|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00072036951465|COLD PREPARED FOODS|DELI|-80.97058|80.97058935057278|475|1
35.03469|55a2898355ae2cd5dd7ab14b5aaaec4bbf11a15f|2.41|2014-12-20 13:24:00|80.970590786568081|4||82|35.079009736394411|0|55|522|-80.994596|64|35.061685|FRESH TOMATOES|0.0|4|RED HOT HOUSE TOMATO, BUNCH|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00204664000004|FRESH PRODUCE|PRODUCE|-80.97058|80.97058935057278|475|1
35.03469|bb60ab31434332a87fe3c4cdec386c2930cdcae0|1.22|2014-11-16 13:06:00|80.970590786568081|4||82|35.079009736394411|0|55|527|-80.994596|64|35.061685|FRESH CARROTS|0.0|4|COO CARROTS, BULK|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00204562000007|FRESH PRODUCE|PRODUCE|-80.97058|80.97058935057278|475|1
35.03469|1a92456e990236820aed46cafcf40aaacb1ab62c|6.99|2014-11-15 16:02:00|80.970590786568081|4|8500004528|82|35.07900972860665|0|55|9938|-80.992182|885|35.103409|NFS POP PINOT GRS/GRIGIO|0.0|13|BAREFOOT PINOT GRIGIO 4PK|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00085000045282|POPULAR (4-$7.99)|WINE|-80.97058|80.970613430786784|88|1
35.03469|58db2dfaaa47b10db6546898a8fba6466e3d02c0|0.85|2014-09-21 20:15:00|1.4132775322775095|4||82|0.6114706929155321|0|58|502|-80.97058|64|35.03469|FRESH BANANAS|0.0|4|BANANAS, YELLOW|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|0.61177642288969325|00204011000008|FRESH PRODUCE|PRODUCE|-80.97058|1.4132032182494703|82|1
35.03469|775481b47bf76dc7f8156e5ffdb3cd29ea60b65f|3.59|2014-12-16 21:49:00|80.970590786568081|4|7357000008|82|35.079009736394411|0|55|317|-80.994596|52|35.061685|CHUNK AND BAR CHEESE|1.59|3|HELUVA GOOD EXTRA SHARP|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00073570000305|CHEESE|DAIRY|-80.97058|80.97058935057278|475|1
35.03469|2e260c3961302cbd1f5bfd5e99991615811d164e|27.98|2014-12-24 09:11:00|80.970590786568081|4|8143431530|82|35.079009736394411|0|55|9962|-80.994596|887|35.061685|NFS-PREM-SAUV/FUME'BLANC|0.0|13|CB-NOBILO SAUVIGNON BLANC|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00081434315304|SUPER PREMIUM ($11-$14.99)|WINE|-80.97058|80.97058935057278|475|2
35.03469|78b6966092644f1c59a6991b2945a4bfdf3a8e58|4.29|2014-12-28 16:24:00|80.970590786568081|4|7565601754|82|35.079009736394411|0|55|6424|-80.994596|1556|35.061685|GAMES|0.0|18|ROTATING TOY|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00075656017542|TOYS|GM|-80.97058|80.97058935057278|475|1
35.03469|c11b462f468719fe739131019800a7c2a7c817be|10.0|2015-02-18 13:03:00|80.970590786568081|4|8500001444|82|35.079009736394411|0|55|9938|-80.994596|885|35.061685|NFS POP PINOT GRS/GRIGIO|0.0|13|CB-BAREFOOT PINOT GRIGIO|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00085000014448|POPULAR (4-$7.99)|WINE|-80.97058|80.97058935057278|475|2
35.03469|68dbd5f28e8d096e6c33725a0ca247318f35a1ec|3.49|2014-11-16 17:00:00|80.970590786568081|4|78142117086|82|35.07900972860665|0|55|1601|-80.992182|371|35.103409|BRANDED BREAD|0.0|14|LA BREA ASIAGO CHEESE FILONE|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00781421170861|BREAD|BAKERY|-80.97058|80.970613430786784|88|1
35.03469|7b1433c64704c7c1286f68f2d7963360b1fc642d|2.99|2014-09-22 12:36:00|80.970590786568081|4|1380004717|82|35.079009695900304|0|55|1278|-80.85753|48|35.116638|SINGLE SERVE NUTRITIONAL|0.0|5|LC SOUTHW CHICKEN PANINI|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00013800156006|FROZEN MEALS|FROZEN|-80.97058|80.970653784086934|204|1
35.03469|f2779abf4c717e1eb17e3fc9a92c2997ea8af8a5|4.98|2014-10-09 16:35:00|80.970590786568081|4|1380017219|82|35.079009695900304|0|55|1278|-80.85753|48|35.116638|SINGLE SERVE NUTRITIONAL|0.0|5|LC SPAGHETTI MEAT SAUCE|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00013800166357|FROZEN MEALS|FROZEN|-80.97058|80.970653784086934|204|2
35.03469|b8d0e5ab101ef45a364681a9844ad946f1ebbb9e|5.38|2015-01-09 16:26:00|80.970590786568081|4|1380016610|82|35.079009736394411|0|55|1278|-80.994596|48|35.061685|SINGLE SERVE NUTRITIONAL|1.38|5|LC CAFE CLSSC MEATLOAF|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00013800166951|FROZEN MEALS|FROZEN|-80.97058|80.97058935057278|475|2
35.03469|4e083d398956220d97557ea74ba854b37da49507|2.49|2014-10-06 11:29:00|80.970590786568081|4|1380017219|82|35.079009695900304|0|55|1278|-80.85753|48|35.116638|SINGLE SERVE NUTRITIONAL|0.49|5|LC SPAGHETTI MEAT SAUCE|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00013800166357|FROZEN MEALS|FROZEN|-80.97058|80.970653784086934|204|1
35.03469|f7165cfc4b5774317c620d321d7e521f3a5a4815|2.49|2014-09-29 09:17:00|80.970590786568081|4|1380017219|82|35.079009695900304|0|55|1278|-80.85753|48|35.116638|SINGLE SERVE NUTRITIONAL|0.0|5|LC SPAGHETTI MEAT SAUCE|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00013800166357|FROZEN MEALS|FROZEN|-80.97058|80.970653784086934|204|1
35.03469|d422328ef44b33c316f14c932275ad2616d43935|4.98|2014-10-02 09:53:00|80.970590786568081|4|1380017219|82|35.079009695900304|0|55|1278|-80.85753|48|35.116638|SINGLE SERVE NUTRITIONAL|0.98|5|LC SPAGHETTI MEAT SAUCE|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00013800166357|FROZEN MEALS|FROZEN|-80.97058|80.970653784086934|204|2
35.03469|0219f8a8d17673c323cd3ff53e3d8eb49a61990c|6.5|2014-11-10 20:29:00|80.970590786568081|4|4127102564|82|35.079009736394411|0|55|341|-80.994596|57|35.061685|CREAMERS|0.5|3|ITNAT'L FRENCH VANILLA|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00041271025644|MILK|DAIRY|-80.97058|80.97058935057278|475|2
35.03469|aa7397691b26d3169798c21f340d2d8af7ecfefa|7.99|2015-01-01 15:35:00|80.970590786568081|4|4775478492|82|35.079009736394411|0|55|6424|-80.994596|1556|35.061685|GAMES|0.0|18|LIC 5IN1 GAME TRAVEL CASE ASST|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00047754784923|TOYS|GM|-80.97058|80.97058935057278|475|1
35.03469|4728612c8643d3997af8b7615e1affa1e7c66d45|3.99|2014-11-08 16:36:00|80.970590786568081|4|7835470843|82|35.07900972860665|0|55|317|-80.992182|52|35.103409|CHUNK AND BAR CHEESE|1.49|3|CABOT EXTRA SHARP WHITE CHEDD|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00078354703182|CHEESE|DAIRY|-80.97058|80.970613430786784|88|1
35.03469|094b66d6fd820c096f1646f5ef342328d7411840|15.49|2014-11-27 12:29:00|80.970590786568081|4|7116005579|82|35.079009736394411|0|55|5811|-80.994596|1534|35.061685|GLASS OVENWARE|0.0|18|PYREX EASY GRAB 3QT OBLONG/CVR|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00071160055797|MEATAL/GLASS BAKEWARE|GM|-80.97058|80.97058935057278|475|1
35.03469|4f58db4935b1b454d58331a996f68434a9172ad0|3.48|2015-01-22 21:03:00|80.970590786568081|4||82|35.079009736394411|0|55|536|-80.994596|64|35.061685|FRESH SQUASH|0.0|4|SPAGHETTI SQUASH|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00204776000008|FRESH PRODUCE|PRODUCE|-80.97058|80.97058935057278|475|1
35.03469|319a1d4e7ee27a624e3e687b3962a535c98235f3|9.3|2015-02-01 19:18:00|80.970590786568081|4|7218063473|82|35.079009736394411|0|55|254|-80.994596|892|35.061685|PREMIUM PIZZA|2.63|5|RED BARON THN CRUST 5 CHEESE|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00072180633217|FROZEN PIZZA|FROZEN|-80.97058|80.97058935057278|475|2
35.03469|911ec647168e4391a945440ca367ddc7de7dcafb|5.78|2015-01-28 11:52:00|80.970590786568081|4|5100019922|82|35.079009736394411|0|55|1261|-80.994596|274|35.061685|MEAL STARTERS|0.0|1|CAMP SKILLETS THAI CUR LMGRASS|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00051000199263|PREP FOODS DINNERS|G1 GROCERY|-80.97058|80.97058935057278|475|2
35.03469|56aa983dd286902b5971a05fc14b6b4f7092832d|2.29|2014-09-10 08:13:00|80.970590786568081|4|1620033500|82|35.079009736394411|0|55|225|-80.994596|35|35.061685|SUGAR-GRANULATED|0.0|1|DIXIE CRYSTAL SUGAR GRANULATE|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00016200335002|SUGAR/SUBSTITUTES|G1 GROCERY|-80.97058|80.97058935057278|475|1
35.03469|54e49036c362d0026f5f3f8ad01a97bacb237843|2.99|2015-02-25 17:03:00|80.970590786568081|4|4470036113|82|35.079009736394411|0|55|659|-80.994596|103|35.061685|CHILDRENS LUNCH SNACKS|0.0|19|FUNPACK LUNCHABLE NACHO|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00044700006795|LUNCH SNACKS|CASE READY MEATS|-80.97058|80.97058935057278|475|1
35.03469|a37ec4829bbb5dd5ad3bcba7f7c88ae2877a4097|2.31|2015-01-31 09:16:00|80.970590786568081|4||82|35.079009736394411|0|55|536|-80.994596|64|35.061685|FRESH SQUASH|0.0|4|COO ZUCCHINI SQUASH, FANCY|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00204067000007|FRESH PRODUCE|PRODUCE|-80.97058|80.97058935057278|475|1
35.03469|6bba59881ea6aad72fad4d718c644df3524c5d21|14.99|2014-11-01 15:28:00|80.970590786568081|4|62901400609|82|35.079009736394411|0|55|1703|-80.994596|387|35.061685|SEASONAL COOKIES|5.0|14|EZ BUILD GINGERBREAD HOUSE KIT|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00629014006091|COOKIES|BAKERY|-80.97058|80.97058935057278|475|1
35.03469|d038a181074d7668ef3d389c1e08d3da6ec6e0e5|0.76|2015-02-25 13:55:00|80.970590786568081|4||82|35.079009736394411|0|55|558|-80.994596|64|35.061685|SPECIALTY-VEGETABLES|0.0|4|COO GINGER ROOT, BULK|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00204612000001|FRESH PRODUCE|PRODUCE|-80.97058|80.97058935057278|475|1
35.03469|15ef8415491377899927f824b48ea9b0dce9f87e|1.48|2014-10-04 16:51:00|80.970590786568081|4||82|35.07900972860665|0|55|558|-80.992182|64|35.103409|SPECIALTY-VEGETABLES|0.0|4|COO GINGER ROOT, BULK|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00204612000001|FRESH PRODUCE|PRODUCE|-80.97058|80.970613430786784|88|1
35.03469|f0e0e4dc231bf5b0fe10ac3d7cccb2a909851d96|2.29|2015-02-28 19:25:00|80.970590786568081|4|7203663996|82|35.079009736394411|0|55|342|-80.994596|57|35.061685|FRESH MILK|0.0|3|HARRIS TEETER FF SKIM MILK|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00072036631299|MILK|DAIRY|-80.97058|80.97058935057278|475|1
35.03469|00975ff4df8071b707093c4205dbb67670499065|3.49|2015-02-14 16:09:00|80.970590786568081|4|7203663995|82|35.079009736394411|0|55|342|-80.994596|57|35.061685|FRESH MILK|0.0|3|HARRIS TEETER 1/2% MILK GALL|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00072036632012|MILK|DAIRY|-80.97058|80.97058935057278|475|1
35.03469|eb31bec48d7e28cfbe2744aebb762f62bf65458e|3.79|2014-09-10 21:45:00|80.970590786568081|4|7203688184|82|35.079009736394411|0|55|555|-80.994596|64|35.061685|PACKAGED SALADS|0.0|4|HTT ASIAN CHOP SALAD KIT|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00072036881847|FRESH PRODUCE|PRODUCE|-80.97058|80.97058935057278|475|1
35.03469|ee3c67dc6b5941f7891380aadc0a37be7cf6ff7f|4.5|2014-11-23 13:54:00|80.970590786568081|4||82|35.079009736394411|0|55|1617|-80.994596|373|35.061685|ROLLS BULK|0.0|14|BULK ROLLS|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00072036955555|ROLLS|BAKERY|-80.97058|80.97058935057278|475|6
35.03469|0a1d81cc0275f72c7cb00acd2891dc00c4e4cc31|1.79|2015-02-10 14:20:00|80.970590786568081|4|7203663157|82|35.079009736394411|0|55|1134|-80.994596|57|35.061685|CARTON MILK|0.0|3|HARRIS TEETER 2% MILK|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00072036631558|MILK|DAIRY|-80.97058|80.97058935057278|475|1
35.03469|ee8958c36cbfdd6f16f194e6983851f4305517de|9.99|2014-11-14 16:54:00|80.970590786568081|4|8427997505|82|35.079009687878134|0|55|9952|-80.806073|886|35.106477|NFS-PREM-PINOT NOIR|0.0|13|LE GRAND PINOT NOIR|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00084279975054|PREMIUM ($8-$10.99)|WINE|-80.97058|80.970660655328672|4|1
35.03469|9310151425118a62e65b2f83b5ce0d65a427eef4|1.87|2015-01-16 22:43:00|80.970590786568081|4|7433610205|82|35.079009736394411|0|55|317|-80.994596|52|35.061685|CHUNK AND BAR CHEESE|0.0|3|HC SHARP CHEDDAR CHEESE|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00074336102059|CHEESE|DAIRY|-80.97058|80.97058935057278|475|1
35.03469|62648c9aff1c627876dab1da0e4dfffd3c0a59cb|9.99|2014-11-28 17:25:00|80.970590786568081|4|1098600250|82|35.079009687878134|0|55|9961|-80.806073|887|35.106477|NFS-S/PREM-MERLOT|0.0|13|KENWOOD MERLOT|3d4c88e4407ba924d8134d1115779175eab2ba70|3.062386802192842|35.077427448337218|00010986002509|SUPER PREMIUM ($11-$14.99)|WINE|-80.97058|80.970660655328672|4|1
35.40953|6bd98d57009020f29538b72a0efb8a5dc44a75df|1.49|2015-02-14 11:38:00|1.4102725052409182|1|4133102785|209|0.6180128850837077|0|1|1214|-80.86175|272|35.40953|AUTHENTIC HISPANIC|0.0|1|GOYA WATER COCONUT|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00041331027854|HISPANIC PREP. FOODS|G1 GROCERY|-80.86175|1.4113037764245249|209|1
35.40953|b3f0210d69bdb736c8b9c046c8a08f743918878a|3.59|2015-02-01 09:16:00|1.4102725052409182|1|4116400022|209|0.6180128850837077|0|1|1469|-80.86175|278|35.40953|REGULAR CUT FRIES|0.59|5|MRS T'S POT/4 CHS MINI PIEROGI|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00041164008419|FROZEN POTATO|FROZEN|-80.86175|1.4113037764245249|209|1
35.40953|8ed874e312673c7213cf0e4f68544a183f056724|2.49|2015-02-21 14:18:00|80.86161257435397|1|4112939640|209|35.433889672079935|1|36|1219|-80.8955|275|35.4437|PASTA SC CORE|0.0|1|CLASSICO PIZZA SAUCE|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|35.472272108304431|00041129396407|PASTA SAUCES|G1 GROCERY|-80.86175|80.861756012753958|272|1
35.40953|28b08690d73c16f2bee4f2c357d066bb40a71e1c|4.19|2015-01-18 10:48:00|1.4102725052409182|1|3800031846|209|0.6180128850837077|0|1|81|-80.86175|9|35.40953|RTE CEREAL KIDS|0.0|1|KELL COCOA KRISPIES|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00038000768620|CEREAL|G1 GROCERY|-80.86175|1.4113037764245249|209|1
35.40953|b28be19494799e504bf26383653cc6414c0c253a|3.49|2015-02-07 09:13:00|1.4102725052409182|1|3800001611|209|0.6180128850837077|0|1|61|-80.86175|9|35.40953|RTE CEREAL ADULT|0.0|1|KELLOGG SPECIAL K RED BERRIES|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00038000599231|CEREAL|G1 GROCERY|-80.86175|1.4113037764245249|209|1
35.40953|38a05060c0ca332d89b3026b90a0e6f9e1d955ff|4.99|2014-09-13 15:57:00|1.4102725052409182|1|4082201114|209|0.6180128850837077|0|1|1878|-80.86175|435|35.40953|HUMMUS|0.0|6|HUMMUS W/ ROASTED PINE NUTS|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00040822011747|SALADS|DELI|-80.86175|1.4113037764245249|209|1
35.40953|2b9a02082b123c9d9f13b287b5d28ac5b7ee8c9a|3.39|2015-01-24 08:45:00|1.4102725052409182|1|3800031829|209|0.6180128850837077|0|1|74|-80.86175|9|35.40953|RTE CEREAL ALL FAMILY|0.89|1|KELL MIN WH STRAWBERRY|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00038000576362|CEREAL|G1 GROCERY|-80.86175|1.4113037764245249|209|1
35.40953|f066475b6ee4785bee6217c2bc9d6b433b8595e7|3.39|2014-12-07 09:04:00|1.4102725052409182|1|3800031829|209|0.6180128850837077|0|1|74|-80.86175|9|35.40953|RTE CEREAL ALL FAMILY|0.0|1|KELL MIN WH STRAWBERRY|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00038000576362|CEREAL|G1 GROCERY|-80.86175|1.4113037764245249|209|1
35.40953|773c9d008a5675c0332bfcc52e3b0bb839cb614a|4.19|2014-12-14 09:40:00|1.4102725052409182|1|3800031846|209|0.6180128850837077|0|1|81|-80.86175|9|35.40953|RTE CEREAL KIDS|1.69|1|KELL COCOA KRISPIES|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00038000768620|CEREAL|G1 GROCERY|-80.86175|1.4113037764245249|209|1
35.40953|fc79e4169e9eff481f527b92cd8b3b477d1c94e4|2.35|2015-01-03 10:12:00|1.4102725052409182|1|4112907700|209|0.6180128850837077|0|1|1219|-80.86175|275|35.40953|PASTA SC CORE|0.35|1|CLASSICO SC SPICY RED PEPPER|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00041129077429|PASTA SAUCES|G1 GROCERY|-80.86175|1.4113037764245249|209|1
35.40953|12001709bf5ef7ab6711d25ebea9752b841fd1c0|3.39|2014-11-15 09:07:00|1.4102725052409182|1|3800031829|209|0.6180128850837077|0|1|74|-80.86175|9|35.40953|RTE CEREAL ALL FAMILY|0.0|1|KELL MIN WH STRAWBERRY|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00038000576362|CEREAL|G1 GROCERY|-80.86175|1.4113037764245249|209|1
35.40953|18b75643185c0eb9a36bb86810f462f4b90bc4bc|3.19|2015-03-08 09:31:00|1.4102725052409182|1|1600027532|209|0.6180128850837077|0|1|81|-80.86175|9|35.40953|RTE CEREAL KIDS|1.6|1|GM TRIX|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00016000275324|CEREAL|G1 GROCERY|-80.86175|1.4113037764245249|209|1
35.40953|27b31035c3a76eb34c19592a31c04e7a0c21eb95|1.07|2014-09-28 14:33:00|1.4102725052409182|1||209|0.6180128850837077|0|1|502|-80.86175|64|35.40953|FRESH BANANAS|0.0|4|BANANAS, YELLOW|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.86175|1.4113037764245249|209|1
35.40953|83174fd52656e98024ab8ce3c645e49c50434ff6|1.76|2014-09-20 09:36:00|1.4102725052409182|1||209|0.6180128850837077|0|1|502|-80.86175|64|35.40953|FRESH BANANAS|0.0|4|BANANAS, YELLOW|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.86175|1.4113037764245249|209|1
35.40953|8df2d0c9b27b6f01650678c9b9f7b364e9cd485e|1.53|2014-11-24 17:42:00|1.4102725052409182|1||209|0.6180128850837077|0|1|502|-80.86175|64|35.40953|FRESH BANANAS|0.0|4|BANANAS, YELLOW|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.86175|1.4113037764245249|209|1
35.40953|281c4cffcd16a5b5bedd2393a91249bbdf723b4d|0.9|2014-12-30 17:22:00|1.4102725052409182|1||209|0.6180128850837077|0|1|502|-80.86175|64|35.40953|FRESH BANANAS|0.0|4|BANANAS, YELLOW|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00204011000008|FRESH PRODUCE|PRODUCE|-80.86175|1.4113037764245249|209|1
35.40953|2648e83c350af18a2a1dd4121c6e1a433d90b4f5|3.99|2015-03-01 09:08:00|1.4102725052409182|1|4610000012|209|0.6180128850837077|0|1|318|-80.86175|52|35.40953|SHREDDED/GRATED CHEESE|2.0|3|SARGENTO OTB MOZZ TRAD CUT|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00046100000120|CHEESE|DAIRY|-80.86175|1.4113037764245249|209|1
35.40953|626a0c09d42b2ef2eafedcf2dcfb97e7f41c8b1f|3.89|2014-10-02 15:36:00|1.4102725052409182|1|3800039118|209|0.6180128850837077|0|1|81|-80.86175|9|35.40953|RTE CEREAL KIDS|1.9|1|KELLOGG APPLE JACKS 12.2|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00038000391347|CEREAL|G1 GROCERY|-80.86175|1.4113037764245249|209|1
35.40953|b5903658aedd3e496f3cec3ab28513662e863922|7.97|2015-02-09 21:32:00|1.4102725052409182|1|4116706651|209|0.6180128850837077|0|1|3202|-80.86175|1015|35.40953|HAND & BODY THERAPEUTIC|0.0|17|GOLD BOND ULT HEALING LOTION|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00041167066515|HAND & BODY LOTION/SUN CARE|HBC|-80.86175|1.4113037764245249|209|1
35.40953|41e7608a78902d7ab0924a48c12943c69ca5c904|3.98|2014-11-26 08:39:00|1.4102725052409182|1|3900004504|209|0.6180128850837077|0|1|114|-80.86175|14|35.40953|PUMPKIN|0.4|1|LIBBY SOLID PACK PUMPKIN|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00039000045049|DESSERTS/GELS/SYRUPS|G1 GROCERY|-80.86175|1.4113037764245249|209|2
35.40953|b23f14b8e100ecb776cebb7ff5a5bf89559a8d03|3.99|2014-12-21 12:53:00|1.4102725052409182|1|3800005220|209|0.6180128850837077|0|1|81|-80.86175|9|35.40953|RTE CEREAL KIDS|0.0|1|KELLOGG FUN PACK 8 CT|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00038000052200|CEREAL|G1 GROCERY|-80.86175|1.4113037764245249|209|1
35.40953|65520d7e858fef28889a2b2eee13de61399e2176|4.59|2014-10-01 22:08:00|1.4102725052409182|1|3800059661|209|0.6180128850837077|0|1|61|-80.86175|9|35.40953|RTE CEREAL ADULT|0.0|1|KELLOGG RAISIN BRAN 23|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00038000596612|CEREAL|G1 GROCERY|-80.86175|1.4113037764245249|209|1
35.40953|7f356b08225caeec1da2f64ba03db9124e2cc861|3.99|2014-09-23 16:54:00|1.4102725052409182|1|3800005220|209|0.6180128850837077|0|1|81|-80.86175|9|35.40953|RTE CEREAL KIDS|0.0|1|KELLOGG FUN PACK 8 CT|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00038000052200|CEREAL|G1 GROCERY|-80.86175|1.4113037764245249|209|1
35.40953|a40d657b17c391ede5cd7e60fbeedec0486e4eee|3.99|2014-11-23 09:46:00|1.4102725052409182|1|7203688076|209|0.6180128850837077|0|1|523|-80.86175|64|35.40953|FRESH POTATOES|0.49|4|HT RUSSET POTATO 5LB BAG|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00072036880765|FRESH PRODUCE|PRODUCE|-80.86175|1.4113037764245249|209|1
35.40953|842b71dc6152d182a09a4a6e1b83ecb20c1e8a77|3.99|2015-02-18 21:03:00|1.4102725052409182|1|3338300005|209|0.6180128850837077|0|1|500|-80.86175|64|35.40953|FRESH APPLES|0.0|4|RED DEL APPLE 3LB BAG|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00072036880116|FRESH PRODUCE|PRODUCE|-80.86175|1.4113037764245249|209|1
35.40953|4ccd7a11603e4d72b511668be214d046777dcec2|5.91|2015-02-12 16:48:00|1.4102725052409182|1|7203656070|209|0.6180128850837077|0|1|316|-80.86175|52|35.40953|CREAM CHEESE|1.41|3|HT LIGHT CREAM CHEESE|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00072036560742|CHEESE|DAIRY|-80.86175|1.4113037764245249|209|3
35.40953|f6968cbd9b0ba7fa200eef26c22d7bddf450088b|6.27|2015-02-25 16:47:00|1.4102725052409182|1|7203676359|209|0.6180128850837077|0|1|345|-80.86175|57|35.40953|ORGANIC MILK|0.0|3|HTO ORGANIC 1% MILK GAL|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00072036763617|MILK|DAIRY|-80.86175|1.4113037764245249|209|1
35.40953|05d9124f1cf217b9a5cad3974033f7a8ce66766a|5.49|2014-10-05 10:32:00|1.4102725052409182|1|7203670737|209|0.6180128850837077|0|1|202|-80.86175|31|35.40953|PRETZELS|0.49|1|HTT PNUT BTR FILL PRETZL|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00072036707376|SNACKS|G1 GROCERY|-80.86175|1.4113037764245249|209|1
35.40953|461720be4e98bb779cbe01618e763a07c4bd1b99|6.58|2015-01-31 13:31:00|1.4102725052409182|1|2840004768|209|0.6180128850837077|0|1|202|-80.86175|31|35.40953|PRETZELS|1.58|1|ROLD GOLD RODS PRETZELS|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00028400012348|SNACKS|G1 GROCERY|-80.86175|1.4113037764245249|209|2
35.40953|cccb363787636fd9449e0053f058a7abb65affaa|1.39|2014-11-09 09:25:00|1.4102725052409182|1|6414404551|209|0.6180128850837077|0|1|179|-80.86175|27|35.40953|CANNED PASTA|0.39|1|CBRD WG BEEFARONI|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00064144041336|PREPARED FOODS-RTS|G1 GROCERY|-80.86175|1.4113037764245249|209|1
35.40953|a03d89ac84cd24895d773a57645e625f466cb4d5|4.99|2015-02-18 16:35:00|1.4102725052409182|1|7203688138|209|0.6180128850837077|0|1|500|-80.86175|64|35.40953|FRESH APPLES|0.0|4|HT CRIPPS PINK APPLE 3LB|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00072036881380|FRESH PRODUCE|PRODUCE|-80.86175|1.4113037764245249|209|1
35.40953|0db50b8b1212fdd83b09c05fe02a67417751041d|4.99|2014-11-20 12:01:00|1.4102725052409182|1|3700039316|209|0.6180128850837077|0|1|726|-80.86175|73|35.40953|NFS-BODY WASHES|1.0|1|OLD SPC FRESH COL FIJI BDYWASH|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00037000267904|PERSONAL SOAP/BATH ADDITIVES|G1 GROCERY|-80.86175|1.4113037764245249|209|1
35.40953|3c3f55389abc3afd6fd4c1d724e7baad528900fb|8.19|2014-10-11 08:21:00|1.4102725052409182|1|2840000288|209|0.6180128850837077|0|1|205|-80.86175|31|35.40953|REMAINING SNACKS|1.2|1|FRITOLAY CLASSIC 20 CTN|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00028400002882|SNACKS|G1 GROCERY|-80.86175|1.4113037764245249|209|1
35.40953|441fa318e36f1b08cfe543bbc90ecd7f2f4fec34|6.97|2014-12-06 20:13:00|1.4102725052409182|1|1150904933|209|0.6180128850837077|0|1|3965|-80.86175|1075|35.40953|HAIR COLORING-MEN|0.0|17|JFM DRK BROWN FACIAL HAIRCOLOR|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00011509049049|SHAVING NEEDS/MEN HAIR|HBC|-80.86175|1.4113037764245249|209|1
35.40953|d20a20ac090b15d06b4aba62f7e76b02b6287650|3.19|2015-01-30 19:19:00|1.4102725052409182|1|9396681150|209|0.6180128850837077|0|1|364|-80.86175|55|35.40953|ORGANIC AND CF EGGS|0.0|3|ORGANIC VALLEY XTRA LARGE EGGS|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00093966811506|EGGS FRESH|DAIRY|-80.86175|1.4113037764245249|209|1
35.40953|c2c492ca44864aedf62026ced4b6e1ab70de6487|3.99|2014-09-26 18:25:00|1.4102725052409182|1|7203602701|209|0.6180128850837077|0|1|1878|-80.86175|435|35.40953|HUMMUS|0.5|6|FFM ARTISAN RED PEPPER HUMMUS|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00072036027030|SALADS|DELI|-80.86175|1.4113037764245249|209|1
35.40953|42bd873c3fb2ea2b2881df199a8b8a0401554f69|1.29|2014-10-09 12:33:00|1.4102725052409182|1|7203670782|209|0.6180128850837077|0|1|725|-80.86175|66|35.40953|NFS-DISHWASHING LIQUID|0.4|1|YH LIQ DISH ORIGINAL 10 OZ|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00072036707826|DETERGENTS|G1 GROCERY|-80.86175|1.4113037764245249|209|1
35.40953|abfacdede8874d9e3507ece36d4b04563ad46de0|1.99|2014-12-20 13:21:00|1.4102725052409182|1|3400000007|209|0.6180128850837077|0|1|48|-80.86175|7|35.40953|REGISTER GUM|0.0|1|ICE BREAKER WINTERGREEN MINTS|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00034000000098|CANDY|G1 GROCERY|-80.86175|1.4113037764245249|209|1
35.40953|baef2bdc9f8efed0db9c2894107a295577707f79|7.99|2014-12-29 21:40:00|1.4102725052409182|1|7203697620|209|0.6180128850837077|0|1|4615|-80.86175|1215|35.40953|VITAMIN-MULTIPLE-ADULT|0.0|17|HT ONE DAILY MENS TABS 97620|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00072036976208|VITAMINS & SUPPLEMENTS|HBC|-80.86175|1.4113037764245249|209|1
35.40953|c8ed8451491fd5099194272323d90f41e9ccc7bc|5.97|2014-11-07 21:09:00|1.4102725052409182|1|7203676359|209|0.6180128850837077|0|1|345|-80.86175|57|35.40953|ORGANIC MILK|0.0|3|HTO ORGANIC FF SKIM GAL|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00072036763624|MILK|DAIRY|-80.86175|1.4113037764245249|209|1
35.40953|ab29e0242bc2f418d3be14c993a07e88b395baab|5.97|2014-10-21 22:16:00|1.4102725052409182|1|7203676359|209|0.6180128850837077|0|1|345|-80.86175|57|35.40953|ORGANIC MILK|0.0|3|HTO ORGANIC FF SKIM GAL|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00072036763624|MILK|DAIRY|-80.86175|1.4113037764245249|209|1
35.40953|3c4c1769712debdc626e68bfc831ec0a27edca11|6.27|2015-03-06 20:42:00|1.4102725052409182|1|7203676359|209|0.6180128850837077|0|1|345|-80.86175|57|35.40953|ORGANIC MILK|0.0|3|HTO ORGANIC FF SKIM GAL|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00072036763624|MILK|DAIRY|-80.86175|1.4113037764245249|209|1
35.40953|ac2d0712d3e6263b032df0d69ad846967b0f0bf7|2.69|2015-02-25 16:52:00|1.4102725052409182|1|1410007660|209|0.6180128850837077|0|1|1031|-80.86175|162|35.40953|ITALIAN|0.0|7|PEP SLICED ITALIAN BRD SD  PP|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00014100076605|SLICED BREAD|COMMERCIAL BAKERY|-80.86175|1.4113037764245249|209|1
35.40953|c15d6768878827d8d9f12aef398369d44cf4e93a|7.38|2014-09-21 10:24:00|1.4102725052409182|1|7127928100|209|0.6180128850837077|0|1|555|-80.86175|64|35.40953|PACKAGED SALADS|0.0|4|F.E. FARMERS GARDEN|40a591ec09cd3340627dbdf5706b92330562806e|1.6831945482722543|0.61833652052202714|00071279281025|FRESH PRODUCE|PRODUCE|-80.86175|1.4113037764245249|209|2
35.096737|24e77c7c589ed59249383c149a9894e542cef7a5|3.79|2015-02-08 17:29:00|80.782094729586973|2|7684010015|30|35.102762219822544|0|27|275|-80.85013|45|35.175855|SUPER PREMIUM ICE CREAM|0.29|5|BEN & JERRY S'MORES|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00076840101771|ICE CREAM|FROZEN|-80.78468|80.784683882857976|218|1
35.096737|be735a0804a3578b6dbe3a4915a6ffd9bad0e5b7|3.89|2014-11-21 12:18:00|80.782094729586973|2|2800011470|30|35.102762218483747|0|27|46|-80.844274|7|35.204336|PKG CHOC|0.0|1|SWEETART CHEWY MINI|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00079200717834|CANDY|G1 GROCERY|-80.78468|80.784686259269677|61|1
35.096737|dd1d8cd6879e16adff59bee640d343456760da7e|2.79|2014-11-26 12:03:00|1.4091206135396188|2|7878390810|30|0.612553617356517|0|47|561|-80.78468|64|35.096737|FR PROD ORGANIC PRODUCE|0.0|4|ORG CARROTS, PETITE 12OZ BAG|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|0.61242566243833529|00078783908103|FRESH PRODUCE|PRODUCE|-80.78468|1.4099586511700126|30|1
35.096737|b864727006c53149adf74649e79999f593de794a|3.79|2014-12-23 11:27:00|1.4091206135396188|2|4850002013|30|0.612553617356517|0|47|335|-80.78468|56|35.096737|ORANGE JUICE-REGRIGERATED|0.79|3|TROPICANA PP W/CALCIUM|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|0.61242566243833529|00048500305690|JUICES & DRINKS-REFRIGERATED|DAIRY|-80.78468|1.4099586511700126|30|1
35.096737|892b1edcd18d59d2e66f9e95c2c2244e16bc7202|1.39|2015-01-06 19:24:00|1.4091206135396188|2|5210076069|30|0.612553617356517|0|47|80|-80.78468|34|35.096737|SEASONING PACKETS|0.0|1|MC GRILL MATE BRW SUGAR BOURBO|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|0.61242566243833529|00052100013848|SPICES/SEASONINGS/EXTRACTS|G1 GROCERY|-80.78468|1.4099586511700126|30|1
35.096737|795f53ebe4e1edb75be8b7e91c548850c8935d15|3.99|2014-12-20 16:58:00|80.782094729586973|2|5783602064|30|35.102762218393444|0|27|522|-80.992182|64|35.103409|FRESH TOMATOES|0.0|4|CAMPARI TOMATO 16 OZ|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00057836020641|FRESH PRODUCE|PRODUCE|-80.78468|80.784686387816123|88|1
35.096737|f34390ce629c3d8a9a5961bff1962b20c377fa44|2.99|2014-10-06 16:24:00|80.782094729586973|2|7203695121|30|35.102762220218196|0|27|1629|-80.849471|373|35.161696|TAKE & BAKE ROLLS|0.0|14|TAKE & BAKE WHEAT PETIT PN RL|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00072036951212|ROLLS|BAKERY|-80.78468|80.784682820269396|35|1
35.096737|ab0fd9bf4d95921b8c1e9cb8d8affe9b8bbd0af8|4.99|2015-01-05 16:30:00|80.782094729586973|2|7203698017|30|35.102762219822544|0|27|1243|-80.85013|21|35.175855|MIXED NUTS CASHEWS|0.5|1|HT SALTED MIXED NUTS|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00072036980175|NUTS|G1 GROCERY|-80.78468|80.784683882857976|218|1
35.096737|01d85295042033165c6dc9dd7bba53b15944cdc2|2.99|2014-12-09 18:38:00|80.782094729586973|2|7203695121|30|35.102762219822544|0|27|1629|-80.85013|373|35.175855|TAKE & BAKE ROLLS|0.0|14|TAKE & BAKE WHEAT PETIT PN RL|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00072036951212|ROLLS|BAKERY|-80.78468|80.784683882857976|218|1
35.096737|1ddbb6f83f62e29438089f77205b4db4468b06ec|6.99|2014-11-08 19:21:00|80.782094729586973|2|89413700203|30|35.102762220614999|0|27|463|-80.85753|84|35.116638|HARD CIDER|0.0|16|CRISPIN CIDER 4PK|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00894137002033|SPECIALTY|BEER|-80.78468|80.78468090022767|204|1
35.096737|000d5d638fa812adfe59046f63a5d50ed9a69ed4|10.99|2014-11-15 09:18:00|80.782094729586973|2|1103450005|30|35.10276222019543|0|27|9983|-80.770346|889|35.052812|NFS-SPARKLING|0.0|13|MARTINI & ROSSI ASTI SPUMANTE|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00011034500053|SPARKLING|WINE|-80.78468|80.784682892026439|40|1
35.096737|4263bac4d8bdf5b87470a56ce52855510d5dbc8e|4.49|2015-01-14 19:28:00|1.4091206135396188|2|4400000430|30|0.612553617356517|0|47|90|-80.78468|13|35.096737|SNACK CRACKERS|0.5|1|WHEAT THINS REDUCED FAT FAMILY|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|0.61242566243833529|00044000004309|CRACKERS|G1 GROCERY|-80.78468|1.4099586511700126|30|1
35.096737|e4566a0f1ded7d0cd51254d9da03528e3c1a1536|2.95|2014-10-20 17:26:00|80.782094729586973|2|4127102591|30|35.102762218483747|0|27|144|-80.844274|229|35.204336|CEAMERS-POWDERED|0.0|1|INT'L DELIGHT CLD STN SWT CRM|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00041271017571|COCOAS CREAMERS SYRUPS|G1 GROCERY|-80.78468|80.784686259269677|61|1
35.096737|c516f92355c5f465ec026e0356617f74863b3a95|3.99|2015-02-03 09:57:00|1.4091206135396188|2|7341001375|30|0.612553617356517|0|47|1026|-80.78468|162|35.096737|WHEAT|0.0|7|ARN 100% WHOLE WHEAT WP  PP|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|0.61242566243833529|00073410013755|SLICED BREAD|COMMERCIAL BAKERY|-80.78468|1.4099586511700126|30|1
35.096737|3d3901a27fd96e55d6e4b9f82b49542fd1d0d47f|10.99|2014-10-16 16:11:00|1.4091206135396188|2|8500001736|30|0.612553617356517|0|47|9939|-80.78468|885|35.096737|NFS POP PINOT NOIR|0.0|13|BAREFOOT PINOT NOIR 1.5L|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|0.61242566243833529|00085000017364|POPULAR (4-$7.99)|WINE|-80.78468|1.4099586511700126|30|1
35.096737|5b99a0b056ae56655ca7a5676fccc2ee7ecb2f4e|10.99|2014-11-29 16:47:00|80.782094729586973|2|8500001736|30|35.102762220463141|0|27|9939|-80.771677|885|35.066546|NFS POP PINOT NOIR|0.0|13|BAREFOOT PINOT NOIR 1.5L|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00085000017364|POPULAR (4-$7.99)|WINE|-80.78468|80.784681882621484|45|1
35.096737|788c07a635eb83a8ccf689d72d3be6d0616a1e2c|9.99|2014-09-23 16:39:00|80.782094729586973|2|8500001736|30|35.102762220659947|0|27|9939|-80.806073|885|35.106477|NFS POP PINOT NOIR|0.0|13|BAREFOOT PINOT NOIR 1.5L|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00085000017364|POPULAR (4-$7.99)|WINE|-80.78468|80.78468003418341|4|1
35.096737|7643e205a29b9f1512ff24cabba362e30cf85121|4.75|2015-01-15 20:24:00|80.782094729586973|2|18685200031|30|35.102762220218196|0|27|275|-80.849471|45|35.161696|SUPER PREMIUM ICE CREAM|0.0|5|TALENTI DBL DRK CHOC GELATO|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00186852000341|ICE CREAM|FROZEN|-80.78468|80.784682820269396|35|1
35.096737|c05ee6b4174d44a7f8cd6427b036e2bc07f2e664|3.49|2014-11-24 17:41:00|80.782094729586973|2|4610000107|30|35.102762218483747|0|27|331|-80.844274|52|35.204336|NATURAL SLICED|0.49|3|SARGENTO MUENSTER CHEESE|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00046100001073|CHEESE|DAIRY|-80.78468|80.784686259269677|61|1
35.096737|549d1385e74e2b78ddf7a665df11c2083d80bcb3|2.35|2014-09-17 20:47:00|80.782094729586973|2|3800030110|30|35.102762218483747|0|27|44|-80.844274|6|35.204336|TOASTER PASTRIES-SHELF STABLE|0.6|1|KELL POPTART BROWN SUGAR|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00038000311109|BREAKFAST FOODS|G1 GROCERY|-80.78468|80.784686259269677|61|1
35.096737|bd05ad4bf322df58430f4fba120c0986295d7a9d|3.49|2014-12-15 16:38:00|80.782094729586973|2|3400000847|30|35.102762220659947|0|27|45|-80.806073|7|35.106477|PEG GUM|0.0|1|ICE BRKRS CUBE SPEARMINT|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00034000008476|CANDY|G1 GROCERY|-80.78468|80.78468003418341|4|1
35.096737|0eb03762e7212307bf3640867ff30848ff525375|4.3|2014-11-01 16:43:00|80.782094729586973|2|3800030110|30|35.102762219822544|0|27|44|-80.85013|6|35.175855|TOASTER PASTRIES-SHELF STABLE|0.3|1|KELL POPTART BROWN SUGAR|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00038000311109|BREAKFAST FOODS|G1 GROCERY|-80.78468|80.784683882857976|218|2
35.096737|df501a6755ac1382463a08c0c2a88f32f8a3ef8c|6.39|2014-10-21 14:49:00|1.4091206135396188|2|4154800385|30|0.612553617356517|0|47|252|-80.78468|45|35.096737|PREMIUM ICE CREAM|3.2|5|EDY'S VANILLA BEAN ICE CREAM|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|0.61242566243833529|00041548003856|ICE CREAM|FROZEN|-80.78468|1.4099586511700126|30|1
35.096737|cca79e77fe975f2099e5158ada0b324c2fa7bddb|3.99|2014-10-10 14:24:00|1.4091206135396188|2|3400000847|30|0.612553617356517|0|47|45|-80.78468|7|35.096737|PEG GUM|0.0|1|ICE BRKRS CUBE SPEARMINT|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|0.61242566243833529|00034000008476|CANDY|G1 GROCERY|-80.78468|1.4099586511700126|30|1
35.096737|4a42a20535a56d2613ff2951e3caa48287a222f7|1.55|2014-10-15 19:29:00|80.782094729586973|2|7203663214|30|35.102762220218196|0|27|330|-80.849471|55|35.161696|EGGS|0.0|3|HT GRADE A    EX-LARGE EGGS|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00072036632142|EGGS FRESH|DAIRY|-80.78468|80.784682820269396|35|1
35.096737|4c5e7b08cbe9b526f9a7aee46787841dc5798207|1.79|2015-02-24 16:48:00|1.4091206135396188|2|7203663214|30|0.612553617356517|0|47|330|-80.78468|55|35.096737|EGGS|0.0|3|HT GRADE A    EX-LARGE EGGS|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|0.61242566243833529|00072036632142|EGGS FRESH|DAIRY|-80.78468|1.4099586511700126|30|1
35.096737|eb585e235e3953a7ded5cebb5ca7bcaf31bdb8f8|0.67|2015-02-16 11:09:00|1.4091206135396188|2|7203698078|30|0.612553617356517|0|47|242|-80.78468|39|35.096737|CANNED BEANS|0.17|1|HT BEANS KIDNEY DARK RED|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|0.61242566243833529|00072036411105|VEGETABLES-CAN/JAR|G1 GROCERY|-80.78468|1.4099586511700126|30|1
35.096737|cd853ed1003d758071be68464fa80217be082ab7|3.25|2014-12-22 18:58:00|80.782094729586973|2|7203656080|30|35.102762220463141|0|27|318|-80.771677|52|35.066546|SHREDDED/GRATED CHEESE|0.0|3|HT FANCY SHRED SWISS CHEESE|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00072036000200|CHEESE|DAIRY|-80.78468|80.784681882621484|45|1
35.096737|5997e23a3188a20771162e8020f00696870dd05f|3.92|2014-11-14 15:42:00|1.4091206135396188|2||30|0.612553617356517|0|47|523|-80.78468|64|35.096737|FRESH POTATOES|1.21|4|COO SWEET POTATOES, BULK|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|0.61242566243833529|00204091000004|FRESH PRODUCE|PRODUCE|-80.78468|1.4099586511700126|30|1
35.096737|9689d021f62a483b84bea69ed572e6a2cc8ef851|1.45|2015-02-23 15:46:00|1.4091206135396188|2||30|0.612553617356517|0|47|502|-80.78468|64|35.096737|FRESH BANANAS|0.0|4|BANANAS, YELLOW|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|0.61242566243833529|00204011000008|FRESH PRODUCE|PRODUCE|-80.78468|1.4099586511700126|30|1
35.096737|6ec1a6d8cec8725e38d090d3854fb32b508e69ab|1.2|2015-02-16 13:27:00|80.782094729586973|2||30|35.102762218483747|0|27|502|-80.844274|64|35.204336|FRESH BANANAS|0.0|4|BANANAS, YELLOW|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00204011000008|FRESH PRODUCE|PRODUCE|-80.78468|80.784686259269677|61|1
35.096737|6afe8fc71c34d7fc8915d2bc2df7993c1bb661ff|1.33|2014-09-30 21:07:00|80.782094729586973|2||30|35.102762220218196|0|27|502|-80.849471|64|35.161696|FRESH BANANAS|0.0|4|BANANAS, YELLOW|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00204011000008|FRESH PRODUCE|PRODUCE|-80.78468|80.784682820269396|35|1
35.096737|122718517a6b3553fb2acd3af0320bef735e8fd7|0.94|2015-02-01 14:03:00|80.782094729586973|2||30|35.102762220659947|0|27|502|-80.806073|64|35.106477|FRESH BANANAS|0.0|4|BANANAS, YELLOW|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00204011000008|FRESH PRODUCE|PRODUCE|-80.78468|80.78468003418341|4|1
35.096737|256573f5d632dae6be0f2ed8ab58bc19cf25b663|0.88|2014-11-10 17:46:00|80.782094729586973|2||30|35.102762219822544|0|27|502|-80.85013|64|35.175855|FRESH BANANAS|0.0|4|BANANAS, YELLOW|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00204011000008|FRESH PRODUCE|PRODUCE|-80.78468|80.784683882857976|218|1
35.096737|94a0a2c52d7e7b7c03969491be44f539dedab3eb|1.5|2015-01-12 16:50:00|80.782094729586973|2||30|35.102762220659947|0|27|502|-80.806073|64|35.106477|FRESH BANANAS|0.0|4|BANANAS, YELLOW|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00204011000008|FRESH PRODUCE|PRODUCE|-80.78468|80.78468003418341|4|1
35.096737|2e5a37354da45c019083e6d8cc362da7517079ae|1.16|2015-03-06 19:57:00|80.782094729586973|2||30|35.102762219822544|0|27|502|-80.85013|64|35.175855|FRESH BANANAS|0.0|4|BANANAS, YELLOW|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00204011000008|FRESH PRODUCE|PRODUCE|-80.78468|80.784683882857976|218|1
35.096737|35a3a92f1aec95f1ef537881568ac3a89a8cd7c0|1.1|2015-01-31 18:47:00|80.782094729586973|2||30|35.102762220218196|0|27|502|-80.849471|64|35.161696|FRESH BANANAS|0.0|4|BANANAS, YELLOW|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00204011000008|FRESH PRODUCE|PRODUCE|-80.78468|80.784682820269396|35|1
35.096737|464f804f6ebc06bfddda4ae6869a83231b33ee3c|1.53|2015-01-05 18:46:00|80.782094729586973|2||30|35.102762219822544|0|27|502|-80.85013|64|35.175855|FRESH BANANAS|0.0|4|BANANAS, YELLOW|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00204011000008|FRESH PRODUCE|PRODUCE|-80.78468|80.784683882857976|218|1
35.096737|8c12a96445c001b4009a307e1f7ec9594708b709|1.39|2014-09-16 13:30:00|80.782094729586973|2|1500007607|30|35.102762220463141|0|27|6|-80.771677|1|35.066546|JARRED BABY FOOD|0.32|1|GERBER 2ND APPL W/CHERIES|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00015000073206|BABY FOOD|G1 GROCERY|-80.78468|80.784681882621484|45|1
35.096737|d4927c18b734e6759d2b2b88bb9a463b307ca141|2.69|2015-02-10 16:14:00|80.782094729586973|2|1450000253|30|35.102762219823973|0|27|1273|-80.816172|50|35.059823|BAG VEG NON STEAM|1.35|5|BE ASPARAGUS STIR FRY|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00014500505033|VEGETABLES-FROZEN|FROZEN|-80.78468|80.784683879540324|66|1
35.096737|48d2b7bc167d914b13d1a43f9b316005577cdf33|1.59|2014-12-05 12:14:00|80.782094729586973|2|78142100127|30|35.102762218483747|0|27|1601|-80.844274|371|35.204336|BRANDED BREAD|0.0|14|LA BREA FRENCH DEMI BAGUETTE|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00781421001271|BREAD|BAKERY|-80.78468|80.784686259269677|61|1
35.096737|3cc58031ff644de4743f74709964c50732086bc3|3.99|2014-12-22 14:03:00|80.782094729586973|2|4400002854|30|35.102762218393444|0|27|1248|-80.992182|12|35.103409|SANDWICH COOKIES|1.49|1|OREO DOUBLE STUFF|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00044000028541|COOKIES|G1 GROCERY|-80.78468|80.784686387816123|88|1
35.096737|adf78bd5a25dbc1d37d675f3dbb21d1e4c416eb9|6.5|2015-01-27 13:27:00|80.782094729586973|2|4157005617|30|35.102762218483747|0|27|1265|-80.844274|57|35.204336|ALMOND MILK|0.75|3|ALMOND BREEZE ORIGINAL|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00041570056172|MILK|DAIRY|-80.78468|80.784686259269677|61|2
35.096737|e814e9f0208d1dd0b5d606b8c88512d2b9dd10ab|6.5|2014-12-23 18:30:00|80.782094729586973|2|4157005617|30|35.102762219822544|0|27|1265|-80.85013|57|35.175855|ALMOND MILK|0.75|3|ALMOND BREEZE ORIGINAL|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00041570056172|MILK|DAIRY|-80.78468|80.784683882857976|218|2
35.096737|69ed321a8f7ed4a69b42bd653554105459e6dee5|3.25|2014-09-24 20:05:00|80.782094729586973|2|4157005617|30|35.102762219822544|0|27|1265|-80.85013|57|35.175855|ALMOND MILK|0.0|3|ALMOND BREEZE ORIGINAL|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00041570056172|MILK|DAIRY|-80.78468|80.784683882857976|218|1
35.096737|43a060b84f3a304945172de07324594abc8c0a37|6.39|2015-01-01 12:22:00|1.4091206135396188|2|4154800385|30|0.612553617356517|0|47|252|-80.78468|45|35.096737|PREMIUM ICE CREAM|1.51|5|EDY'S SLOW CHURNED  VANILLA|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|0.61242566243833529|00041548001869|ICE CREAM|FROZEN|-80.78468|1.4099586511700126|30|1
35.096737|accb1b9fd6d7d43dcabbcef333d7bc5030c343da|5.62|2014-11-01 19:29:00|1.4091206135396188|2||30|0.612553617356517|0|47|522|-80.78468|64|35.096737|FRESH TOMATOES|0.0|4|RED H/H TOMATOES, BULK|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|0.61242566243833529|00204799000009|FRESH PRODUCE|PRODUCE|-80.78468|1.4099586511700126|30|1
35.096737|8bac05acc241a3df64c558b0775416263d83c55c|3.29|2015-01-26 15:58:00|80.782094729586973|2|4000024947|30|35.102762218483747|0|27|52|-80.844274|7|35.204336|PKG NON CHOC|0.79|1|STARBURST ORIGINAL FRUITS|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00040000249474|CANDY|G1 GROCERY|-80.78468|80.784686259269677|61|1
35.096737|032b1b56507db4c7f1ac429827fe8a8f0b5bdef2|8.99|2015-03-01 12:36:00|1.4091206135396188|2|2400039329|30|0.612553617356517|0|47|578|-80.78468|136|35.096737|FRESH JARRED FRUIT|0.0|4|DM RED GRAPEFRUIT 64OZ|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|0.61242566243833529|00024000393290|OTHER MERCHANDISE|PRODUCE|-80.78468|1.4099586511700126|30|1
35.096737|d04fe6e2df5ddfa788c5c0f233533991fc05fa8e|3.97|2014-09-21 18:13:00|1.4091206135396188|2|7203663218|30|0.612553617356517|0|47|330|-80.78468|55|35.096737|EGGS|0.0|3|(U)HT LARGE GRADE A LARGE EGGS|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|0.61242566243833529|00072036632180|EGGS FRESH|DAIRY|-80.78468|1.4099586511700126|30|1
35.096737|3dcac83a730d589d238511127395eb027fabbd48|6.39|2014-12-10 15:44:00|1.4091206135396188|2|4154800385|30|0.612553617356517|0|47|252|-80.78468|45|35.096737|PREMIUM ICE CREAM|3.19|5|EDY'S LIGHT VANILLA BEAN|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|0.61242566243833529|00041548003863|ICE CREAM|FROZEN|-80.78468|1.4099586511700126|30|1
35.096737|d659876b9ef3c17dcc839eb194d2503eb4030d4d|6.5|2015-02-17 14:53:00|80.782094729586973|2|4157005617|30|35.102762219822544|0|27|1265|-80.85013|57|35.175855|ALMOND MILK|1.5|3|ALMOND BREEZE UNSWEET ORIGINAL|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00041570056707|MILK|DAIRY|-80.78468|80.784683882857976|218|2
35.096737|c7ffd4c896db8562c7ab0655abc5995456116fe4|1.45|2014-09-25 18:13:00|1.4091206135396188|2|7203663220|30|0.612553617356517|0|47|330|-80.78468|55|35.096737|EGGS|0.0|3|HT GRADE A    LARGE EGGS|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|0.61242566243833529|00072036632203|EGGS FRESH|DAIRY|-80.78468|1.4099586511700126|30|1
35.096737|ec615a28ec0d1d4d16643d290d78b1b6726d9df3|4.99|2015-01-08 14:21:00|80.782094729586973|2|3000006442|30|35.102762218483747|0|27|61|-80.844274|9|35.204336|RTE CEREAL ADULT|0.0|1|QUAKER OATMEAL SQ BROWN SUG|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00030000064412|CEREAL|G1 GROCERY|-80.78468|80.784686259269677|61|1
35.096737|e7f4fc24dbdca83774199376da06f87ffa172b18|5.49|2014-11-19 12:19:00|80.782094729586973|2|88513162808|30|35.102762219822544|0|27|5164|-80.85013|1300|35.175855|PACIFIER|0.0|17|NUK TRNDLINE W/B SILI PAC SZ1|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00885131628091|BABY ACCESSORY|HBC|-80.78468|80.784683882857976|218|1
35.096737|1630537c45803f31ce5dd7e93d372c6a1bb5a383|10.99|2014-12-26 12:44:00|80.782094729586973|2|1008610047|30|35.102762218903614|0|27|9983|-80.80146|889|35.17739|NFS-SPARKLING|0.0|13|CB-RIONDO PROSECCO 750ml|4393c53a2bd19d6352d3f144e3e4c8c985e8fda2|0.4163281972199689|35.102887530186244|00010086100471|SPARKLING|WINE|-80.78468|80.784685623149485|208|1